magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -4931 1140 4931 1174
rect -4931 -1140 -4897 1140
rect 4897 -1140 4931 1140
rect -4931 -1174 4931 -1140
<< nmos >>
rect -4767 -1000 -4737 1000
rect -4671 -1000 -4641 1000
rect -4575 -1000 -4545 1000
rect -4479 -1000 -4449 1000
rect -4383 -1000 -4353 1000
rect -4287 -1000 -4257 1000
rect -4191 -1000 -4161 1000
rect -4095 -1000 -4065 1000
rect -3999 -1000 -3969 1000
rect -3903 -1000 -3873 1000
rect -3807 -1000 -3777 1000
rect -3711 -1000 -3681 1000
rect -3615 -1000 -3585 1000
rect -3519 -1000 -3489 1000
rect -3423 -1000 -3393 1000
rect -3327 -1000 -3297 1000
rect -3231 -1000 -3201 1000
rect -3135 -1000 -3105 1000
rect -3039 -1000 -3009 1000
rect -2943 -1000 -2913 1000
rect -2847 -1000 -2817 1000
rect -2751 -1000 -2721 1000
rect -2655 -1000 -2625 1000
rect -2559 -1000 -2529 1000
rect -2463 -1000 -2433 1000
rect -2367 -1000 -2337 1000
rect -2271 -1000 -2241 1000
rect -2175 -1000 -2145 1000
rect -2079 -1000 -2049 1000
rect -1983 -1000 -1953 1000
rect -1887 -1000 -1857 1000
rect -1791 -1000 -1761 1000
rect -1695 -1000 -1665 1000
rect -1599 -1000 -1569 1000
rect -1503 -1000 -1473 1000
rect -1407 -1000 -1377 1000
rect -1311 -1000 -1281 1000
rect -1215 -1000 -1185 1000
rect -1119 -1000 -1089 1000
rect -1023 -1000 -993 1000
rect -927 -1000 -897 1000
rect -831 -1000 -801 1000
rect -735 -1000 -705 1000
rect -639 -1000 -609 1000
rect -543 -1000 -513 1000
rect -447 -1000 -417 1000
rect -351 -1000 -321 1000
rect -255 -1000 -225 1000
rect -159 -1000 -129 1000
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
rect 129 -1000 159 1000
rect 225 -1000 255 1000
rect 321 -1000 351 1000
rect 417 -1000 447 1000
rect 513 -1000 543 1000
rect 609 -1000 639 1000
rect 705 -1000 735 1000
rect 801 -1000 831 1000
rect 897 -1000 927 1000
rect 993 -1000 1023 1000
rect 1089 -1000 1119 1000
rect 1185 -1000 1215 1000
rect 1281 -1000 1311 1000
rect 1377 -1000 1407 1000
rect 1473 -1000 1503 1000
rect 1569 -1000 1599 1000
rect 1665 -1000 1695 1000
rect 1761 -1000 1791 1000
rect 1857 -1000 1887 1000
rect 1953 -1000 1983 1000
rect 2049 -1000 2079 1000
rect 2145 -1000 2175 1000
rect 2241 -1000 2271 1000
rect 2337 -1000 2367 1000
rect 2433 -1000 2463 1000
rect 2529 -1000 2559 1000
rect 2625 -1000 2655 1000
rect 2721 -1000 2751 1000
rect 2817 -1000 2847 1000
rect 2913 -1000 2943 1000
rect 3009 -1000 3039 1000
rect 3105 -1000 3135 1000
rect 3201 -1000 3231 1000
rect 3297 -1000 3327 1000
rect 3393 -1000 3423 1000
rect 3489 -1000 3519 1000
rect 3585 -1000 3615 1000
rect 3681 -1000 3711 1000
rect 3777 -1000 3807 1000
rect 3873 -1000 3903 1000
rect 3969 -1000 3999 1000
rect 4065 -1000 4095 1000
rect 4161 -1000 4191 1000
rect 4257 -1000 4287 1000
rect 4353 -1000 4383 1000
rect 4449 -1000 4479 1000
rect 4545 -1000 4575 1000
rect 4641 -1000 4671 1000
rect 4737 -1000 4767 1000
<< ndiff >>
rect -4829 969 -4767 1000
rect -4829 935 -4817 969
rect -4783 935 -4767 969
rect -4829 901 -4767 935
rect -4829 867 -4817 901
rect -4783 867 -4767 901
rect -4829 833 -4767 867
rect -4829 799 -4817 833
rect -4783 799 -4767 833
rect -4829 765 -4767 799
rect -4829 731 -4817 765
rect -4783 731 -4767 765
rect -4829 697 -4767 731
rect -4829 663 -4817 697
rect -4783 663 -4767 697
rect -4829 629 -4767 663
rect -4829 595 -4817 629
rect -4783 595 -4767 629
rect -4829 561 -4767 595
rect -4829 527 -4817 561
rect -4783 527 -4767 561
rect -4829 493 -4767 527
rect -4829 459 -4817 493
rect -4783 459 -4767 493
rect -4829 425 -4767 459
rect -4829 391 -4817 425
rect -4783 391 -4767 425
rect -4829 357 -4767 391
rect -4829 323 -4817 357
rect -4783 323 -4767 357
rect -4829 289 -4767 323
rect -4829 255 -4817 289
rect -4783 255 -4767 289
rect -4829 221 -4767 255
rect -4829 187 -4817 221
rect -4783 187 -4767 221
rect -4829 153 -4767 187
rect -4829 119 -4817 153
rect -4783 119 -4767 153
rect -4829 85 -4767 119
rect -4829 51 -4817 85
rect -4783 51 -4767 85
rect -4829 17 -4767 51
rect -4829 -17 -4817 17
rect -4783 -17 -4767 17
rect -4829 -51 -4767 -17
rect -4829 -85 -4817 -51
rect -4783 -85 -4767 -51
rect -4829 -119 -4767 -85
rect -4829 -153 -4817 -119
rect -4783 -153 -4767 -119
rect -4829 -187 -4767 -153
rect -4829 -221 -4817 -187
rect -4783 -221 -4767 -187
rect -4829 -255 -4767 -221
rect -4829 -289 -4817 -255
rect -4783 -289 -4767 -255
rect -4829 -323 -4767 -289
rect -4829 -357 -4817 -323
rect -4783 -357 -4767 -323
rect -4829 -391 -4767 -357
rect -4829 -425 -4817 -391
rect -4783 -425 -4767 -391
rect -4829 -459 -4767 -425
rect -4829 -493 -4817 -459
rect -4783 -493 -4767 -459
rect -4829 -527 -4767 -493
rect -4829 -561 -4817 -527
rect -4783 -561 -4767 -527
rect -4829 -595 -4767 -561
rect -4829 -629 -4817 -595
rect -4783 -629 -4767 -595
rect -4829 -663 -4767 -629
rect -4829 -697 -4817 -663
rect -4783 -697 -4767 -663
rect -4829 -731 -4767 -697
rect -4829 -765 -4817 -731
rect -4783 -765 -4767 -731
rect -4829 -799 -4767 -765
rect -4829 -833 -4817 -799
rect -4783 -833 -4767 -799
rect -4829 -867 -4767 -833
rect -4829 -901 -4817 -867
rect -4783 -901 -4767 -867
rect -4829 -935 -4767 -901
rect -4829 -969 -4817 -935
rect -4783 -969 -4767 -935
rect -4829 -1000 -4767 -969
rect -4737 969 -4671 1000
rect -4737 935 -4721 969
rect -4687 935 -4671 969
rect -4737 901 -4671 935
rect -4737 867 -4721 901
rect -4687 867 -4671 901
rect -4737 833 -4671 867
rect -4737 799 -4721 833
rect -4687 799 -4671 833
rect -4737 765 -4671 799
rect -4737 731 -4721 765
rect -4687 731 -4671 765
rect -4737 697 -4671 731
rect -4737 663 -4721 697
rect -4687 663 -4671 697
rect -4737 629 -4671 663
rect -4737 595 -4721 629
rect -4687 595 -4671 629
rect -4737 561 -4671 595
rect -4737 527 -4721 561
rect -4687 527 -4671 561
rect -4737 493 -4671 527
rect -4737 459 -4721 493
rect -4687 459 -4671 493
rect -4737 425 -4671 459
rect -4737 391 -4721 425
rect -4687 391 -4671 425
rect -4737 357 -4671 391
rect -4737 323 -4721 357
rect -4687 323 -4671 357
rect -4737 289 -4671 323
rect -4737 255 -4721 289
rect -4687 255 -4671 289
rect -4737 221 -4671 255
rect -4737 187 -4721 221
rect -4687 187 -4671 221
rect -4737 153 -4671 187
rect -4737 119 -4721 153
rect -4687 119 -4671 153
rect -4737 85 -4671 119
rect -4737 51 -4721 85
rect -4687 51 -4671 85
rect -4737 17 -4671 51
rect -4737 -17 -4721 17
rect -4687 -17 -4671 17
rect -4737 -51 -4671 -17
rect -4737 -85 -4721 -51
rect -4687 -85 -4671 -51
rect -4737 -119 -4671 -85
rect -4737 -153 -4721 -119
rect -4687 -153 -4671 -119
rect -4737 -187 -4671 -153
rect -4737 -221 -4721 -187
rect -4687 -221 -4671 -187
rect -4737 -255 -4671 -221
rect -4737 -289 -4721 -255
rect -4687 -289 -4671 -255
rect -4737 -323 -4671 -289
rect -4737 -357 -4721 -323
rect -4687 -357 -4671 -323
rect -4737 -391 -4671 -357
rect -4737 -425 -4721 -391
rect -4687 -425 -4671 -391
rect -4737 -459 -4671 -425
rect -4737 -493 -4721 -459
rect -4687 -493 -4671 -459
rect -4737 -527 -4671 -493
rect -4737 -561 -4721 -527
rect -4687 -561 -4671 -527
rect -4737 -595 -4671 -561
rect -4737 -629 -4721 -595
rect -4687 -629 -4671 -595
rect -4737 -663 -4671 -629
rect -4737 -697 -4721 -663
rect -4687 -697 -4671 -663
rect -4737 -731 -4671 -697
rect -4737 -765 -4721 -731
rect -4687 -765 -4671 -731
rect -4737 -799 -4671 -765
rect -4737 -833 -4721 -799
rect -4687 -833 -4671 -799
rect -4737 -867 -4671 -833
rect -4737 -901 -4721 -867
rect -4687 -901 -4671 -867
rect -4737 -935 -4671 -901
rect -4737 -969 -4721 -935
rect -4687 -969 -4671 -935
rect -4737 -1000 -4671 -969
rect -4641 969 -4575 1000
rect -4641 935 -4625 969
rect -4591 935 -4575 969
rect -4641 901 -4575 935
rect -4641 867 -4625 901
rect -4591 867 -4575 901
rect -4641 833 -4575 867
rect -4641 799 -4625 833
rect -4591 799 -4575 833
rect -4641 765 -4575 799
rect -4641 731 -4625 765
rect -4591 731 -4575 765
rect -4641 697 -4575 731
rect -4641 663 -4625 697
rect -4591 663 -4575 697
rect -4641 629 -4575 663
rect -4641 595 -4625 629
rect -4591 595 -4575 629
rect -4641 561 -4575 595
rect -4641 527 -4625 561
rect -4591 527 -4575 561
rect -4641 493 -4575 527
rect -4641 459 -4625 493
rect -4591 459 -4575 493
rect -4641 425 -4575 459
rect -4641 391 -4625 425
rect -4591 391 -4575 425
rect -4641 357 -4575 391
rect -4641 323 -4625 357
rect -4591 323 -4575 357
rect -4641 289 -4575 323
rect -4641 255 -4625 289
rect -4591 255 -4575 289
rect -4641 221 -4575 255
rect -4641 187 -4625 221
rect -4591 187 -4575 221
rect -4641 153 -4575 187
rect -4641 119 -4625 153
rect -4591 119 -4575 153
rect -4641 85 -4575 119
rect -4641 51 -4625 85
rect -4591 51 -4575 85
rect -4641 17 -4575 51
rect -4641 -17 -4625 17
rect -4591 -17 -4575 17
rect -4641 -51 -4575 -17
rect -4641 -85 -4625 -51
rect -4591 -85 -4575 -51
rect -4641 -119 -4575 -85
rect -4641 -153 -4625 -119
rect -4591 -153 -4575 -119
rect -4641 -187 -4575 -153
rect -4641 -221 -4625 -187
rect -4591 -221 -4575 -187
rect -4641 -255 -4575 -221
rect -4641 -289 -4625 -255
rect -4591 -289 -4575 -255
rect -4641 -323 -4575 -289
rect -4641 -357 -4625 -323
rect -4591 -357 -4575 -323
rect -4641 -391 -4575 -357
rect -4641 -425 -4625 -391
rect -4591 -425 -4575 -391
rect -4641 -459 -4575 -425
rect -4641 -493 -4625 -459
rect -4591 -493 -4575 -459
rect -4641 -527 -4575 -493
rect -4641 -561 -4625 -527
rect -4591 -561 -4575 -527
rect -4641 -595 -4575 -561
rect -4641 -629 -4625 -595
rect -4591 -629 -4575 -595
rect -4641 -663 -4575 -629
rect -4641 -697 -4625 -663
rect -4591 -697 -4575 -663
rect -4641 -731 -4575 -697
rect -4641 -765 -4625 -731
rect -4591 -765 -4575 -731
rect -4641 -799 -4575 -765
rect -4641 -833 -4625 -799
rect -4591 -833 -4575 -799
rect -4641 -867 -4575 -833
rect -4641 -901 -4625 -867
rect -4591 -901 -4575 -867
rect -4641 -935 -4575 -901
rect -4641 -969 -4625 -935
rect -4591 -969 -4575 -935
rect -4641 -1000 -4575 -969
rect -4545 969 -4479 1000
rect -4545 935 -4529 969
rect -4495 935 -4479 969
rect -4545 901 -4479 935
rect -4545 867 -4529 901
rect -4495 867 -4479 901
rect -4545 833 -4479 867
rect -4545 799 -4529 833
rect -4495 799 -4479 833
rect -4545 765 -4479 799
rect -4545 731 -4529 765
rect -4495 731 -4479 765
rect -4545 697 -4479 731
rect -4545 663 -4529 697
rect -4495 663 -4479 697
rect -4545 629 -4479 663
rect -4545 595 -4529 629
rect -4495 595 -4479 629
rect -4545 561 -4479 595
rect -4545 527 -4529 561
rect -4495 527 -4479 561
rect -4545 493 -4479 527
rect -4545 459 -4529 493
rect -4495 459 -4479 493
rect -4545 425 -4479 459
rect -4545 391 -4529 425
rect -4495 391 -4479 425
rect -4545 357 -4479 391
rect -4545 323 -4529 357
rect -4495 323 -4479 357
rect -4545 289 -4479 323
rect -4545 255 -4529 289
rect -4495 255 -4479 289
rect -4545 221 -4479 255
rect -4545 187 -4529 221
rect -4495 187 -4479 221
rect -4545 153 -4479 187
rect -4545 119 -4529 153
rect -4495 119 -4479 153
rect -4545 85 -4479 119
rect -4545 51 -4529 85
rect -4495 51 -4479 85
rect -4545 17 -4479 51
rect -4545 -17 -4529 17
rect -4495 -17 -4479 17
rect -4545 -51 -4479 -17
rect -4545 -85 -4529 -51
rect -4495 -85 -4479 -51
rect -4545 -119 -4479 -85
rect -4545 -153 -4529 -119
rect -4495 -153 -4479 -119
rect -4545 -187 -4479 -153
rect -4545 -221 -4529 -187
rect -4495 -221 -4479 -187
rect -4545 -255 -4479 -221
rect -4545 -289 -4529 -255
rect -4495 -289 -4479 -255
rect -4545 -323 -4479 -289
rect -4545 -357 -4529 -323
rect -4495 -357 -4479 -323
rect -4545 -391 -4479 -357
rect -4545 -425 -4529 -391
rect -4495 -425 -4479 -391
rect -4545 -459 -4479 -425
rect -4545 -493 -4529 -459
rect -4495 -493 -4479 -459
rect -4545 -527 -4479 -493
rect -4545 -561 -4529 -527
rect -4495 -561 -4479 -527
rect -4545 -595 -4479 -561
rect -4545 -629 -4529 -595
rect -4495 -629 -4479 -595
rect -4545 -663 -4479 -629
rect -4545 -697 -4529 -663
rect -4495 -697 -4479 -663
rect -4545 -731 -4479 -697
rect -4545 -765 -4529 -731
rect -4495 -765 -4479 -731
rect -4545 -799 -4479 -765
rect -4545 -833 -4529 -799
rect -4495 -833 -4479 -799
rect -4545 -867 -4479 -833
rect -4545 -901 -4529 -867
rect -4495 -901 -4479 -867
rect -4545 -935 -4479 -901
rect -4545 -969 -4529 -935
rect -4495 -969 -4479 -935
rect -4545 -1000 -4479 -969
rect -4449 969 -4383 1000
rect -4449 935 -4433 969
rect -4399 935 -4383 969
rect -4449 901 -4383 935
rect -4449 867 -4433 901
rect -4399 867 -4383 901
rect -4449 833 -4383 867
rect -4449 799 -4433 833
rect -4399 799 -4383 833
rect -4449 765 -4383 799
rect -4449 731 -4433 765
rect -4399 731 -4383 765
rect -4449 697 -4383 731
rect -4449 663 -4433 697
rect -4399 663 -4383 697
rect -4449 629 -4383 663
rect -4449 595 -4433 629
rect -4399 595 -4383 629
rect -4449 561 -4383 595
rect -4449 527 -4433 561
rect -4399 527 -4383 561
rect -4449 493 -4383 527
rect -4449 459 -4433 493
rect -4399 459 -4383 493
rect -4449 425 -4383 459
rect -4449 391 -4433 425
rect -4399 391 -4383 425
rect -4449 357 -4383 391
rect -4449 323 -4433 357
rect -4399 323 -4383 357
rect -4449 289 -4383 323
rect -4449 255 -4433 289
rect -4399 255 -4383 289
rect -4449 221 -4383 255
rect -4449 187 -4433 221
rect -4399 187 -4383 221
rect -4449 153 -4383 187
rect -4449 119 -4433 153
rect -4399 119 -4383 153
rect -4449 85 -4383 119
rect -4449 51 -4433 85
rect -4399 51 -4383 85
rect -4449 17 -4383 51
rect -4449 -17 -4433 17
rect -4399 -17 -4383 17
rect -4449 -51 -4383 -17
rect -4449 -85 -4433 -51
rect -4399 -85 -4383 -51
rect -4449 -119 -4383 -85
rect -4449 -153 -4433 -119
rect -4399 -153 -4383 -119
rect -4449 -187 -4383 -153
rect -4449 -221 -4433 -187
rect -4399 -221 -4383 -187
rect -4449 -255 -4383 -221
rect -4449 -289 -4433 -255
rect -4399 -289 -4383 -255
rect -4449 -323 -4383 -289
rect -4449 -357 -4433 -323
rect -4399 -357 -4383 -323
rect -4449 -391 -4383 -357
rect -4449 -425 -4433 -391
rect -4399 -425 -4383 -391
rect -4449 -459 -4383 -425
rect -4449 -493 -4433 -459
rect -4399 -493 -4383 -459
rect -4449 -527 -4383 -493
rect -4449 -561 -4433 -527
rect -4399 -561 -4383 -527
rect -4449 -595 -4383 -561
rect -4449 -629 -4433 -595
rect -4399 -629 -4383 -595
rect -4449 -663 -4383 -629
rect -4449 -697 -4433 -663
rect -4399 -697 -4383 -663
rect -4449 -731 -4383 -697
rect -4449 -765 -4433 -731
rect -4399 -765 -4383 -731
rect -4449 -799 -4383 -765
rect -4449 -833 -4433 -799
rect -4399 -833 -4383 -799
rect -4449 -867 -4383 -833
rect -4449 -901 -4433 -867
rect -4399 -901 -4383 -867
rect -4449 -935 -4383 -901
rect -4449 -969 -4433 -935
rect -4399 -969 -4383 -935
rect -4449 -1000 -4383 -969
rect -4353 969 -4287 1000
rect -4353 935 -4337 969
rect -4303 935 -4287 969
rect -4353 901 -4287 935
rect -4353 867 -4337 901
rect -4303 867 -4287 901
rect -4353 833 -4287 867
rect -4353 799 -4337 833
rect -4303 799 -4287 833
rect -4353 765 -4287 799
rect -4353 731 -4337 765
rect -4303 731 -4287 765
rect -4353 697 -4287 731
rect -4353 663 -4337 697
rect -4303 663 -4287 697
rect -4353 629 -4287 663
rect -4353 595 -4337 629
rect -4303 595 -4287 629
rect -4353 561 -4287 595
rect -4353 527 -4337 561
rect -4303 527 -4287 561
rect -4353 493 -4287 527
rect -4353 459 -4337 493
rect -4303 459 -4287 493
rect -4353 425 -4287 459
rect -4353 391 -4337 425
rect -4303 391 -4287 425
rect -4353 357 -4287 391
rect -4353 323 -4337 357
rect -4303 323 -4287 357
rect -4353 289 -4287 323
rect -4353 255 -4337 289
rect -4303 255 -4287 289
rect -4353 221 -4287 255
rect -4353 187 -4337 221
rect -4303 187 -4287 221
rect -4353 153 -4287 187
rect -4353 119 -4337 153
rect -4303 119 -4287 153
rect -4353 85 -4287 119
rect -4353 51 -4337 85
rect -4303 51 -4287 85
rect -4353 17 -4287 51
rect -4353 -17 -4337 17
rect -4303 -17 -4287 17
rect -4353 -51 -4287 -17
rect -4353 -85 -4337 -51
rect -4303 -85 -4287 -51
rect -4353 -119 -4287 -85
rect -4353 -153 -4337 -119
rect -4303 -153 -4287 -119
rect -4353 -187 -4287 -153
rect -4353 -221 -4337 -187
rect -4303 -221 -4287 -187
rect -4353 -255 -4287 -221
rect -4353 -289 -4337 -255
rect -4303 -289 -4287 -255
rect -4353 -323 -4287 -289
rect -4353 -357 -4337 -323
rect -4303 -357 -4287 -323
rect -4353 -391 -4287 -357
rect -4353 -425 -4337 -391
rect -4303 -425 -4287 -391
rect -4353 -459 -4287 -425
rect -4353 -493 -4337 -459
rect -4303 -493 -4287 -459
rect -4353 -527 -4287 -493
rect -4353 -561 -4337 -527
rect -4303 -561 -4287 -527
rect -4353 -595 -4287 -561
rect -4353 -629 -4337 -595
rect -4303 -629 -4287 -595
rect -4353 -663 -4287 -629
rect -4353 -697 -4337 -663
rect -4303 -697 -4287 -663
rect -4353 -731 -4287 -697
rect -4353 -765 -4337 -731
rect -4303 -765 -4287 -731
rect -4353 -799 -4287 -765
rect -4353 -833 -4337 -799
rect -4303 -833 -4287 -799
rect -4353 -867 -4287 -833
rect -4353 -901 -4337 -867
rect -4303 -901 -4287 -867
rect -4353 -935 -4287 -901
rect -4353 -969 -4337 -935
rect -4303 -969 -4287 -935
rect -4353 -1000 -4287 -969
rect -4257 969 -4191 1000
rect -4257 935 -4241 969
rect -4207 935 -4191 969
rect -4257 901 -4191 935
rect -4257 867 -4241 901
rect -4207 867 -4191 901
rect -4257 833 -4191 867
rect -4257 799 -4241 833
rect -4207 799 -4191 833
rect -4257 765 -4191 799
rect -4257 731 -4241 765
rect -4207 731 -4191 765
rect -4257 697 -4191 731
rect -4257 663 -4241 697
rect -4207 663 -4191 697
rect -4257 629 -4191 663
rect -4257 595 -4241 629
rect -4207 595 -4191 629
rect -4257 561 -4191 595
rect -4257 527 -4241 561
rect -4207 527 -4191 561
rect -4257 493 -4191 527
rect -4257 459 -4241 493
rect -4207 459 -4191 493
rect -4257 425 -4191 459
rect -4257 391 -4241 425
rect -4207 391 -4191 425
rect -4257 357 -4191 391
rect -4257 323 -4241 357
rect -4207 323 -4191 357
rect -4257 289 -4191 323
rect -4257 255 -4241 289
rect -4207 255 -4191 289
rect -4257 221 -4191 255
rect -4257 187 -4241 221
rect -4207 187 -4191 221
rect -4257 153 -4191 187
rect -4257 119 -4241 153
rect -4207 119 -4191 153
rect -4257 85 -4191 119
rect -4257 51 -4241 85
rect -4207 51 -4191 85
rect -4257 17 -4191 51
rect -4257 -17 -4241 17
rect -4207 -17 -4191 17
rect -4257 -51 -4191 -17
rect -4257 -85 -4241 -51
rect -4207 -85 -4191 -51
rect -4257 -119 -4191 -85
rect -4257 -153 -4241 -119
rect -4207 -153 -4191 -119
rect -4257 -187 -4191 -153
rect -4257 -221 -4241 -187
rect -4207 -221 -4191 -187
rect -4257 -255 -4191 -221
rect -4257 -289 -4241 -255
rect -4207 -289 -4191 -255
rect -4257 -323 -4191 -289
rect -4257 -357 -4241 -323
rect -4207 -357 -4191 -323
rect -4257 -391 -4191 -357
rect -4257 -425 -4241 -391
rect -4207 -425 -4191 -391
rect -4257 -459 -4191 -425
rect -4257 -493 -4241 -459
rect -4207 -493 -4191 -459
rect -4257 -527 -4191 -493
rect -4257 -561 -4241 -527
rect -4207 -561 -4191 -527
rect -4257 -595 -4191 -561
rect -4257 -629 -4241 -595
rect -4207 -629 -4191 -595
rect -4257 -663 -4191 -629
rect -4257 -697 -4241 -663
rect -4207 -697 -4191 -663
rect -4257 -731 -4191 -697
rect -4257 -765 -4241 -731
rect -4207 -765 -4191 -731
rect -4257 -799 -4191 -765
rect -4257 -833 -4241 -799
rect -4207 -833 -4191 -799
rect -4257 -867 -4191 -833
rect -4257 -901 -4241 -867
rect -4207 -901 -4191 -867
rect -4257 -935 -4191 -901
rect -4257 -969 -4241 -935
rect -4207 -969 -4191 -935
rect -4257 -1000 -4191 -969
rect -4161 969 -4095 1000
rect -4161 935 -4145 969
rect -4111 935 -4095 969
rect -4161 901 -4095 935
rect -4161 867 -4145 901
rect -4111 867 -4095 901
rect -4161 833 -4095 867
rect -4161 799 -4145 833
rect -4111 799 -4095 833
rect -4161 765 -4095 799
rect -4161 731 -4145 765
rect -4111 731 -4095 765
rect -4161 697 -4095 731
rect -4161 663 -4145 697
rect -4111 663 -4095 697
rect -4161 629 -4095 663
rect -4161 595 -4145 629
rect -4111 595 -4095 629
rect -4161 561 -4095 595
rect -4161 527 -4145 561
rect -4111 527 -4095 561
rect -4161 493 -4095 527
rect -4161 459 -4145 493
rect -4111 459 -4095 493
rect -4161 425 -4095 459
rect -4161 391 -4145 425
rect -4111 391 -4095 425
rect -4161 357 -4095 391
rect -4161 323 -4145 357
rect -4111 323 -4095 357
rect -4161 289 -4095 323
rect -4161 255 -4145 289
rect -4111 255 -4095 289
rect -4161 221 -4095 255
rect -4161 187 -4145 221
rect -4111 187 -4095 221
rect -4161 153 -4095 187
rect -4161 119 -4145 153
rect -4111 119 -4095 153
rect -4161 85 -4095 119
rect -4161 51 -4145 85
rect -4111 51 -4095 85
rect -4161 17 -4095 51
rect -4161 -17 -4145 17
rect -4111 -17 -4095 17
rect -4161 -51 -4095 -17
rect -4161 -85 -4145 -51
rect -4111 -85 -4095 -51
rect -4161 -119 -4095 -85
rect -4161 -153 -4145 -119
rect -4111 -153 -4095 -119
rect -4161 -187 -4095 -153
rect -4161 -221 -4145 -187
rect -4111 -221 -4095 -187
rect -4161 -255 -4095 -221
rect -4161 -289 -4145 -255
rect -4111 -289 -4095 -255
rect -4161 -323 -4095 -289
rect -4161 -357 -4145 -323
rect -4111 -357 -4095 -323
rect -4161 -391 -4095 -357
rect -4161 -425 -4145 -391
rect -4111 -425 -4095 -391
rect -4161 -459 -4095 -425
rect -4161 -493 -4145 -459
rect -4111 -493 -4095 -459
rect -4161 -527 -4095 -493
rect -4161 -561 -4145 -527
rect -4111 -561 -4095 -527
rect -4161 -595 -4095 -561
rect -4161 -629 -4145 -595
rect -4111 -629 -4095 -595
rect -4161 -663 -4095 -629
rect -4161 -697 -4145 -663
rect -4111 -697 -4095 -663
rect -4161 -731 -4095 -697
rect -4161 -765 -4145 -731
rect -4111 -765 -4095 -731
rect -4161 -799 -4095 -765
rect -4161 -833 -4145 -799
rect -4111 -833 -4095 -799
rect -4161 -867 -4095 -833
rect -4161 -901 -4145 -867
rect -4111 -901 -4095 -867
rect -4161 -935 -4095 -901
rect -4161 -969 -4145 -935
rect -4111 -969 -4095 -935
rect -4161 -1000 -4095 -969
rect -4065 969 -3999 1000
rect -4065 935 -4049 969
rect -4015 935 -3999 969
rect -4065 901 -3999 935
rect -4065 867 -4049 901
rect -4015 867 -3999 901
rect -4065 833 -3999 867
rect -4065 799 -4049 833
rect -4015 799 -3999 833
rect -4065 765 -3999 799
rect -4065 731 -4049 765
rect -4015 731 -3999 765
rect -4065 697 -3999 731
rect -4065 663 -4049 697
rect -4015 663 -3999 697
rect -4065 629 -3999 663
rect -4065 595 -4049 629
rect -4015 595 -3999 629
rect -4065 561 -3999 595
rect -4065 527 -4049 561
rect -4015 527 -3999 561
rect -4065 493 -3999 527
rect -4065 459 -4049 493
rect -4015 459 -3999 493
rect -4065 425 -3999 459
rect -4065 391 -4049 425
rect -4015 391 -3999 425
rect -4065 357 -3999 391
rect -4065 323 -4049 357
rect -4015 323 -3999 357
rect -4065 289 -3999 323
rect -4065 255 -4049 289
rect -4015 255 -3999 289
rect -4065 221 -3999 255
rect -4065 187 -4049 221
rect -4015 187 -3999 221
rect -4065 153 -3999 187
rect -4065 119 -4049 153
rect -4015 119 -3999 153
rect -4065 85 -3999 119
rect -4065 51 -4049 85
rect -4015 51 -3999 85
rect -4065 17 -3999 51
rect -4065 -17 -4049 17
rect -4015 -17 -3999 17
rect -4065 -51 -3999 -17
rect -4065 -85 -4049 -51
rect -4015 -85 -3999 -51
rect -4065 -119 -3999 -85
rect -4065 -153 -4049 -119
rect -4015 -153 -3999 -119
rect -4065 -187 -3999 -153
rect -4065 -221 -4049 -187
rect -4015 -221 -3999 -187
rect -4065 -255 -3999 -221
rect -4065 -289 -4049 -255
rect -4015 -289 -3999 -255
rect -4065 -323 -3999 -289
rect -4065 -357 -4049 -323
rect -4015 -357 -3999 -323
rect -4065 -391 -3999 -357
rect -4065 -425 -4049 -391
rect -4015 -425 -3999 -391
rect -4065 -459 -3999 -425
rect -4065 -493 -4049 -459
rect -4015 -493 -3999 -459
rect -4065 -527 -3999 -493
rect -4065 -561 -4049 -527
rect -4015 -561 -3999 -527
rect -4065 -595 -3999 -561
rect -4065 -629 -4049 -595
rect -4015 -629 -3999 -595
rect -4065 -663 -3999 -629
rect -4065 -697 -4049 -663
rect -4015 -697 -3999 -663
rect -4065 -731 -3999 -697
rect -4065 -765 -4049 -731
rect -4015 -765 -3999 -731
rect -4065 -799 -3999 -765
rect -4065 -833 -4049 -799
rect -4015 -833 -3999 -799
rect -4065 -867 -3999 -833
rect -4065 -901 -4049 -867
rect -4015 -901 -3999 -867
rect -4065 -935 -3999 -901
rect -4065 -969 -4049 -935
rect -4015 -969 -3999 -935
rect -4065 -1000 -3999 -969
rect -3969 969 -3903 1000
rect -3969 935 -3953 969
rect -3919 935 -3903 969
rect -3969 901 -3903 935
rect -3969 867 -3953 901
rect -3919 867 -3903 901
rect -3969 833 -3903 867
rect -3969 799 -3953 833
rect -3919 799 -3903 833
rect -3969 765 -3903 799
rect -3969 731 -3953 765
rect -3919 731 -3903 765
rect -3969 697 -3903 731
rect -3969 663 -3953 697
rect -3919 663 -3903 697
rect -3969 629 -3903 663
rect -3969 595 -3953 629
rect -3919 595 -3903 629
rect -3969 561 -3903 595
rect -3969 527 -3953 561
rect -3919 527 -3903 561
rect -3969 493 -3903 527
rect -3969 459 -3953 493
rect -3919 459 -3903 493
rect -3969 425 -3903 459
rect -3969 391 -3953 425
rect -3919 391 -3903 425
rect -3969 357 -3903 391
rect -3969 323 -3953 357
rect -3919 323 -3903 357
rect -3969 289 -3903 323
rect -3969 255 -3953 289
rect -3919 255 -3903 289
rect -3969 221 -3903 255
rect -3969 187 -3953 221
rect -3919 187 -3903 221
rect -3969 153 -3903 187
rect -3969 119 -3953 153
rect -3919 119 -3903 153
rect -3969 85 -3903 119
rect -3969 51 -3953 85
rect -3919 51 -3903 85
rect -3969 17 -3903 51
rect -3969 -17 -3953 17
rect -3919 -17 -3903 17
rect -3969 -51 -3903 -17
rect -3969 -85 -3953 -51
rect -3919 -85 -3903 -51
rect -3969 -119 -3903 -85
rect -3969 -153 -3953 -119
rect -3919 -153 -3903 -119
rect -3969 -187 -3903 -153
rect -3969 -221 -3953 -187
rect -3919 -221 -3903 -187
rect -3969 -255 -3903 -221
rect -3969 -289 -3953 -255
rect -3919 -289 -3903 -255
rect -3969 -323 -3903 -289
rect -3969 -357 -3953 -323
rect -3919 -357 -3903 -323
rect -3969 -391 -3903 -357
rect -3969 -425 -3953 -391
rect -3919 -425 -3903 -391
rect -3969 -459 -3903 -425
rect -3969 -493 -3953 -459
rect -3919 -493 -3903 -459
rect -3969 -527 -3903 -493
rect -3969 -561 -3953 -527
rect -3919 -561 -3903 -527
rect -3969 -595 -3903 -561
rect -3969 -629 -3953 -595
rect -3919 -629 -3903 -595
rect -3969 -663 -3903 -629
rect -3969 -697 -3953 -663
rect -3919 -697 -3903 -663
rect -3969 -731 -3903 -697
rect -3969 -765 -3953 -731
rect -3919 -765 -3903 -731
rect -3969 -799 -3903 -765
rect -3969 -833 -3953 -799
rect -3919 -833 -3903 -799
rect -3969 -867 -3903 -833
rect -3969 -901 -3953 -867
rect -3919 -901 -3903 -867
rect -3969 -935 -3903 -901
rect -3969 -969 -3953 -935
rect -3919 -969 -3903 -935
rect -3969 -1000 -3903 -969
rect -3873 969 -3807 1000
rect -3873 935 -3857 969
rect -3823 935 -3807 969
rect -3873 901 -3807 935
rect -3873 867 -3857 901
rect -3823 867 -3807 901
rect -3873 833 -3807 867
rect -3873 799 -3857 833
rect -3823 799 -3807 833
rect -3873 765 -3807 799
rect -3873 731 -3857 765
rect -3823 731 -3807 765
rect -3873 697 -3807 731
rect -3873 663 -3857 697
rect -3823 663 -3807 697
rect -3873 629 -3807 663
rect -3873 595 -3857 629
rect -3823 595 -3807 629
rect -3873 561 -3807 595
rect -3873 527 -3857 561
rect -3823 527 -3807 561
rect -3873 493 -3807 527
rect -3873 459 -3857 493
rect -3823 459 -3807 493
rect -3873 425 -3807 459
rect -3873 391 -3857 425
rect -3823 391 -3807 425
rect -3873 357 -3807 391
rect -3873 323 -3857 357
rect -3823 323 -3807 357
rect -3873 289 -3807 323
rect -3873 255 -3857 289
rect -3823 255 -3807 289
rect -3873 221 -3807 255
rect -3873 187 -3857 221
rect -3823 187 -3807 221
rect -3873 153 -3807 187
rect -3873 119 -3857 153
rect -3823 119 -3807 153
rect -3873 85 -3807 119
rect -3873 51 -3857 85
rect -3823 51 -3807 85
rect -3873 17 -3807 51
rect -3873 -17 -3857 17
rect -3823 -17 -3807 17
rect -3873 -51 -3807 -17
rect -3873 -85 -3857 -51
rect -3823 -85 -3807 -51
rect -3873 -119 -3807 -85
rect -3873 -153 -3857 -119
rect -3823 -153 -3807 -119
rect -3873 -187 -3807 -153
rect -3873 -221 -3857 -187
rect -3823 -221 -3807 -187
rect -3873 -255 -3807 -221
rect -3873 -289 -3857 -255
rect -3823 -289 -3807 -255
rect -3873 -323 -3807 -289
rect -3873 -357 -3857 -323
rect -3823 -357 -3807 -323
rect -3873 -391 -3807 -357
rect -3873 -425 -3857 -391
rect -3823 -425 -3807 -391
rect -3873 -459 -3807 -425
rect -3873 -493 -3857 -459
rect -3823 -493 -3807 -459
rect -3873 -527 -3807 -493
rect -3873 -561 -3857 -527
rect -3823 -561 -3807 -527
rect -3873 -595 -3807 -561
rect -3873 -629 -3857 -595
rect -3823 -629 -3807 -595
rect -3873 -663 -3807 -629
rect -3873 -697 -3857 -663
rect -3823 -697 -3807 -663
rect -3873 -731 -3807 -697
rect -3873 -765 -3857 -731
rect -3823 -765 -3807 -731
rect -3873 -799 -3807 -765
rect -3873 -833 -3857 -799
rect -3823 -833 -3807 -799
rect -3873 -867 -3807 -833
rect -3873 -901 -3857 -867
rect -3823 -901 -3807 -867
rect -3873 -935 -3807 -901
rect -3873 -969 -3857 -935
rect -3823 -969 -3807 -935
rect -3873 -1000 -3807 -969
rect -3777 969 -3711 1000
rect -3777 935 -3761 969
rect -3727 935 -3711 969
rect -3777 901 -3711 935
rect -3777 867 -3761 901
rect -3727 867 -3711 901
rect -3777 833 -3711 867
rect -3777 799 -3761 833
rect -3727 799 -3711 833
rect -3777 765 -3711 799
rect -3777 731 -3761 765
rect -3727 731 -3711 765
rect -3777 697 -3711 731
rect -3777 663 -3761 697
rect -3727 663 -3711 697
rect -3777 629 -3711 663
rect -3777 595 -3761 629
rect -3727 595 -3711 629
rect -3777 561 -3711 595
rect -3777 527 -3761 561
rect -3727 527 -3711 561
rect -3777 493 -3711 527
rect -3777 459 -3761 493
rect -3727 459 -3711 493
rect -3777 425 -3711 459
rect -3777 391 -3761 425
rect -3727 391 -3711 425
rect -3777 357 -3711 391
rect -3777 323 -3761 357
rect -3727 323 -3711 357
rect -3777 289 -3711 323
rect -3777 255 -3761 289
rect -3727 255 -3711 289
rect -3777 221 -3711 255
rect -3777 187 -3761 221
rect -3727 187 -3711 221
rect -3777 153 -3711 187
rect -3777 119 -3761 153
rect -3727 119 -3711 153
rect -3777 85 -3711 119
rect -3777 51 -3761 85
rect -3727 51 -3711 85
rect -3777 17 -3711 51
rect -3777 -17 -3761 17
rect -3727 -17 -3711 17
rect -3777 -51 -3711 -17
rect -3777 -85 -3761 -51
rect -3727 -85 -3711 -51
rect -3777 -119 -3711 -85
rect -3777 -153 -3761 -119
rect -3727 -153 -3711 -119
rect -3777 -187 -3711 -153
rect -3777 -221 -3761 -187
rect -3727 -221 -3711 -187
rect -3777 -255 -3711 -221
rect -3777 -289 -3761 -255
rect -3727 -289 -3711 -255
rect -3777 -323 -3711 -289
rect -3777 -357 -3761 -323
rect -3727 -357 -3711 -323
rect -3777 -391 -3711 -357
rect -3777 -425 -3761 -391
rect -3727 -425 -3711 -391
rect -3777 -459 -3711 -425
rect -3777 -493 -3761 -459
rect -3727 -493 -3711 -459
rect -3777 -527 -3711 -493
rect -3777 -561 -3761 -527
rect -3727 -561 -3711 -527
rect -3777 -595 -3711 -561
rect -3777 -629 -3761 -595
rect -3727 -629 -3711 -595
rect -3777 -663 -3711 -629
rect -3777 -697 -3761 -663
rect -3727 -697 -3711 -663
rect -3777 -731 -3711 -697
rect -3777 -765 -3761 -731
rect -3727 -765 -3711 -731
rect -3777 -799 -3711 -765
rect -3777 -833 -3761 -799
rect -3727 -833 -3711 -799
rect -3777 -867 -3711 -833
rect -3777 -901 -3761 -867
rect -3727 -901 -3711 -867
rect -3777 -935 -3711 -901
rect -3777 -969 -3761 -935
rect -3727 -969 -3711 -935
rect -3777 -1000 -3711 -969
rect -3681 969 -3615 1000
rect -3681 935 -3665 969
rect -3631 935 -3615 969
rect -3681 901 -3615 935
rect -3681 867 -3665 901
rect -3631 867 -3615 901
rect -3681 833 -3615 867
rect -3681 799 -3665 833
rect -3631 799 -3615 833
rect -3681 765 -3615 799
rect -3681 731 -3665 765
rect -3631 731 -3615 765
rect -3681 697 -3615 731
rect -3681 663 -3665 697
rect -3631 663 -3615 697
rect -3681 629 -3615 663
rect -3681 595 -3665 629
rect -3631 595 -3615 629
rect -3681 561 -3615 595
rect -3681 527 -3665 561
rect -3631 527 -3615 561
rect -3681 493 -3615 527
rect -3681 459 -3665 493
rect -3631 459 -3615 493
rect -3681 425 -3615 459
rect -3681 391 -3665 425
rect -3631 391 -3615 425
rect -3681 357 -3615 391
rect -3681 323 -3665 357
rect -3631 323 -3615 357
rect -3681 289 -3615 323
rect -3681 255 -3665 289
rect -3631 255 -3615 289
rect -3681 221 -3615 255
rect -3681 187 -3665 221
rect -3631 187 -3615 221
rect -3681 153 -3615 187
rect -3681 119 -3665 153
rect -3631 119 -3615 153
rect -3681 85 -3615 119
rect -3681 51 -3665 85
rect -3631 51 -3615 85
rect -3681 17 -3615 51
rect -3681 -17 -3665 17
rect -3631 -17 -3615 17
rect -3681 -51 -3615 -17
rect -3681 -85 -3665 -51
rect -3631 -85 -3615 -51
rect -3681 -119 -3615 -85
rect -3681 -153 -3665 -119
rect -3631 -153 -3615 -119
rect -3681 -187 -3615 -153
rect -3681 -221 -3665 -187
rect -3631 -221 -3615 -187
rect -3681 -255 -3615 -221
rect -3681 -289 -3665 -255
rect -3631 -289 -3615 -255
rect -3681 -323 -3615 -289
rect -3681 -357 -3665 -323
rect -3631 -357 -3615 -323
rect -3681 -391 -3615 -357
rect -3681 -425 -3665 -391
rect -3631 -425 -3615 -391
rect -3681 -459 -3615 -425
rect -3681 -493 -3665 -459
rect -3631 -493 -3615 -459
rect -3681 -527 -3615 -493
rect -3681 -561 -3665 -527
rect -3631 -561 -3615 -527
rect -3681 -595 -3615 -561
rect -3681 -629 -3665 -595
rect -3631 -629 -3615 -595
rect -3681 -663 -3615 -629
rect -3681 -697 -3665 -663
rect -3631 -697 -3615 -663
rect -3681 -731 -3615 -697
rect -3681 -765 -3665 -731
rect -3631 -765 -3615 -731
rect -3681 -799 -3615 -765
rect -3681 -833 -3665 -799
rect -3631 -833 -3615 -799
rect -3681 -867 -3615 -833
rect -3681 -901 -3665 -867
rect -3631 -901 -3615 -867
rect -3681 -935 -3615 -901
rect -3681 -969 -3665 -935
rect -3631 -969 -3615 -935
rect -3681 -1000 -3615 -969
rect -3585 969 -3519 1000
rect -3585 935 -3569 969
rect -3535 935 -3519 969
rect -3585 901 -3519 935
rect -3585 867 -3569 901
rect -3535 867 -3519 901
rect -3585 833 -3519 867
rect -3585 799 -3569 833
rect -3535 799 -3519 833
rect -3585 765 -3519 799
rect -3585 731 -3569 765
rect -3535 731 -3519 765
rect -3585 697 -3519 731
rect -3585 663 -3569 697
rect -3535 663 -3519 697
rect -3585 629 -3519 663
rect -3585 595 -3569 629
rect -3535 595 -3519 629
rect -3585 561 -3519 595
rect -3585 527 -3569 561
rect -3535 527 -3519 561
rect -3585 493 -3519 527
rect -3585 459 -3569 493
rect -3535 459 -3519 493
rect -3585 425 -3519 459
rect -3585 391 -3569 425
rect -3535 391 -3519 425
rect -3585 357 -3519 391
rect -3585 323 -3569 357
rect -3535 323 -3519 357
rect -3585 289 -3519 323
rect -3585 255 -3569 289
rect -3535 255 -3519 289
rect -3585 221 -3519 255
rect -3585 187 -3569 221
rect -3535 187 -3519 221
rect -3585 153 -3519 187
rect -3585 119 -3569 153
rect -3535 119 -3519 153
rect -3585 85 -3519 119
rect -3585 51 -3569 85
rect -3535 51 -3519 85
rect -3585 17 -3519 51
rect -3585 -17 -3569 17
rect -3535 -17 -3519 17
rect -3585 -51 -3519 -17
rect -3585 -85 -3569 -51
rect -3535 -85 -3519 -51
rect -3585 -119 -3519 -85
rect -3585 -153 -3569 -119
rect -3535 -153 -3519 -119
rect -3585 -187 -3519 -153
rect -3585 -221 -3569 -187
rect -3535 -221 -3519 -187
rect -3585 -255 -3519 -221
rect -3585 -289 -3569 -255
rect -3535 -289 -3519 -255
rect -3585 -323 -3519 -289
rect -3585 -357 -3569 -323
rect -3535 -357 -3519 -323
rect -3585 -391 -3519 -357
rect -3585 -425 -3569 -391
rect -3535 -425 -3519 -391
rect -3585 -459 -3519 -425
rect -3585 -493 -3569 -459
rect -3535 -493 -3519 -459
rect -3585 -527 -3519 -493
rect -3585 -561 -3569 -527
rect -3535 -561 -3519 -527
rect -3585 -595 -3519 -561
rect -3585 -629 -3569 -595
rect -3535 -629 -3519 -595
rect -3585 -663 -3519 -629
rect -3585 -697 -3569 -663
rect -3535 -697 -3519 -663
rect -3585 -731 -3519 -697
rect -3585 -765 -3569 -731
rect -3535 -765 -3519 -731
rect -3585 -799 -3519 -765
rect -3585 -833 -3569 -799
rect -3535 -833 -3519 -799
rect -3585 -867 -3519 -833
rect -3585 -901 -3569 -867
rect -3535 -901 -3519 -867
rect -3585 -935 -3519 -901
rect -3585 -969 -3569 -935
rect -3535 -969 -3519 -935
rect -3585 -1000 -3519 -969
rect -3489 969 -3423 1000
rect -3489 935 -3473 969
rect -3439 935 -3423 969
rect -3489 901 -3423 935
rect -3489 867 -3473 901
rect -3439 867 -3423 901
rect -3489 833 -3423 867
rect -3489 799 -3473 833
rect -3439 799 -3423 833
rect -3489 765 -3423 799
rect -3489 731 -3473 765
rect -3439 731 -3423 765
rect -3489 697 -3423 731
rect -3489 663 -3473 697
rect -3439 663 -3423 697
rect -3489 629 -3423 663
rect -3489 595 -3473 629
rect -3439 595 -3423 629
rect -3489 561 -3423 595
rect -3489 527 -3473 561
rect -3439 527 -3423 561
rect -3489 493 -3423 527
rect -3489 459 -3473 493
rect -3439 459 -3423 493
rect -3489 425 -3423 459
rect -3489 391 -3473 425
rect -3439 391 -3423 425
rect -3489 357 -3423 391
rect -3489 323 -3473 357
rect -3439 323 -3423 357
rect -3489 289 -3423 323
rect -3489 255 -3473 289
rect -3439 255 -3423 289
rect -3489 221 -3423 255
rect -3489 187 -3473 221
rect -3439 187 -3423 221
rect -3489 153 -3423 187
rect -3489 119 -3473 153
rect -3439 119 -3423 153
rect -3489 85 -3423 119
rect -3489 51 -3473 85
rect -3439 51 -3423 85
rect -3489 17 -3423 51
rect -3489 -17 -3473 17
rect -3439 -17 -3423 17
rect -3489 -51 -3423 -17
rect -3489 -85 -3473 -51
rect -3439 -85 -3423 -51
rect -3489 -119 -3423 -85
rect -3489 -153 -3473 -119
rect -3439 -153 -3423 -119
rect -3489 -187 -3423 -153
rect -3489 -221 -3473 -187
rect -3439 -221 -3423 -187
rect -3489 -255 -3423 -221
rect -3489 -289 -3473 -255
rect -3439 -289 -3423 -255
rect -3489 -323 -3423 -289
rect -3489 -357 -3473 -323
rect -3439 -357 -3423 -323
rect -3489 -391 -3423 -357
rect -3489 -425 -3473 -391
rect -3439 -425 -3423 -391
rect -3489 -459 -3423 -425
rect -3489 -493 -3473 -459
rect -3439 -493 -3423 -459
rect -3489 -527 -3423 -493
rect -3489 -561 -3473 -527
rect -3439 -561 -3423 -527
rect -3489 -595 -3423 -561
rect -3489 -629 -3473 -595
rect -3439 -629 -3423 -595
rect -3489 -663 -3423 -629
rect -3489 -697 -3473 -663
rect -3439 -697 -3423 -663
rect -3489 -731 -3423 -697
rect -3489 -765 -3473 -731
rect -3439 -765 -3423 -731
rect -3489 -799 -3423 -765
rect -3489 -833 -3473 -799
rect -3439 -833 -3423 -799
rect -3489 -867 -3423 -833
rect -3489 -901 -3473 -867
rect -3439 -901 -3423 -867
rect -3489 -935 -3423 -901
rect -3489 -969 -3473 -935
rect -3439 -969 -3423 -935
rect -3489 -1000 -3423 -969
rect -3393 969 -3327 1000
rect -3393 935 -3377 969
rect -3343 935 -3327 969
rect -3393 901 -3327 935
rect -3393 867 -3377 901
rect -3343 867 -3327 901
rect -3393 833 -3327 867
rect -3393 799 -3377 833
rect -3343 799 -3327 833
rect -3393 765 -3327 799
rect -3393 731 -3377 765
rect -3343 731 -3327 765
rect -3393 697 -3327 731
rect -3393 663 -3377 697
rect -3343 663 -3327 697
rect -3393 629 -3327 663
rect -3393 595 -3377 629
rect -3343 595 -3327 629
rect -3393 561 -3327 595
rect -3393 527 -3377 561
rect -3343 527 -3327 561
rect -3393 493 -3327 527
rect -3393 459 -3377 493
rect -3343 459 -3327 493
rect -3393 425 -3327 459
rect -3393 391 -3377 425
rect -3343 391 -3327 425
rect -3393 357 -3327 391
rect -3393 323 -3377 357
rect -3343 323 -3327 357
rect -3393 289 -3327 323
rect -3393 255 -3377 289
rect -3343 255 -3327 289
rect -3393 221 -3327 255
rect -3393 187 -3377 221
rect -3343 187 -3327 221
rect -3393 153 -3327 187
rect -3393 119 -3377 153
rect -3343 119 -3327 153
rect -3393 85 -3327 119
rect -3393 51 -3377 85
rect -3343 51 -3327 85
rect -3393 17 -3327 51
rect -3393 -17 -3377 17
rect -3343 -17 -3327 17
rect -3393 -51 -3327 -17
rect -3393 -85 -3377 -51
rect -3343 -85 -3327 -51
rect -3393 -119 -3327 -85
rect -3393 -153 -3377 -119
rect -3343 -153 -3327 -119
rect -3393 -187 -3327 -153
rect -3393 -221 -3377 -187
rect -3343 -221 -3327 -187
rect -3393 -255 -3327 -221
rect -3393 -289 -3377 -255
rect -3343 -289 -3327 -255
rect -3393 -323 -3327 -289
rect -3393 -357 -3377 -323
rect -3343 -357 -3327 -323
rect -3393 -391 -3327 -357
rect -3393 -425 -3377 -391
rect -3343 -425 -3327 -391
rect -3393 -459 -3327 -425
rect -3393 -493 -3377 -459
rect -3343 -493 -3327 -459
rect -3393 -527 -3327 -493
rect -3393 -561 -3377 -527
rect -3343 -561 -3327 -527
rect -3393 -595 -3327 -561
rect -3393 -629 -3377 -595
rect -3343 -629 -3327 -595
rect -3393 -663 -3327 -629
rect -3393 -697 -3377 -663
rect -3343 -697 -3327 -663
rect -3393 -731 -3327 -697
rect -3393 -765 -3377 -731
rect -3343 -765 -3327 -731
rect -3393 -799 -3327 -765
rect -3393 -833 -3377 -799
rect -3343 -833 -3327 -799
rect -3393 -867 -3327 -833
rect -3393 -901 -3377 -867
rect -3343 -901 -3327 -867
rect -3393 -935 -3327 -901
rect -3393 -969 -3377 -935
rect -3343 -969 -3327 -935
rect -3393 -1000 -3327 -969
rect -3297 969 -3231 1000
rect -3297 935 -3281 969
rect -3247 935 -3231 969
rect -3297 901 -3231 935
rect -3297 867 -3281 901
rect -3247 867 -3231 901
rect -3297 833 -3231 867
rect -3297 799 -3281 833
rect -3247 799 -3231 833
rect -3297 765 -3231 799
rect -3297 731 -3281 765
rect -3247 731 -3231 765
rect -3297 697 -3231 731
rect -3297 663 -3281 697
rect -3247 663 -3231 697
rect -3297 629 -3231 663
rect -3297 595 -3281 629
rect -3247 595 -3231 629
rect -3297 561 -3231 595
rect -3297 527 -3281 561
rect -3247 527 -3231 561
rect -3297 493 -3231 527
rect -3297 459 -3281 493
rect -3247 459 -3231 493
rect -3297 425 -3231 459
rect -3297 391 -3281 425
rect -3247 391 -3231 425
rect -3297 357 -3231 391
rect -3297 323 -3281 357
rect -3247 323 -3231 357
rect -3297 289 -3231 323
rect -3297 255 -3281 289
rect -3247 255 -3231 289
rect -3297 221 -3231 255
rect -3297 187 -3281 221
rect -3247 187 -3231 221
rect -3297 153 -3231 187
rect -3297 119 -3281 153
rect -3247 119 -3231 153
rect -3297 85 -3231 119
rect -3297 51 -3281 85
rect -3247 51 -3231 85
rect -3297 17 -3231 51
rect -3297 -17 -3281 17
rect -3247 -17 -3231 17
rect -3297 -51 -3231 -17
rect -3297 -85 -3281 -51
rect -3247 -85 -3231 -51
rect -3297 -119 -3231 -85
rect -3297 -153 -3281 -119
rect -3247 -153 -3231 -119
rect -3297 -187 -3231 -153
rect -3297 -221 -3281 -187
rect -3247 -221 -3231 -187
rect -3297 -255 -3231 -221
rect -3297 -289 -3281 -255
rect -3247 -289 -3231 -255
rect -3297 -323 -3231 -289
rect -3297 -357 -3281 -323
rect -3247 -357 -3231 -323
rect -3297 -391 -3231 -357
rect -3297 -425 -3281 -391
rect -3247 -425 -3231 -391
rect -3297 -459 -3231 -425
rect -3297 -493 -3281 -459
rect -3247 -493 -3231 -459
rect -3297 -527 -3231 -493
rect -3297 -561 -3281 -527
rect -3247 -561 -3231 -527
rect -3297 -595 -3231 -561
rect -3297 -629 -3281 -595
rect -3247 -629 -3231 -595
rect -3297 -663 -3231 -629
rect -3297 -697 -3281 -663
rect -3247 -697 -3231 -663
rect -3297 -731 -3231 -697
rect -3297 -765 -3281 -731
rect -3247 -765 -3231 -731
rect -3297 -799 -3231 -765
rect -3297 -833 -3281 -799
rect -3247 -833 -3231 -799
rect -3297 -867 -3231 -833
rect -3297 -901 -3281 -867
rect -3247 -901 -3231 -867
rect -3297 -935 -3231 -901
rect -3297 -969 -3281 -935
rect -3247 -969 -3231 -935
rect -3297 -1000 -3231 -969
rect -3201 969 -3135 1000
rect -3201 935 -3185 969
rect -3151 935 -3135 969
rect -3201 901 -3135 935
rect -3201 867 -3185 901
rect -3151 867 -3135 901
rect -3201 833 -3135 867
rect -3201 799 -3185 833
rect -3151 799 -3135 833
rect -3201 765 -3135 799
rect -3201 731 -3185 765
rect -3151 731 -3135 765
rect -3201 697 -3135 731
rect -3201 663 -3185 697
rect -3151 663 -3135 697
rect -3201 629 -3135 663
rect -3201 595 -3185 629
rect -3151 595 -3135 629
rect -3201 561 -3135 595
rect -3201 527 -3185 561
rect -3151 527 -3135 561
rect -3201 493 -3135 527
rect -3201 459 -3185 493
rect -3151 459 -3135 493
rect -3201 425 -3135 459
rect -3201 391 -3185 425
rect -3151 391 -3135 425
rect -3201 357 -3135 391
rect -3201 323 -3185 357
rect -3151 323 -3135 357
rect -3201 289 -3135 323
rect -3201 255 -3185 289
rect -3151 255 -3135 289
rect -3201 221 -3135 255
rect -3201 187 -3185 221
rect -3151 187 -3135 221
rect -3201 153 -3135 187
rect -3201 119 -3185 153
rect -3151 119 -3135 153
rect -3201 85 -3135 119
rect -3201 51 -3185 85
rect -3151 51 -3135 85
rect -3201 17 -3135 51
rect -3201 -17 -3185 17
rect -3151 -17 -3135 17
rect -3201 -51 -3135 -17
rect -3201 -85 -3185 -51
rect -3151 -85 -3135 -51
rect -3201 -119 -3135 -85
rect -3201 -153 -3185 -119
rect -3151 -153 -3135 -119
rect -3201 -187 -3135 -153
rect -3201 -221 -3185 -187
rect -3151 -221 -3135 -187
rect -3201 -255 -3135 -221
rect -3201 -289 -3185 -255
rect -3151 -289 -3135 -255
rect -3201 -323 -3135 -289
rect -3201 -357 -3185 -323
rect -3151 -357 -3135 -323
rect -3201 -391 -3135 -357
rect -3201 -425 -3185 -391
rect -3151 -425 -3135 -391
rect -3201 -459 -3135 -425
rect -3201 -493 -3185 -459
rect -3151 -493 -3135 -459
rect -3201 -527 -3135 -493
rect -3201 -561 -3185 -527
rect -3151 -561 -3135 -527
rect -3201 -595 -3135 -561
rect -3201 -629 -3185 -595
rect -3151 -629 -3135 -595
rect -3201 -663 -3135 -629
rect -3201 -697 -3185 -663
rect -3151 -697 -3135 -663
rect -3201 -731 -3135 -697
rect -3201 -765 -3185 -731
rect -3151 -765 -3135 -731
rect -3201 -799 -3135 -765
rect -3201 -833 -3185 -799
rect -3151 -833 -3135 -799
rect -3201 -867 -3135 -833
rect -3201 -901 -3185 -867
rect -3151 -901 -3135 -867
rect -3201 -935 -3135 -901
rect -3201 -969 -3185 -935
rect -3151 -969 -3135 -935
rect -3201 -1000 -3135 -969
rect -3105 969 -3039 1000
rect -3105 935 -3089 969
rect -3055 935 -3039 969
rect -3105 901 -3039 935
rect -3105 867 -3089 901
rect -3055 867 -3039 901
rect -3105 833 -3039 867
rect -3105 799 -3089 833
rect -3055 799 -3039 833
rect -3105 765 -3039 799
rect -3105 731 -3089 765
rect -3055 731 -3039 765
rect -3105 697 -3039 731
rect -3105 663 -3089 697
rect -3055 663 -3039 697
rect -3105 629 -3039 663
rect -3105 595 -3089 629
rect -3055 595 -3039 629
rect -3105 561 -3039 595
rect -3105 527 -3089 561
rect -3055 527 -3039 561
rect -3105 493 -3039 527
rect -3105 459 -3089 493
rect -3055 459 -3039 493
rect -3105 425 -3039 459
rect -3105 391 -3089 425
rect -3055 391 -3039 425
rect -3105 357 -3039 391
rect -3105 323 -3089 357
rect -3055 323 -3039 357
rect -3105 289 -3039 323
rect -3105 255 -3089 289
rect -3055 255 -3039 289
rect -3105 221 -3039 255
rect -3105 187 -3089 221
rect -3055 187 -3039 221
rect -3105 153 -3039 187
rect -3105 119 -3089 153
rect -3055 119 -3039 153
rect -3105 85 -3039 119
rect -3105 51 -3089 85
rect -3055 51 -3039 85
rect -3105 17 -3039 51
rect -3105 -17 -3089 17
rect -3055 -17 -3039 17
rect -3105 -51 -3039 -17
rect -3105 -85 -3089 -51
rect -3055 -85 -3039 -51
rect -3105 -119 -3039 -85
rect -3105 -153 -3089 -119
rect -3055 -153 -3039 -119
rect -3105 -187 -3039 -153
rect -3105 -221 -3089 -187
rect -3055 -221 -3039 -187
rect -3105 -255 -3039 -221
rect -3105 -289 -3089 -255
rect -3055 -289 -3039 -255
rect -3105 -323 -3039 -289
rect -3105 -357 -3089 -323
rect -3055 -357 -3039 -323
rect -3105 -391 -3039 -357
rect -3105 -425 -3089 -391
rect -3055 -425 -3039 -391
rect -3105 -459 -3039 -425
rect -3105 -493 -3089 -459
rect -3055 -493 -3039 -459
rect -3105 -527 -3039 -493
rect -3105 -561 -3089 -527
rect -3055 -561 -3039 -527
rect -3105 -595 -3039 -561
rect -3105 -629 -3089 -595
rect -3055 -629 -3039 -595
rect -3105 -663 -3039 -629
rect -3105 -697 -3089 -663
rect -3055 -697 -3039 -663
rect -3105 -731 -3039 -697
rect -3105 -765 -3089 -731
rect -3055 -765 -3039 -731
rect -3105 -799 -3039 -765
rect -3105 -833 -3089 -799
rect -3055 -833 -3039 -799
rect -3105 -867 -3039 -833
rect -3105 -901 -3089 -867
rect -3055 -901 -3039 -867
rect -3105 -935 -3039 -901
rect -3105 -969 -3089 -935
rect -3055 -969 -3039 -935
rect -3105 -1000 -3039 -969
rect -3009 969 -2943 1000
rect -3009 935 -2993 969
rect -2959 935 -2943 969
rect -3009 901 -2943 935
rect -3009 867 -2993 901
rect -2959 867 -2943 901
rect -3009 833 -2943 867
rect -3009 799 -2993 833
rect -2959 799 -2943 833
rect -3009 765 -2943 799
rect -3009 731 -2993 765
rect -2959 731 -2943 765
rect -3009 697 -2943 731
rect -3009 663 -2993 697
rect -2959 663 -2943 697
rect -3009 629 -2943 663
rect -3009 595 -2993 629
rect -2959 595 -2943 629
rect -3009 561 -2943 595
rect -3009 527 -2993 561
rect -2959 527 -2943 561
rect -3009 493 -2943 527
rect -3009 459 -2993 493
rect -2959 459 -2943 493
rect -3009 425 -2943 459
rect -3009 391 -2993 425
rect -2959 391 -2943 425
rect -3009 357 -2943 391
rect -3009 323 -2993 357
rect -2959 323 -2943 357
rect -3009 289 -2943 323
rect -3009 255 -2993 289
rect -2959 255 -2943 289
rect -3009 221 -2943 255
rect -3009 187 -2993 221
rect -2959 187 -2943 221
rect -3009 153 -2943 187
rect -3009 119 -2993 153
rect -2959 119 -2943 153
rect -3009 85 -2943 119
rect -3009 51 -2993 85
rect -2959 51 -2943 85
rect -3009 17 -2943 51
rect -3009 -17 -2993 17
rect -2959 -17 -2943 17
rect -3009 -51 -2943 -17
rect -3009 -85 -2993 -51
rect -2959 -85 -2943 -51
rect -3009 -119 -2943 -85
rect -3009 -153 -2993 -119
rect -2959 -153 -2943 -119
rect -3009 -187 -2943 -153
rect -3009 -221 -2993 -187
rect -2959 -221 -2943 -187
rect -3009 -255 -2943 -221
rect -3009 -289 -2993 -255
rect -2959 -289 -2943 -255
rect -3009 -323 -2943 -289
rect -3009 -357 -2993 -323
rect -2959 -357 -2943 -323
rect -3009 -391 -2943 -357
rect -3009 -425 -2993 -391
rect -2959 -425 -2943 -391
rect -3009 -459 -2943 -425
rect -3009 -493 -2993 -459
rect -2959 -493 -2943 -459
rect -3009 -527 -2943 -493
rect -3009 -561 -2993 -527
rect -2959 -561 -2943 -527
rect -3009 -595 -2943 -561
rect -3009 -629 -2993 -595
rect -2959 -629 -2943 -595
rect -3009 -663 -2943 -629
rect -3009 -697 -2993 -663
rect -2959 -697 -2943 -663
rect -3009 -731 -2943 -697
rect -3009 -765 -2993 -731
rect -2959 -765 -2943 -731
rect -3009 -799 -2943 -765
rect -3009 -833 -2993 -799
rect -2959 -833 -2943 -799
rect -3009 -867 -2943 -833
rect -3009 -901 -2993 -867
rect -2959 -901 -2943 -867
rect -3009 -935 -2943 -901
rect -3009 -969 -2993 -935
rect -2959 -969 -2943 -935
rect -3009 -1000 -2943 -969
rect -2913 969 -2847 1000
rect -2913 935 -2897 969
rect -2863 935 -2847 969
rect -2913 901 -2847 935
rect -2913 867 -2897 901
rect -2863 867 -2847 901
rect -2913 833 -2847 867
rect -2913 799 -2897 833
rect -2863 799 -2847 833
rect -2913 765 -2847 799
rect -2913 731 -2897 765
rect -2863 731 -2847 765
rect -2913 697 -2847 731
rect -2913 663 -2897 697
rect -2863 663 -2847 697
rect -2913 629 -2847 663
rect -2913 595 -2897 629
rect -2863 595 -2847 629
rect -2913 561 -2847 595
rect -2913 527 -2897 561
rect -2863 527 -2847 561
rect -2913 493 -2847 527
rect -2913 459 -2897 493
rect -2863 459 -2847 493
rect -2913 425 -2847 459
rect -2913 391 -2897 425
rect -2863 391 -2847 425
rect -2913 357 -2847 391
rect -2913 323 -2897 357
rect -2863 323 -2847 357
rect -2913 289 -2847 323
rect -2913 255 -2897 289
rect -2863 255 -2847 289
rect -2913 221 -2847 255
rect -2913 187 -2897 221
rect -2863 187 -2847 221
rect -2913 153 -2847 187
rect -2913 119 -2897 153
rect -2863 119 -2847 153
rect -2913 85 -2847 119
rect -2913 51 -2897 85
rect -2863 51 -2847 85
rect -2913 17 -2847 51
rect -2913 -17 -2897 17
rect -2863 -17 -2847 17
rect -2913 -51 -2847 -17
rect -2913 -85 -2897 -51
rect -2863 -85 -2847 -51
rect -2913 -119 -2847 -85
rect -2913 -153 -2897 -119
rect -2863 -153 -2847 -119
rect -2913 -187 -2847 -153
rect -2913 -221 -2897 -187
rect -2863 -221 -2847 -187
rect -2913 -255 -2847 -221
rect -2913 -289 -2897 -255
rect -2863 -289 -2847 -255
rect -2913 -323 -2847 -289
rect -2913 -357 -2897 -323
rect -2863 -357 -2847 -323
rect -2913 -391 -2847 -357
rect -2913 -425 -2897 -391
rect -2863 -425 -2847 -391
rect -2913 -459 -2847 -425
rect -2913 -493 -2897 -459
rect -2863 -493 -2847 -459
rect -2913 -527 -2847 -493
rect -2913 -561 -2897 -527
rect -2863 -561 -2847 -527
rect -2913 -595 -2847 -561
rect -2913 -629 -2897 -595
rect -2863 -629 -2847 -595
rect -2913 -663 -2847 -629
rect -2913 -697 -2897 -663
rect -2863 -697 -2847 -663
rect -2913 -731 -2847 -697
rect -2913 -765 -2897 -731
rect -2863 -765 -2847 -731
rect -2913 -799 -2847 -765
rect -2913 -833 -2897 -799
rect -2863 -833 -2847 -799
rect -2913 -867 -2847 -833
rect -2913 -901 -2897 -867
rect -2863 -901 -2847 -867
rect -2913 -935 -2847 -901
rect -2913 -969 -2897 -935
rect -2863 -969 -2847 -935
rect -2913 -1000 -2847 -969
rect -2817 969 -2751 1000
rect -2817 935 -2801 969
rect -2767 935 -2751 969
rect -2817 901 -2751 935
rect -2817 867 -2801 901
rect -2767 867 -2751 901
rect -2817 833 -2751 867
rect -2817 799 -2801 833
rect -2767 799 -2751 833
rect -2817 765 -2751 799
rect -2817 731 -2801 765
rect -2767 731 -2751 765
rect -2817 697 -2751 731
rect -2817 663 -2801 697
rect -2767 663 -2751 697
rect -2817 629 -2751 663
rect -2817 595 -2801 629
rect -2767 595 -2751 629
rect -2817 561 -2751 595
rect -2817 527 -2801 561
rect -2767 527 -2751 561
rect -2817 493 -2751 527
rect -2817 459 -2801 493
rect -2767 459 -2751 493
rect -2817 425 -2751 459
rect -2817 391 -2801 425
rect -2767 391 -2751 425
rect -2817 357 -2751 391
rect -2817 323 -2801 357
rect -2767 323 -2751 357
rect -2817 289 -2751 323
rect -2817 255 -2801 289
rect -2767 255 -2751 289
rect -2817 221 -2751 255
rect -2817 187 -2801 221
rect -2767 187 -2751 221
rect -2817 153 -2751 187
rect -2817 119 -2801 153
rect -2767 119 -2751 153
rect -2817 85 -2751 119
rect -2817 51 -2801 85
rect -2767 51 -2751 85
rect -2817 17 -2751 51
rect -2817 -17 -2801 17
rect -2767 -17 -2751 17
rect -2817 -51 -2751 -17
rect -2817 -85 -2801 -51
rect -2767 -85 -2751 -51
rect -2817 -119 -2751 -85
rect -2817 -153 -2801 -119
rect -2767 -153 -2751 -119
rect -2817 -187 -2751 -153
rect -2817 -221 -2801 -187
rect -2767 -221 -2751 -187
rect -2817 -255 -2751 -221
rect -2817 -289 -2801 -255
rect -2767 -289 -2751 -255
rect -2817 -323 -2751 -289
rect -2817 -357 -2801 -323
rect -2767 -357 -2751 -323
rect -2817 -391 -2751 -357
rect -2817 -425 -2801 -391
rect -2767 -425 -2751 -391
rect -2817 -459 -2751 -425
rect -2817 -493 -2801 -459
rect -2767 -493 -2751 -459
rect -2817 -527 -2751 -493
rect -2817 -561 -2801 -527
rect -2767 -561 -2751 -527
rect -2817 -595 -2751 -561
rect -2817 -629 -2801 -595
rect -2767 -629 -2751 -595
rect -2817 -663 -2751 -629
rect -2817 -697 -2801 -663
rect -2767 -697 -2751 -663
rect -2817 -731 -2751 -697
rect -2817 -765 -2801 -731
rect -2767 -765 -2751 -731
rect -2817 -799 -2751 -765
rect -2817 -833 -2801 -799
rect -2767 -833 -2751 -799
rect -2817 -867 -2751 -833
rect -2817 -901 -2801 -867
rect -2767 -901 -2751 -867
rect -2817 -935 -2751 -901
rect -2817 -969 -2801 -935
rect -2767 -969 -2751 -935
rect -2817 -1000 -2751 -969
rect -2721 969 -2655 1000
rect -2721 935 -2705 969
rect -2671 935 -2655 969
rect -2721 901 -2655 935
rect -2721 867 -2705 901
rect -2671 867 -2655 901
rect -2721 833 -2655 867
rect -2721 799 -2705 833
rect -2671 799 -2655 833
rect -2721 765 -2655 799
rect -2721 731 -2705 765
rect -2671 731 -2655 765
rect -2721 697 -2655 731
rect -2721 663 -2705 697
rect -2671 663 -2655 697
rect -2721 629 -2655 663
rect -2721 595 -2705 629
rect -2671 595 -2655 629
rect -2721 561 -2655 595
rect -2721 527 -2705 561
rect -2671 527 -2655 561
rect -2721 493 -2655 527
rect -2721 459 -2705 493
rect -2671 459 -2655 493
rect -2721 425 -2655 459
rect -2721 391 -2705 425
rect -2671 391 -2655 425
rect -2721 357 -2655 391
rect -2721 323 -2705 357
rect -2671 323 -2655 357
rect -2721 289 -2655 323
rect -2721 255 -2705 289
rect -2671 255 -2655 289
rect -2721 221 -2655 255
rect -2721 187 -2705 221
rect -2671 187 -2655 221
rect -2721 153 -2655 187
rect -2721 119 -2705 153
rect -2671 119 -2655 153
rect -2721 85 -2655 119
rect -2721 51 -2705 85
rect -2671 51 -2655 85
rect -2721 17 -2655 51
rect -2721 -17 -2705 17
rect -2671 -17 -2655 17
rect -2721 -51 -2655 -17
rect -2721 -85 -2705 -51
rect -2671 -85 -2655 -51
rect -2721 -119 -2655 -85
rect -2721 -153 -2705 -119
rect -2671 -153 -2655 -119
rect -2721 -187 -2655 -153
rect -2721 -221 -2705 -187
rect -2671 -221 -2655 -187
rect -2721 -255 -2655 -221
rect -2721 -289 -2705 -255
rect -2671 -289 -2655 -255
rect -2721 -323 -2655 -289
rect -2721 -357 -2705 -323
rect -2671 -357 -2655 -323
rect -2721 -391 -2655 -357
rect -2721 -425 -2705 -391
rect -2671 -425 -2655 -391
rect -2721 -459 -2655 -425
rect -2721 -493 -2705 -459
rect -2671 -493 -2655 -459
rect -2721 -527 -2655 -493
rect -2721 -561 -2705 -527
rect -2671 -561 -2655 -527
rect -2721 -595 -2655 -561
rect -2721 -629 -2705 -595
rect -2671 -629 -2655 -595
rect -2721 -663 -2655 -629
rect -2721 -697 -2705 -663
rect -2671 -697 -2655 -663
rect -2721 -731 -2655 -697
rect -2721 -765 -2705 -731
rect -2671 -765 -2655 -731
rect -2721 -799 -2655 -765
rect -2721 -833 -2705 -799
rect -2671 -833 -2655 -799
rect -2721 -867 -2655 -833
rect -2721 -901 -2705 -867
rect -2671 -901 -2655 -867
rect -2721 -935 -2655 -901
rect -2721 -969 -2705 -935
rect -2671 -969 -2655 -935
rect -2721 -1000 -2655 -969
rect -2625 969 -2559 1000
rect -2625 935 -2609 969
rect -2575 935 -2559 969
rect -2625 901 -2559 935
rect -2625 867 -2609 901
rect -2575 867 -2559 901
rect -2625 833 -2559 867
rect -2625 799 -2609 833
rect -2575 799 -2559 833
rect -2625 765 -2559 799
rect -2625 731 -2609 765
rect -2575 731 -2559 765
rect -2625 697 -2559 731
rect -2625 663 -2609 697
rect -2575 663 -2559 697
rect -2625 629 -2559 663
rect -2625 595 -2609 629
rect -2575 595 -2559 629
rect -2625 561 -2559 595
rect -2625 527 -2609 561
rect -2575 527 -2559 561
rect -2625 493 -2559 527
rect -2625 459 -2609 493
rect -2575 459 -2559 493
rect -2625 425 -2559 459
rect -2625 391 -2609 425
rect -2575 391 -2559 425
rect -2625 357 -2559 391
rect -2625 323 -2609 357
rect -2575 323 -2559 357
rect -2625 289 -2559 323
rect -2625 255 -2609 289
rect -2575 255 -2559 289
rect -2625 221 -2559 255
rect -2625 187 -2609 221
rect -2575 187 -2559 221
rect -2625 153 -2559 187
rect -2625 119 -2609 153
rect -2575 119 -2559 153
rect -2625 85 -2559 119
rect -2625 51 -2609 85
rect -2575 51 -2559 85
rect -2625 17 -2559 51
rect -2625 -17 -2609 17
rect -2575 -17 -2559 17
rect -2625 -51 -2559 -17
rect -2625 -85 -2609 -51
rect -2575 -85 -2559 -51
rect -2625 -119 -2559 -85
rect -2625 -153 -2609 -119
rect -2575 -153 -2559 -119
rect -2625 -187 -2559 -153
rect -2625 -221 -2609 -187
rect -2575 -221 -2559 -187
rect -2625 -255 -2559 -221
rect -2625 -289 -2609 -255
rect -2575 -289 -2559 -255
rect -2625 -323 -2559 -289
rect -2625 -357 -2609 -323
rect -2575 -357 -2559 -323
rect -2625 -391 -2559 -357
rect -2625 -425 -2609 -391
rect -2575 -425 -2559 -391
rect -2625 -459 -2559 -425
rect -2625 -493 -2609 -459
rect -2575 -493 -2559 -459
rect -2625 -527 -2559 -493
rect -2625 -561 -2609 -527
rect -2575 -561 -2559 -527
rect -2625 -595 -2559 -561
rect -2625 -629 -2609 -595
rect -2575 -629 -2559 -595
rect -2625 -663 -2559 -629
rect -2625 -697 -2609 -663
rect -2575 -697 -2559 -663
rect -2625 -731 -2559 -697
rect -2625 -765 -2609 -731
rect -2575 -765 -2559 -731
rect -2625 -799 -2559 -765
rect -2625 -833 -2609 -799
rect -2575 -833 -2559 -799
rect -2625 -867 -2559 -833
rect -2625 -901 -2609 -867
rect -2575 -901 -2559 -867
rect -2625 -935 -2559 -901
rect -2625 -969 -2609 -935
rect -2575 -969 -2559 -935
rect -2625 -1000 -2559 -969
rect -2529 969 -2463 1000
rect -2529 935 -2513 969
rect -2479 935 -2463 969
rect -2529 901 -2463 935
rect -2529 867 -2513 901
rect -2479 867 -2463 901
rect -2529 833 -2463 867
rect -2529 799 -2513 833
rect -2479 799 -2463 833
rect -2529 765 -2463 799
rect -2529 731 -2513 765
rect -2479 731 -2463 765
rect -2529 697 -2463 731
rect -2529 663 -2513 697
rect -2479 663 -2463 697
rect -2529 629 -2463 663
rect -2529 595 -2513 629
rect -2479 595 -2463 629
rect -2529 561 -2463 595
rect -2529 527 -2513 561
rect -2479 527 -2463 561
rect -2529 493 -2463 527
rect -2529 459 -2513 493
rect -2479 459 -2463 493
rect -2529 425 -2463 459
rect -2529 391 -2513 425
rect -2479 391 -2463 425
rect -2529 357 -2463 391
rect -2529 323 -2513 357
rect -2479 323 -2463 357
rect -2529 289 -2463 323
rect -2529 255 -2513 289
rect -2479 255 -2463 289
rect -2529 221 -2463 255
rect -2529 187 -2513 221
rect -2479 187 -2463 221
rect -2529 153 -2463 187
rect -2529 119 -2513 153
rect -2479 119 -2463 153
rect -2529 85 -2463 119
rect -2529 51 -2513 85
rect -2479 51 -2463 85
rect -2529 17 -2463 51
rect -2529 -17 -2513 17
rect -2479 -17 -2463 17
rect -2529 -51 -2463 -17
rect -2529 -85 -2513 -51
rect -2479 -85 -2463 -51
rect -2529 -119 -2463 -85
rect -2529 -153 -2513 -119
rect -2479 -153 -2463 -119
rect -2529 -187 -2463 -153
rect -2529 -221 -2513 -187
rect -2479 -221 -2463 -187
rect -2529 -255 -2463 -221
rect -2529 -289 -2513 -255
rect -2479 -289 -2463 -255
rect -2529 -323 -2463 -289
rect -2529 -357 -2513 -323
rect -2479 -357 -2463 -323
rect -2529 -391 -2463 -357
rect -2529 -425 -2513 -391
rect -2479 -425 -2463 -391
rect -2529 -459 -2463 -425
rect -2529 -493 -2513 -459
rect -2479 -493 -2463 -459
rect -2529 -527 -2463 -493
rect -2529 -561 -2513 -527
rect -2479 -561 -2463 -527
rect -2529 -595 -2463 -561
rect -2529 -629 -2513 -595
rect -2479 -629 -2463 -595
rect -2529 -663 -2463 -629
rect -2529 -697 -2513 -663
rect -2479 -697 -2463 -663
rect -2529 -731 -2463 -697
rect -2529 -765 -2513 -731
rect -2479 -765 -2463 -731
rect -2529 -799 -2463 -765
rect -2529 -833 -2513 -799
rect -2479 -833 -2463 -799
rect -2529 -867 -2463 -833
rect -2529 -901 -2513 -867
rect -2479 -901 -2463 -867
rect -2529 -935 -2463 -901
rect -2529 -969 -2513 -935
rect -2479 -969 -2463 -935
rect -2529 -1000 -2463 -969
rect -2433 969 -2367 1000
rect -2433 935 -2417 969
rect -2383 935 -2367 969
rect -2433 901 -2367 935
rect -2433 867 -2417 901
rect -2383 867 -2367 901
rect -2433 833 -2367 867
rect -2433 799 -2417 833
rect -2383 799 -2367 833
rect -2433 765 -2367 799
rect -2433 731 -2417 765
rect -2383 731 -2367 765
rect -2433 697 -2367 731
rect -2433 663 -2417 697
rect -2383 663 -2367 697
rect -2433 629 -2367 663
rect -2433 595 -2417 629
rect -2383 595 -2367 629
rect -2433 561 -2367 595
rect -2433 527 -2417 561
rect -2383 527 -2367 561
rect -2433 493 -2367 527
rect -2433 459 -2417 493
rect -2383 459 -2367 493
rect -2433 425 -2367 459
rect -2433 391 -2417 425
rect -2383 391 -2367 425
rect -2433 357 -2367 391
rect -2433 323 -2417 357
rect -2383 323 -2367 357
rect -2433 289 -2367 323
rect -2433 255 -2417 289
rect -2383 255 -2367 289
rect -2433 221 -2367 255
rect -2433 187 -2417 221
rect -2383 187 -2367 221
rect -2433 153 -2367 187
rect -2433 119 -2417 153
rect -2383 119 -2367 153
rect -2433 85 -2367 119
rect -2433 51 -2417 85
rect -2383 51 -2367 85
rect -2433 17 -2367 51
rect -2433 -17 -2417 17
rect -2383 -17 -2367 17
rect -2433 -51 -2367 -17
rect -2433 -85 -2417 -51
rect -2383 -85 -2367 -51
rect -2433 -119 -2367 -85
rect -2433 -153 -2417 -119
rect -2383 -153 -2367 -119
rect -2433 -187 -2367 -153
rect -2433 -221 -2417 -187
rect -2383 -221 -2367 -187
rect -2433 -255 -2367 -221
rect -2433 -289 -2417 -255
rect -2383 -289 -2367 -255
rect -2433 -323 -2367 -289
rect -2433 -357 -2417 -323
rect -2383 -357 -2367 -323
rect -2433 -391 -2367 -357
rect -2433 -425 -2417 -391
rect -2383 -425 -2367 -391
rect -2433 -459 -2367 -425
rect -2433 -493 -2417 -459
rect -2383 -493 -2367 -459
rect -2433 -527 -2367 -493
rect -2433 -561 -2417 -527
rect -2383 -561 -2367 -527
rect -2433 -595 -2367 -561
rect -2433 -629 -2417 -595
rect -2383 -629 -2367 -595
rect -2433 -663 -2367 -629
rect -2433 -697 -2417 -663
rect -2383 -697 -2367 -663
rect -2433 -731 -2367 -697
rect -2433 -765 -2417 -731
rect -2383 -765 -2367 -731
rect -2433 -799 -2367 -765
rect -2433 -833 -2417 -799
rect -2383 -833 -2367 -799
rect -2433 -867 -2367 -833
rect -2433 -901 -2417 -867
rect -2383 -901 -2367 -867
rect -2433 -935 -2367 -901
rect -2433 -969 -2417 -935
rect -2383 -969 -2367 -935
rect -2433 -1000 -2367 -969
rect -2337 969 -2271 1000
rect -2337 935 -2321 969
rect -2287 935 -2271 969
rect -2337 901 -2271 935
rect -2337 867 -2321 901
rect -2287 867 -2271 901
rect -2337 833 -2271 867
rect -2337 799 -2321 833
rect -2287 799 -2271 833
rect -2337 765 -2271 799
rect -2337 731 -2321 765
rect -2287 731 -2271 765
rect -2337 697 -2271 731
rect -2337 663 -2321 697
rect -2287 663 -2271 697
rect -2337 629 -2271 663
rect -2337 595 -2321 629
rect -2287 595 -2271 629
rect -2337 561 -2271 595
rect -2337 527 -2321 561
rect -2287 527 -2271 561
rect -2337 493 -2271 527
rect -2337 459 -2321 493
rect -2287 459 -2271 493
rect -2337 425 -2271 459
rect -2337 391 -2321 425
rect -2287 391 -2271 425
rect -2337 357 -2271 391
rect -2337 323 -2321 357
rect -2287 323 -2271 357
rect -2337 289 -2271 323
rect -2337 255 -2321 289
rect -2287 255 -2271 289
rect -2337 221 -2271 255
rect -2337 187 -2321 221
rect -2287 187 -2271 221
rect -2337 153 -2271 187
rect -2337 119 -2321 153
rect -2287 119 -2271 153
rect -2337 85 -2271 119
rect -2337 51 -2321 85
rect -2287 51 -2271 85
rect -2337 17 -2271 51
rect -2337 -17 -2321 17
rect -2287 -17 -2271 17
rect -2337 -51 -2271 -17
rect -2337 -85 -2321 -51
rect -2287 -85 -2271 -51
rect -2337 -119 -2271 -85
rect -2337 -153 -2321 -119
rect -2287 -153 -2271 -119
rect -2337 -187 -2271 -153
rect -2337 -221 -2321 -187
rect -2287 -221 -2271 -187
rect -2337 -255 -2271 -221
rect -2337 -289 -2321 -255
rect -2287 -289 -2271 -255
rect -2337 -323 -2271 -289
rect -2337 -357 -2321 -323
rect -2287 -357 -2271 -323
rect -2337 -391 -2271 -357
rect -2337 -425 -2321 -391
rect -2287 -425 -2271 -391
rect -2337 -459 -2271 -425
rect -2337 -493 -2321 -459
rect -2287 -493 -2271 -459
rect -2337 -527 -2271 -493
rect -2337 -561 -2321 -527
rect -2287 -561 -2271 -527
rect -2337 -595 -2271 -561
rect -2337 -629 -2321 -595
rect -2287 -629 -2271 -595
rect -2337 -663 -2271 -629
rect -2337 -697 -2321 -663
rect -2287 -697 -2271 -663
rect -2337 -731 -2271 -697
rect -2337 -765 -2321 -731
rect -2287 -765 -2271 -731
rect -2337 -799 -2271 -765
rect -2337 -833 -2321 -799
rect -2287 -833 -2271 -799
rect -2337 -867 -2271 -833
rect -2337 -901 -2321 -867
rect -2287 -901 -2271 -867
rect -2337 -935 -2271 -901
rect -2337 -969 -2321 -935
rect -2287 -969 -2271 -935
rect -2337 -1000 -2271 -969
rect -2241 969 -2175 1000
rect -2241 935 -2225 969
rect -2191 935 -2175 969
rect -2241 901 -2175 935
rect -2241 867 -2225 901
rect -2191 867 -2175 901
rect -2241 833 -2175 867
rect -2241 799 -2225 833
rect -2191 799 -2175 833
rect -2241 765 -2175 799
rect -2241 731 -2225 765
rect -2191 731 -2175 765
rect -2241 697 -2175 731
rect -2241 663 -2225 697
rect -2191 663 -2175 697
rect -2241 629 -2175 663
rect -2241 595 -2225 629
rect -2191 595 -2175 629
rect -2241 561 -2175 595
rect -2241 527 -2225 561
rect -2191 527 -2175 561
rect -2241 493 -2175 527
rect -2241 459 -2225 493
rect -2191 459 -2175 493
rect -2241 425 -2175 459
rect -2241 391 -2225 425
rect -2191 391 -2175 425
rect -2241 357 -2175 391
rect -2241 323 -2225 357
rect -2191 323 -2175 357
rect -2241 289 -2175 323
rect -2241 255 -2225 289
rect -2191 255 -2175 289
rect -2241 221 -2175 255
rect -2241 187 -2225 221
rect -2191 187 -2175 221
rect -2241 153 -2175 187
rect -2241 119 -2225 153
rect -2191 119 -2175 153
rect -2241 85 -2175 119
rect -2241 51 -2225 85
rect -2191 51 -2175 85
rect -2241 17 -2175 51
rect -2241 -17 -2225 17
rect -2191 -17 -2175 17
rect -2241 -51 -2175 -17
rect -2241 -85 -2225 -51
rect -2191 -85 -2175 -51
rect -2241 -119 -2175 -85
rect -2241 -153 -2225 -119
rect -2191 -153 -2175 -119
rect -2241 -187 -2175 -153
rect -2241 -221 -2225 -187
rect -2191 -221 -2175 -187
rect -2241 -255 -2175 -221
rect -2241 -289 -2225 -255
rect -2191 -289 -2175 -255
rect -2241 -323 -2175 -289
rect -2241 -357 -2225 -323
rect -2191 -357 -2175 -323
rect -2241 -391 -2175 -357
rect -2241 -425 -2225 -391
rect -2191 -425 -2175 -391
rect -2241 -459 -2175 -425
rect -2241 -493 -2225 -459
rect -2191 -493 -2175 -459
rect -2241 -527 -2175 -493
rect -2241 -561 -2225 -527
rect -2191 -561 -2175 -527
rect -2241 -595 -2175 -561
rect -2241 -629 -2225 -595
rect -2191 -629 -2175 -595
rect -2241 -663 -2175 -629
rect -2241 -697 -2225 -663
rect -2191 -697 -2175 -663
rect -2241 -731 -2175 -697
rect -2241 -765 -2225 -731
rect -2191 -765 -2175 -731
rect -2241 -799 -2175 -765
rect -2241 -833 -2225 -799
rect -2191 -833 -2175 -799
rect -2241 -867 -2175 -833
rect -2241 -901 -2225 -867
rect -2191 -901 -2175 -867
rect -2241 -935 -2175 -901
rect -2241 -969 -2225 -935
rect -2191 -969 -2175 -935
rect -2241 -1000 -2175 -969
rect -2145 969 -2079 1000
rect -2145 935 -2129 969
rect -2095 935 -2079 969
rect -2145 901 -2079 935
rect -2145 867 -2129 901
rect -2095 867 -2079 901
rect -2145 833 -2079 867
rect -2145 799 -2129 833
rect -2095 799 -2079 833
rect -2145 765 -2079 799
rect -2145 731 -2129 765
rect -2095 731 -2079 765
rect -2145 697 -2079 731
rect -2145 663 -2129 697
rect -2095 663 -2079 697
rect -2145 629 -2079 663
rect -2145 595 -2129 629
rect -2095 595 -2079 629
rect -2145 561 -2079 595
rect -2145 527 -2129 561
rect -2095 527 -2079 561
rect -2145 493 -2079 527
rect -2145 459 -2129 493
rect -2095 459 -2079 493
rect -2145 425 -2079 459
rect -2145 391 -2129 425
rect -2095 391 -2079 425
rect -2145 357 -2079 391
rect -2145 323 -2129 357
rect -2095 323 -2079 357
rect -2145 289 -2079 323
rect -2145 255 -2129 289
rect -2095 255 -2079 289
rect -2145 221 -2079 255
rect -2145 187 -2129 221
rect -2095 187 -2079 221
rect -2145 153 -2079 187
rect -2145 119 -2129 153
rect -2095 119 -2079 153
rect -2145 85 -2079 119
rect -2145 51 -2129 85
rect -2095 51 -2079 85
rect -2145 17 -2079 51
rect -2145 -17 -2129 17
rect -2095 -17 -2079 17
rect -2145 -51 -2079 -17
rect -2145 -85 -2129 -51
rect -2095 -85 -2079 -51
rect -2145 -119 -2079 -85
rect -2145 -153 -2129 -119
rect -2095 -153 -2079 -119
rect -2145 -187 -2079 -153
rect -2145 -221 -2129 -187
rect -2095 -221 -2079 -187
rect -2145 -255 -2079 -221
rect -2145 -289 -2129 -255
rect -2095 -289 -2079 -255
rect -2145 -323 -2079 -289
rect -2145 -357 -2129 -323
rect -2095 -357 -2079 -323
rect -2145 -391 -2079 -357
rect -2145 -425 -2129 -391
rect -2095 -425 -2079 -391
rect -2145 -459 -2079 -425
rect -2145 -493 -2129 -459
rect -2095 -493 -2079 -459
rect -2145 -527 -2079 -493
rect -2145 -561 -2129 -527
rect -2095 -561 -2079 -527
rect -2145 -595 -2079 -561
rect -2145 -629 -2129 -595
rect -2095 -629 -2079 -595
rect -2145 -663 -2079 -629
rect -2145 -697 -2129 -663
rect -2095 -697 -2079 -663
rect -2145 -731 -2079 -697
rect -2145 -765 -2129 -731
rect -2095 -765 -2079 -731
rect -2145 -799 -2079 -765
rect -2145 -833 -2129 -799
rect -2095 -833 -2079 -799
rect -2145 -867 -2079 -833
rect -2145 -901 -2129 -867
rect -2095 -901 -2079 -867
rect -2145 -935 -2079 -901
rect -2145 -969 -2129 -935
rect -2095 -969 -2079 -935
rect -2145 -1000 -2079 -969
rect -2049 969 -1983 1000
rect -2049 935 -2033 969
rect -1999 935 -1983 969
rect -2049 901 -1983 935
rect -2049 867 -2033 901
rect -1999 867 -1983 901
rect -2049 833 -1983 867
rect -2049 799 -2033 833
rect -1999 799 -1983 833
rect -2049 765 -1983 799
rect -2049 731 -2033 765
rect -1999 731 -1983 765
rect -2049 697 -1983 731
rect -2049 663 -2033 697
rect -1999 663 -1983 697
rect -2049 629 -1983 663
rect -2049 595 -2033 629
rect -1999 595 -1983 629
rect -2049 561 -1983 595
rect -2049 527 -2033 561
rect -1999 527 -1983 561
rect -2049 493 -1983 527
rect -2049 459 -2033 493
rect -1999 459 -1983 493
rect -2049 425 -1983 459
rect -2049 391 -2033 425
rect -1999 391 -1983 425
rect -2049 357 -1983 391
rect -2049 323 -2033 357
rect -1999 323 -1983 357
rect -2049 289 -1983 323
rect -2049 255 -2033 289
rect -1999 255 -1983 289
rect -2049 221 -1983 255
rect -2049 187 -2033 221
rect -1999 187 -1983 221
rect -2049 153 -1983 187
rect -2049 119 -2033 153
rect -1999 119 -1983 153
rect -2049 85 -1983 119
rect -2049 51 -2033 85
rect -1999 51 -1983 85
rect -2049 17 -1983 51
rect -2049 -17 -2033 17
rect -1999 -17 -1983 17
rect -2049 -51 -1983 -17
rect -2049 -85 -2033 -51
rect -1999 -85 -1983 -51
rect -2049 -119 -1983 -85
rect -2049 -153 -2033 -119
rect -1999 -153 -1983 -119
rect -2049 -187 -1983 -153
rect -2049 -221 -2033 -187
rect -1999 -221 -1983 -187
rect -2049 -255 -1983 -221
rect -2049 -289 -2033 -255
rect -1999 -289 -1983 -255
rect -2049 -323 -1983 -289
rect -2049 -357 -2033 -323
rect -1999 -357 -1983 -323
rect -2049 -391 -1983 -357
rect -2049 -425 -2033 -391
rect -1999 -425 -1983 -391
rect -2049 -459 -1983 -425
rect -2049 -493 -2033 -459
rect -1999 -493 -1983 -459
rect -2049 -527 -1983 -493
rect -2049 -561 -2033 -527
rect -1999 -561 -1983 -527
rect -2049 -595 -1983 -561
rect -2049 -629 -2033 -595
rect -1999 -629 -1983 -595
rect -2049 -663 -1983 -629
rect -2049 -697 -2033 -663
rect -1999 -697 -1983 -663
rect -2049 -731 -1983 -697
rect -2049 -765 -2033 -731
rect -1999 -765 -1983 -731
rect -2049 -799 -1983 -765
rect -2049 -833 -2033 -799
rect -1999 -833 -1983 -799
rect -2049 -867 -1983 -833
rect -2049 -901 -2033 -867
rect -1999 -901 -1983 -867
rect -2049 -935 -1983 -901
rect -2049 -969 -2033 -935
rect -1999 -969 -1983 -935
rect -2049 -1000 -1983 -969
rect -1953 969 -1887 1000
rect -1953 935 -1937 969
rect -1903 935 -1887 969
rect -1953 901 -1887 935
rect -1953 867 -1937 901
rect -1903 867 -1887 901
rect -1953 833 -1887 867
rect -1953 799 -1937 833
rect -1903 799 -1887 833
rect -1953 765 -1887 799
rect -1953 731 -1937 765
rect -1903 731 -1887 765
rect -1953 697 -1887 731
rect -1953 663 -1937 697
rect -1903 663 -1887 697
rect -1953 629 -1887 663
rect -1953 595 -1937 629
rect -1903 595 -1887 629
rect -1953 561 -1887 595
rect -1953 527 -1937 561
rect -1903 527 -1887 561
rect -1953 493 -1887 527
rect -1953 459 -1937 493
rect -1903 459 -1887 493
rect -1953 425 -1887 459
rect -1953 391 -1937 425
rect -1903 391 -1887 425
rect -1953 357 -1887 391
rect -1953 323 -1937 357
rect -1903 323 -1887 357
rect -1953 289 -1887 323
rect -1953 255 -1937 289
rect -1903 255 -1887 289
rect -1953 221 -1887 255
rect -1953 187 -1937 221
rect -1903 187 -1887 221
rect -1953 153 -1887 187
rect -1953 119 -1937 153
rect -1903 119 -1887 153
rect -1953 85 -1887 119
rect -1953 51 -1937 85
rect -1903 51 -1887 85
rect -1953 17 -1887 51
rect -1953 -17 -1937 17
rect -1903 -17 -1887 17
rect -1953 -51 -1887 -17
rect -1953 -85 -1937 -51
rect -1903 -85 -1887 -51
rect -1953 -119 -1887 -85
rect -1953 -153 -1937 -119
rect -1903 -153 -1887 -119
rect -1953 -187 -1887 -153
rect -1953 -221 -1937 -187
rect -1903 -221 -1887 -187
rect -1953 -255 -1887 -221
rect -1953 -289 -1937 -255
rect -1903 -289 -1887 -255
rect -1953 -323 -1887 -289
rect -1953 -357 -1937 -323
rect -1903 -357 -1887 -323
rect -1953 -391 -1887 -357
rect -1953 -425 -1937 -391
rect -1903 -425 -1887 -391
rect -1953 -459 -1887 -425
rect -1953 -493 -1937 -459
rect -1903 -493 -1887 -459
rect -1953 -527 -1887 -493
rect -1953 -561 -1937 -527
rect -1903 -561 -1887 -527
rect -1953 -595 -1887 -561
rect -1953 -629 -1937 -595
rect -1903 -629 -1887 -595
rect -1953 -663 -1887 -629
rect -1953 -697 -1937 -663
rect -1903 -697 -1887 -663
rect -1953 -731 -1887 -697
rect -1953 -765 -1937 -731
rect -1903 -765 -1887 -731
rect -1953 -799 -1887 -765
rect -1953 -833 -1937 -799
rect -1903 -833 -1887 -799
rect -1953 -867 -1887 -833
rect -1953 -901 -1937 -867
rect -1903 -901 -1887 -867
rect -1953 -935 -1887 -901
rect -1953 -969 -1937 -935
rect -1903 -969 -1887 -935
rect -1953 -1000 -1887 -969
rect -1857 969 -1791 1000
rect -1857 935 -1841 969
rect -1807 935 -1791 969
rect -1857 901 -1791 935
rect -1857 867 -1841 901
rect -1807 867 -1791 901
rect -1857 833 -1791 867
rect -1857 799 -1841 833
rect -1807 799 -1791 833
rect -1857 765 -1791 799
rect -1857 731 -1841 765
rect -1807 731 -1791 765
rect -1857 697 -1791 731
rect -1857 663 -1841 697
rect -1807 663 -1791 697
rect -1857 629 -1791 663
rect -1857 595 -1841 629
rect -1807 595 -1791 629
rect -1857 561 -1791 595
rect -1857 527 -1841 561
rect -1807 527 -1791 561
rect -1857 493 -1791 527
rect -1857 459 -1841 493
rect -1807 459 -1791 493
rect -1857 425 -1791 459
rect -1857 391 -1841 425
rect -1807 391 -1791 425
rect -1857 357 -1791 391
rect -1857 323 -1841 357
rect -1807 323 -1791 357
rect -1857 289 -1791 323
rect -1857 255 -1841 289
rect -1807 255 -1791 289
rect -1857 221 -1791 255
rect -1857 187 -1841 221
rect -1807 187 -1791 221
rect -1857 153 -1791 187
rect -1857 119 -1841 153
rect -1807 119 -1791 153
rect -1857 85 -1791 119
rect -1857 51 -1841 85
rect -1807 51 -1791 85
rect -1857 17 -1791 51
rect -1857 -17 -1841 17
rect -1807 -17 -1791 17
rect -1857 -51 -1791 -17
rect -1857 -85 -1841 -51
rect -1807 -85 -1791 -51
rect -1857 -119 -1791 -85
rect -1857 -153 -1841 -119
rect -1807 -153 -1791 -119
rect -1857 -187 -1791 -153
rect -1857 -221 -1841 -187
rect -1807 -221 -1791 -187
rect -1857 -255 -1791 -221
rect -1857 -289 -1841 -255
rect -1807 -289 -1791 -255
rect -1857 -323 -1791 -289
rect -1857 -357 -1841 -323
rect -1807 -357 -1791 -323
rect -1857 -391 -1791 -357
rect -1857 -425 -1841 -391
rect -1807 -425 -1791 -391
rect -1857 -459 -1791 -425
rect -1857 -493 -1841 -459
rect -1807 -493 -1791 -459
rect -1857 -527 -1791 -493
rect -1857 -561 -1841 -527
rect -1807 -561 -1791 -527
rect -1857 -595 -1791 -561
rect -1857 -629 -1841 -595
rect -1807 -629 -1791 -595
rect -1857 -663 -1791 -629
rect -1857 -697 -1841 -663
rect -1807 -697 -1791 -663
rect -1857 -731 -1791 -697
rect -1857 -765 -1841 -731
rect -1807 -765 -1791 -731
rect -1857 -799 -1791 -765
rect -1857 -833 -1841 -799
rect -1807 -833 -1791 -799
rect -1857 -867 -1791 -833
rect -1857 -901 -1841 -867
rect -1807 -901 -1791 -867
rect -1857 -935 -1791 -901
rect -1857 -969 -1841 -935
rect -1807 -969 -1791 -935
rect -1857 -1000 -1791 -969
rect -1761 969 -1695 1000
rect -1761 935 -1745 969
rect -1711 935 -1695 969
rect -1761 901 -1695 935
rect -1761 867 -1745 901
rect -1711 867 -1695 901
rect -1761 833 -1695 867
rect -1761 799 -1745 833
rect -1711 799 -1695 833
rect -1761 765 -1695 799
rect -1761 731 -1745 765
rect -1711 731 -1695 765
rect -1761 697 -1695 731
rect -1761 663 -1745 697
rect -1711 663 -1695 697
rect -1761 629 -1695 663
rect -1761 595 -1745 629
rect -1711 595 -1695 629
rect -1761 561 -1695 595
rect -1761 527 -1745 561
rect -1711 527 -1695 561
rect -1761 493 -1695 527
rect -1761 459 -1745 493
rect -1711 459 -1695 493
rect -1761 425 -1695 459
rect -1761 391 -1745 425
rect -1711 391 -1695 425
rect -1761 357 -1695 391
rect -1761 323 -1745 357
rect -1711 323 -1695 357
rect -1761 289 -1695 323
rect -1761 255 -1745 289
rect -1711 255 -1695 289
rect -1761 221 -1695 255
rect -1761 187 -1745 221
rect -1711 187 -1695 221
rect -1761 153 -1695 187
rect -1761 119 -1745 153
rect -1711 119 -1695 153
rect -1761 85 -1695 119
rect -1761 51 -1745 85
rect -1711 51 -1695 85
rect -1761 17 -1695 51
rect -1761 -17 -1745 17
rect -1711 -17 -1695 17
rect -1761 -51 -1695 -17
rect -1761 -85 -1745 -51
rect -1711 -85 -1695 -51
rect -1761 -119 -1695 -85
rect -1761 -153 -1745 -119
rect -1711 -153 -1695 -119
rect -1761 -187 -1695 -153
rect -1761 -221 -1745 -187
rect -1711 -221 -1695 -187
rect -1761 -255 -1695 -221
rect -1761 -289 -1745 -255
rect -1711 -289 -1695 -255
rect -1761 -323 -1695 -289
rect -1761 -357 -1745 -323
rect -1711 -357 -1695 -323
rect -1761 -391 -1695 -357
rect -1761 -425 -1745 -391
rect -1711 -425 -1695 -391
rect -1761 -459 -1695 -425
rect -1761 -493 -1745 -459
rect -1711 -493 -1695 -459
rect -1761 -527 -1695 -493
rect -1761 -561 -1745 -527
rect -1711 -561 -1695 -527
rect -1761 -595 -1695 -561
rect -1761 -629 -1745 -595
rect -1711 -629 -1695 -595
rect -1761 -663 -1695 -629
rect -1761 -697 -1745 -663
rect -1711 -697 -1695 -663
rect -1761 -731 -1695 -697
rect -1761 -765 -1745 -731
rect -1711 -765 -1695 -731
rect -1761 -799 -1695 -765
rect -1761 -833 -1745 -799
rect -1711 -833 -1695 -799
rect -1761 -867 -1695 -833
rect -1761 -901 -1745 -867
rect -1711 -901 -1695 -867
rect -1761 -935 -1695 -901
rect -1761 -969 -1745 -935
rect -1711 -969 -1695 -935
rect -1761 -1000 -1695 -969
rect -1665 969 -1599 1000
rect -1665 935 -1649 969
rect -1615 935 -1599 969
rect -1665 901 -1599 935
rect -1665 867 -1649 901
rect -1615 867 -1599 901
rect -1665 833 -1599 867
rect -1665 799 -1649 833
rect -1615 799 -1599 833
rect -1665 765 -1599 799
rect -1665 731 -1649 765
rect -1615 731 -1599 765
rect -1665 697 -1599 731
rect -1665 663 -1649 697
rect -1615 663 -1599 697
rect -1665 629 -1599 663
rect -1665 595 -1649 629
rect -1615 595 -1599 629
rect -1665 561 -1599 595
rect -1665 527 -1649 561
rect -1615 527 -1599 561
rect -1665 493 -1599 527
rect -1665 459 -1649 493
rect -1615 459 -1599 493
rect -1665 425 -1599 459
rect -1665 391 -1649 425
rect -1615 391 -1599 425
rect -1665 357 -1599 391
rect -1665 323 -1649 357
rect -1615 323 -1599 357
rect -1665 289 -1599 323
rect -1665 255 -1649 289
rect -1615 255 -1599 289
rect -1665 221 -1599 255
rect -1665 187 -1649 221
rect -1615 187 -1599 221
rect -1665 153 -1599 187
rect -1665 119 -1649 153
rect -1615 119 -1599 153
rect -1665 85 -1599 119
rect -1665 51 -1649 85
rect -1615 51 -1599 85
rect -1665 17 -1599 51
rect -1665 -17 -1649 17
rect -1615 -17 -1599 17
rect -1665 -51 -1599 -17
rect -1665 -85 -1649 -51
rect -1615 -85 -1599 -51
rect -1665 -119 -1599 -85
rect -1665 -153 -1649 -119
rect -1615 -153 -1599 -119
rect -1665 -187 -1599 -153
rect -1665 -221 -1649 -187
rect -1615 -221 -1599 -187
rect -1665 -255 -1599 -221
rect -1665 -289 -1649 -255
rect -1615 -289 -1599 -255
rect -1665 -323 -1599 -289
rect -1665 -357 -1649 -323
rect -1615 -357 -1599 -323
rect -1665 -391 -1599 -357
rect -1665 -425 -1649 -391
rect -1615 -425 -1599 -391
rect -1665 -459 -1599 -425
rect -1665 -493 -1649 -459
rect -1615 -493 -1599 -459
rect -1665 -527 -1599 -493
rect -1665 -561 -1649 -527
rect -1615 -561 -1599 -527
rect -1665 -595 -1599 -561
rect -1665 -629 -1649 -595
rect -1615 -629 -1599 -595
rect -1665 -663 -1599 -629
rect -1665 -697 -1649 -663
rect -1615 -697 -1599 -663
rect -1665 -731 -1599 -697
rect -1665 -765 -1649 -731
rect -1615 -765 -1599 -731
rect -1665 -799 -1599 -765
rect -1665 -833 -1649 -799
rect -1615 -833 -1599 -799
rect -1665 -867 -1599 -833
rect -1665 -901 -1649 -867
rect -1615 -901 -1599 -867
rect -1665 -935 -1599 -901
rect -1665 -969 -1649 -935
rect -1615 -969 -1599 -935
rect -1665 -1000 -1599 -969
rect -1569 969 -1503 1000
rect -1569 935 -1553 969
rect -1519 935 -1503 969
rect -1569 901 -1503 935
rect -1569 867 -1553 901
rect -1519 867 -1503 901
rect -1569 833 -1503 867
rect -1569 799 -1553 833
rect -1519 799 -1503 833
rect -1569 765 -1503 799
rect -1569 731 -1553 765
rect -1519 731 -1503 765
rect -1569 697 -1503 731
rect -1569 663 -1553 697
rect -1519 663 -1503 697
rect -1569 629 -1503 663
rect -1569 595 -1553 629
rect -1519 595 -1503 629
rect -1569 561 -1503 595
rect -1569 527 -1553 561
rect -1519 527 -1503 561
rect -1569 493 -1503 527
rect -1569 459 -1553 493
rect -1519 459 -1503 493
rect -1569 425 -1503 459
rect -1569 391 -1553 425
rect -1519 391 -1503 425
rect -1569 357 -1503 391
rect -1569 323 -1553 357
rect -1519 323 -1503 357
rect -1569 289 -1503 323
rect -1569 255 -1553 289
rect -1519 255 -1503 289
rect -1569 221 -1503 255
rect -1569 187 -1553 221
rect -1519 187 -1503 221
rect -1569 153 -1503 187
rect -1569 119 -1553 153
rect -1519 119 -1503 153
rect -1569 85 -1503 119
rect -1569 51 -1553 85
rect -1519 51 -1503 85
rect -1569 17 -1503 51
rect -1569 -17 -1553 17
rect -1519 -17 -1503 17
rect -1569 -51 -1503 -17
rect -1569 -85 -1553 -51
rect -1519 -85 -1503 -51
rect -1569 -119 -1503 -85
rect -1569 -153 -1553 -119
rect -1519 -153 -1503 -119
rect -1569 -187 -1503 -153
rect -1569 -221 -1553 -187
rect -1519 -221 -1503 -187
rect -1569 -255 -1503 -221
rect -1569 -289 -1553 -255
rect -1519 -289 -1503 -255
rect -1569 -323 -1503 -289
rect -1569 -357 -1553 -323
rect -1519 -357 -1503 -323
rect -1569 -391 -1503 -357
rect -1569 -425 -1553 -391
rect -1519 -425 -1503 -391
rect -1569 -459 -1503 -425
rect -1569 -493 -1553 -459
rect -1519 -493 -1503 -459
rect -1569 -527 -1503 -493
rect -1569 -561 -1553 -527
rect -1519 -561 -1503 -527
rect -1569 -595 -1503 -561
rect -1569 -629 -1553 -595
rect -1519 -629 -1503 -595
rect -1569 -663 -1503 -629
rect -1569 -697 -1553 -663
rect -1519 -697 -1503 -663
rect -1569 -731 -1503 -697
rect -1569 -765 -1553 -731
rect -1519 -765 -1503 -731
rect -1569 -799 -1503 -765
rect -1569 -833 -1553 -799
rect -1519 -833 -1503 -799
rect -1569 -867 -1503 -833
rect -1569 -901 -1553 -867
rect -1519 -901 -1503 -867
rect -1569 -935 -1503 -901
rect -1569 -969 -1553 -935
rect -1519 -969 -1503 -935
rect -1569 -1000 -1503 -969
rect -1473 969 -1407 1000
rect -1473 935 -1457 969
rect -1423 935 -1407 969
rect -1473 901 -1407 935
rect -1473 867 -1457 901
rect -1423 867 -1407 901
rect -1473 833 -1407 867
rect -1473 799 -1457 833
rect -1423 799 -1407 833
rect -1473 765 -1407 799
rect -1473 731 -1457 765
rect -1423 731 -1407 765
rect -1473 697 -1407 731
rect -1473 663 -1457 697
rect -1423 663 -1407 697
rect -1473 629 -1407 663
rect -1473 595 -1457 629
rect -1423 595 -1407 629
rect -1473 561 -1407 595
rect -1473 527 -1457 561
rect -1423 527 -1407 561
rect -1473 493 -1407 527
rect -1473 459 -1457 493
rect -1423 459 -1407 493
rect -1473 425 -1407 459
rect -1473 391 -1457 425
rect -1423 391 -1407 425
rect -1473 357 -1407 391
rect -1473 323 -1457 357
rect -1423 323 -1407 357
rect -1473 289 -1407 323
rect -1473 255 -1457 289
rect -1423 255 -1407 289
rect -1473 221 -1407 255
rect -1473 187 -1457 221
rect -1423 187 -1407 221
rect -1473 153 -1407 187
rect -1473 119 -1457 153
rect -1423 119 -1407 153
rect -1473 85 -1407 119
rect -1473 51 -1457 85
rect -1423 51 -1407 85
rect -1473 17 -1407 51
rect -1473 -17 -1457 17
rect -1423 -17 -1407 17
rect -1473 -51 -1407 -17
rect -1473 -85 -1457 -51
rect -1423 -85 -1407 -51
rect -1473 -119 -1407 -85
rect -1473 -153 -1457 -119
rect -1423 -153 -1407 -119
rect -1473 -187 -1407 -153
rect -1473 -221 -1457 -187
rect -1423 -221 -1407 -187
rect -1473 -255 -1407 -221
rect -1473 -289 -1457 -255
rect -1423 -289 -1407 -255
rect -1473 -323 -1407 -289
rect -1473 -357 -1457 -323
rect -1423 -357 -1407 -323
rect -1473 -391 -1407 -357
rect -1473 -425 -1457 -391
rect -1423 -425 -1407 -391
rect -1473 -459 -1407 -425
rect -1473 -493 -1457 -459
rect -1423 -493 -1407 -459
rect -1473 -527 -1407 -493
rect -1473 -561 -1457 -527
rect -1423 -561 -1407 -527
rect -1473 -595 -1407 -561
rect -1473 -629 -1457 -595
rect -1423 -629 -1407 -595
rect -1473 -663 -1407 -629
rect -1473 -697 -1457 -663
rect -1423 -697 -1407 -663
rect -1473 -731 -1407 -697
rect -1473 -765 -1457 -731
rect -1423 -765 -1407 -731
rect -1473 -799 -1407 -765
rect -1473 -833 -1457 -799
rect -1423 -833 -1407 -799
rect -1473 -867 -1407 -833
rect -1473 -901 -1457 -867
rect -1423 -901 -1407 -867
rect -1473 -935 -1407 -901
rect -1473 -969 -1457 -935
rect -1423 -969 -1407 -935
rect -1473 -1000 -1407 -969
rect -1377 969 -1311 1000
rect -1377 935 -1361 969
rect -1327 935 -1311 969
rect -1377 901 -1311 935
rect -1377 867 -1361 901
rect -1327 867 -1311 901
rect -1377 833 -1311 867
rect -1377 799 -1361 833
rect -1327 799 -1311 833
rect -1377 765 -1311 799
rect -1377 731 -1361 765
rect -1327 731 -1311 765
rect -1377 697 -1311 731
rect -1377 663 -1361 697
rect -1327 663 -1311 697
rect -1377 629 -1311 663
rect -1377 595 -1361 629
rect -1327 595 -1311 629
rect -1377 561 -1311 595
rect -1377 527 -1361 561
rect -1327 527 -1311 561
rect -1377 493 -1311 527
rect -1377 459 -1361 493
rect -1327 459 -1311 493
rect -1377 425 -1311 459
rect -1377 391 -1361 425
rect -1327 391 -1311 425
rect -1377 357 -1311 391
rect -1377 323 -1361 357
rect -1327 323 -1311 357
rect -1377 289 -1311 323
rect -1377 255 -1361 289
rect -1327 255 -1311 289
rect -1377 221 -1311 255
rect -1377 187 -1361 221
rect -1327 187 -1311 221
rect -1377 153 -1311 187
rect -1377 119 -1361 153
rect -1327 119 -1311 153
rect -1377 85 -1311 119
rect -1377 51 -1361 85
rect -1327 51 -1311 85
rect -1377 17 -1311 51
rect -1377 -17 -1361 17
rect -1327 -17 -1311 17
rect -1377 -51 -1311 -17
rect -1377 -85 -1361 -51
rect -1327 -85 -1311 -51
rect -1377 -119 -1311 -85
rect -1377 -153 -1361 -119
rect -1327 -153 -1311 -119
rect -1377 -187 -1311 -153
rect -1377 -221 -1361 -187
rect -1327 -221 -1311 -187
rect -1377 -255 -1311 -221
rect -1377 -289 -1361 -255
rect -1327 -289 -1311 -255
rect -1377 -323 -1311 -289
rect -1377 -357 -1361 -323
rect -1327 -357 -1311 -323
rect -1377 -391 -1311 -357
rect -1377 -425 -1361 -391
rect -1327 -425 -1311 -391
rect -1377 -459 -1311 -425
rect -1377 -493 -1361 -459
rect -1327 -493 -1311 -459
rect -1377 -527 -1311 -493
rect -1377 -561 -1361 -527
rect -1327 -561 -1311 -527
rect -1377 -595 -1311 -561
rect -1377 -629 -1361 -595
rect -1327 -629 -1311 -595
rect -1377 -663 -1311 -629
rect -1377 -697 -1361 -663
rect -1327 -697 -1311 -663
rect -1377 -731 -1311 -697
rect -1377 -765 -1361 -731
rect -1327 -765 -1311 -731
rect -1377 -799 -1311 -765
rect -1377 -833 -1361 -799
rect -1327 -833 -1311 -799
rect -1377 -867 -1311 -833
rect -1377 -901 -1361 -867
rect -1327 -901 -1311 -867
rect -1377 -935 -1311 -901
rect -1377 -969 -1361 -935
rect -1327 -969 -1311 -935
rect -1377 -1000 -1311 -969
rect -1281 969 -1215 1000
rect -1281 935 -1265 969
rect -1231 935 -1215 969
rect -1281 901 -1215 935
rect -1281 867 -1265 901
rect -1231 867 -1215 901
rect -1281 833 -1215 867
rect -1281 799 -1265 833
rect -1231 799 -1215 833
rect -1281 765 -1215 799
rect -1281 731 -1265 765
rect -1231 731 -1215 765
rect -1281 697 -1215 731
rect -1281 663 -1265 697
rect -1231 663 -1215 697
rect -1281 629 -1215 663
rect -1281 595 -1265 629
rect -1231 595 -1215 629
rect -1281 561 -1215 595
rect -1281 527 -1265 561
rect -1231 527 -1215 561
rect -1281 493 -1215 527
rect -1281 459 -1265 493
rect -1231 459 -1215 493
rect -1281 425 -1215 459
rect -1281 391 -1265 425
rect -1231 391 -1215 425
rect -1281 357 -1215 391
rect -1281 323 -1265 357
rect -1231 323 -1215 357
rect -1281 289 -1215 323
rect -1281 255 -1265 289
rect -1231 255 -1215 289
rect -1281 221 -1215 255
rect -1281 187 -1265 221
rect -1231 187 -1215 221
rect -1281 153 -1215 187
rect -1281 119 -1265 153
rect -1231 119 -1215 153
rect -1281 85 -1215 119
rect -1281 51 -1265 85
rect -1231 51 -1215 85
rect -1281 17 -1215 51
rect -1281 -17 -1265 17
rect -1231 -17 -1215 17
rect -1281 -51 -1215 -17
rect -1281 -85 -1265 -51
rect -1231 -85 -1215 -51
rect -1281 -119 -1215 -85
rect -1281 -153 -1265 -119
rect -1231 -153 -1215 -119
rect -1281 -187 -1215 -153
rect -1281 -221 -1265 -187
rect -1231 -221 -1215 -187
rect -1281 -255 -1215 -221
rect -1281 -289 -1265 -255
rect -1231 -289 -1215 -255
rect -1281 -323 -1215 -289
rect -1281 -357 -1265 -323
rect -1231 -357 -1215 -323
rect -1281 -391 -1215 -357
rect -1281 -425 -1265 -391
rect -1231 -425 -1215 -391
rect -1281 -459 -1215 -425
rect -1281 -493 -1265 -459
rect -1231 -493 -1215 -459
rect -1281 -527 -1215 -493
rect -1281 -561 -1265 -527
rect -1231 -561 -1215 -527
rect -1281 -595 -1215 -561
rect -1281 -629 -1265 -595
rect -1231 -629 -1215 -595
rect -1281 -663 -1215 -629
rect -1281 -697 -1265 -663
rect -1231 -697 -1215 -663
rect -1281 -731 -1215 -697
rect -1281 -765 -1265 -731
rect -1231 -765 -1215 -731
rect -1281 -799 -1215 -765
rect -1281 -833 -1265 -799
rect -1231 -833 -1215 -799
rect -1281 -867 -1215 -833
rect -1281 -901 -1265 -867
rect -1231 -901 -1215 -867
rect -1281 -935 -1215 -901
rect -1281 -969 -1265 -935
rect -1231 -969 -1215 -935
rect -1281 -1000 -1215 -969
rect -1185 969 -1119 1000
rect -1185 935 -1169 969
rect -1135 935 -1119 969
rect -1185 901 -1119 935
rect -1185 867 -1169 901
rect -1135 867 -1119 901
rect -1185 833 -1119 867
rect -1185 799 -1169 833
rect -1135 799 -1119 833
rect -1185 765 -1119 799
rect -1185 731 -1169 765
rect -1135 731 -1119 765
rect -1185 697 -1119 731
rect -1185 663 -1169 697
rect -1135 663 -1119 697
rect -1185 629 -1119 663
rect -1185 595 -1169 629
rect -1135 595 -1119 629
rect -1185 561 -1119 595
rect -1185 527 -1169 561
rect -1135 527 -1119 561
rect -1185 493 -1119 527
rect -1185 459 -1169 493
rect -1135 459 -1119 493
rect -1185 425 -1119 459
rect -1185 391 -1169 425
rect -1135 391 -1119 425
rect -1185 357 -1119 391
rect -1185 323 -1169 357
rect -1135 323 -1119 357
rect -1185 289 -1119 323
rect -1185 255 -1169 289
rect -1135 255 -1119 289
rect -1185 221 -1119 255
rect -1185 187 -1169 221
rect -1135 187 -1119 221
rect -1185 153 -1119 187
rect -1185 119 -1169 153
rect -1135 119 -1119 153
rect -1185 85 -1119 119
rect -1185 51 -1169 85
rect -1135 51 -1119 85
rect -1185 17 -1119 51
rect -1185 -17 -1169 17
rect -1135 -17 -1119 17
rect -1185 -51 -1119 -17
rect -1185 -85 -1169 -51
rect -1135 -85 -1119 -51
rect -1185 -119 -1119 -85
rect -1185 -153 -1169 -119
rect -1135 -153 -1119 -119
rect -1185 -187 -1119 -153
rect -1185 -221 -1169 -187
rect -1135 -221 -1119 -187
rect -1185 -255 -1119 -221
rect -1185 -289 -1169 -255
rect -1135 -289 -1119 -255
rect -1185 -323 -1119 -289
rect -1185 -357 -1169 -323
rect -1135 -357 -1119 -323
rect -1185 -391 -1119 -357
rect -1185 -425 -1169 -391
rect -1135 -425 -1119 -391
rect -1185 -459 -1119 -425
rect -1185 -493 -1169 -459
rect -1135 -493 -1119 -459
rect -1185 -527 -1119 -493
rect -1185 -561 -1169 -527
rect -1135 -561 -1119 -527
rect -1185 -595 -1119 -561
rect -1185 -629 -1169 -595
rect -1135 -629 -1119 -595
rect -1185 -663 -1119 -629
rect -1185 -697 -1169 -663
rect -1135 -697 -1119 -663
rect -1185 -731 -1119 -697
rect -1185 -765 -1169 -731
rect -1135 -765 -1119 -731
rect -1185 -799 -1119 -765
rect -1185 -833 -1169 -799
rect -1135 -833 -1119 -799
rect -1185 -867 -1119 -833
rect -1185 -901 -1169 -867
rect -1135 -901 -1119 -867
rect -1185 -935 -1119 -901
rect -1185 -969 -1169 -935
rect -1135 -969 -1119 -935
rect -1185 -1000 -1119 -969
rect -1089 969 -1023 1000
rect -1089 935 -1073 969
rect -1039 935 -1023 969
rect -1089 901 -1023 935
rect -1089 867 -1073 901
rect -1039 867 -1023 901
rect -1089 833 -1023 867
rect -1089 799 -1073 833
rect -1039 799 -1023 833
rect -1089 765 -1023 799
rect -1089 731 -1073 765
rect -1039 731 -1023 765
rect -1089 697 -1023 731
rect -1089 663 -1073 697
rect -1039 663 -1023 697
rect -1089 629 -1023 663
rect -1089 595 -1073 629
rect -1039 595 -1023 629
rect -1089 561 -1023 595
rect -1089 527 -1073 561
rect -1039 527 -1023 561
rect -1089 493 -1023 527
rect -1089 459 -1073 493
rect -1039 459 -1023 493
rect -1089 425 -1023 459
rect -1089 391 -1073 425
rect -1039 391 -1023 425
rect -1089 357 -1023 391
rect -1089 323 -1073 357
rect -1039 323 -1023 357
rect -1089 289 -1023 323
rect -1089 255 -1073 289
rect -1039 255 -1023 289
rect -1089 221 -1023 255
rect -1089 187 -1073 221
rect -1039 187 -1023 221
rect -1089 153 -1023 187
rect -1089 119 -1073 153
rect -1039 119 -1023 153
rect -1089 85 -1023 119
rect -1089 51 -1073 85
rect -1039 51 -1023 85
rect -1089 17 -1023 51
rect -1089 -17 -1073 17
rect -1039 -17 -1023 17
rect -1089 -51 -1023 -17
rect -1089 -85 -1073 -51
rect -1039 -85 -1023 -51
rect -1089 -119 -1023 -85
rect -1089 -153 -1073 -119
rect -1039 -153 -1023 -119
rect -1089 -187 -1023 -153
rect -1089 -221 -1073 -187
rect -1039 -221 -1023 -187
rect -1089 -255 -1023 -221
rect -1089 -289 -1073 -255
rect -1039 -289 -1023 -255
rect -1089 -323 -1023 -289
rect -1089 -357 -1073 -323
rect -1039 -357 -1023 -323
rect -1089 -391 -1023 -357
rect -1089 -425 -1073 -391
rect -1039 -425 -1023 -391
rect -1089 -459 -1023 -425
rect -1089 -493 -1073 -459
rect -1039 -493 -1023 -459
rect -1089 -527 -1023 -493
rect -1089 -561 -1073 -527
rect -1039 -561 -1023 -527
rect -1089 -595 -1023 -561
rect -1089 -629 -1073 -595
rect -1039 -629 -1023 -595
rect -1089 -663 -1023 -629
rect -1089 -697 -1073 -663
rect -1039 -697 -1023 -663
rect -1089 -731 -1023 -697
rect -1089 -765 -1073 -731
rect -1039 -765 -1023 -731
rect -1089 -799 -1023 -765
rect -1089 -833 -1073 -799
rect -1039 -833 -1023 -799
rect -1089 -867 -1023 -833
rect -1089 -901 -1073 -867
rect -1039 -901 -1023 -867
rect -1089 -935 -1023 -901
rect -1089 -969 -1073 -935
rect -1039 -969 -1023 -935
rect -1089 -1000 -1023 -969
rect -993 969 -927 1000
rect -993 935 -977 969
rect -943 935 -927 969
rect -993 901 -927 935
rect -993 867 -977 901
rect -943 867 -927 901
rect -993 833 -927 867
rect -993 799 -977 833
rect -943 799 -927 833
rect -993 765 -927 799
rect -993 731 -977 765
rect -943 731 -927 765
rect -993 697 -927 731
rect -993 663 -977 697
rect -943 663 -927 697
rect -993 629 -927 663
rect -993 595 -977 629
rect -943 595 -927 629
rect -993 561 -927 595
rect -993 527 -977 561
rect -943 527 -927 561
rect -993 493 -927 527
rect -993 459 -977 493
rect -943 459 -927 493
rect -993 425 -927 459
rect -993 391 -977 425
rect -943 391 -927 425
rect -993 357 -927 391
rect -993 323 -977 357
rect -943 323 -927 357
rect -993 289 -927 323
rect -993 255 -977 289
rect -943 255 -927 289
rect -993 221 -927 255
rect -993 187 -977 221
rect -943 187 -927 221
rect -993 153 -927 187
rect -993 119 -977 153
rect -943 119 -927 153
rect -993 85 -927 119
rect -993 51 -977 85
rect -943 51 -927 85
rect -993 17 -927 51
rect -993 -17 -977 17
rect -943 -17 -927 17
rect -993 -51 -927 -17
rect -993 -85 -977 -51
rect -943 -85 -927 -51
rect -993 -119 -927 -85
rect -993 -153 -977 -119
rect -943 -153 -927 -119
rect -993 -187 -927 -153
rect -993 -221 -977 -187
rect -943 -221 -927 -187
rect -993 -255 -927 -221
rect -993 -289 -977 -255
rect -943 -289 -927 -255
rect -993 -323 -927 -289
rect -993 -357 -977 -323
rect -943 -357 -927 -323
rect -993 -391 -927 -357
rect -993 -425 -977 -391
rect -943 -425 -927 -391
rect -993 -459 -927 -425
rect -993 -493 -977 -459
rect -943 -493 -927 -459
rect -993 -527 -927 -493
rect -993 -561 -977 -527
rect -943 -561 -927 -527
rect -993 -595 -927 -561
rect -993 -629 -977 -595
rect -943 -629 -927 -595
rect -993 -663 -927 -629
rect -993 -697 -977 -663
rect -943 -697 -927 -663
rect -993 -731 -927 -697
rect -993 -765 -977 -731
rect -943 -765 -927 -731
rect -993 -799 -927 -765
rect -993 -833 -977 -799
rect -943 -833 -927 -799
rect -993 -867 -927 -833
rect -993 -901 -977 -867
rect -943 -901 -927 -867
rect -993 -935 -927 -901
rect -993 -969 -977 -935
rect -943 -969 -927 -935
rect -993 -1000 -927 -969
rect -897 969 -831 1000
rect -897 935 -881 969
rect -847 935 -831 969
rect -897 901 -831 935
rect -897 867 -881 901
rect -847 867 -831 901
rect -897 833 -831 867
rect -897 799 -881 833
rect -847 799 -831 833
rect -897 765 -831 799
rect -897 731 -881 765
rect -847 731 -831 765
rect -897 697 -831 731
rect -897 663 -881 697
rect -847 663 -831 697
rect -897 629 -831 663
rect -897 595 -881 629
rect -847 595 -831 629
rect -897 561 -831 595
rect -897 527 -881 561
rect -847 527 -831 561
rect -897 493 -831 527
rect -897 459 -881 493
rect -847 459 -831 493
rect -897 425 -831 459
rect -897 391 -881 425
rect -847 391 -831 425
rect -897 357 -831 391
rect -897 323 -881 357
rect -847 323 -831 357
rect -897 289 -831 323
rect -897 255 -881 289
rect -847 255 -831 289
rect -897 221 -831 255
rect -897 187 -881 221
rect -847 187 -831 221
rect -897 153 -831 187
rect -897 119 -881 153
rect -847 119 -831 153
rect -897 85 -831 119
rect -897 51 -881 85
rect -847 51 -831 85
rect -897 17 -831 51
rect -897 -17 -881 17
rect -847 -17 -831 17
rect -897 -51 -831 -17
rect -897 -85 -881 -51
rect -847 -85 -831 -51
rect -897 -119 -831 -85
rect -897 -153 -881 -119
rect -847 -153 -831 -119
rect -897 -187 -831 -153
rect -897 -221 -881 -187
rect -847 -221 -831 -187
rect -897 -255 -831 -221
rect -897 -289 -881 -255
rect -847 -289 -831 -255
rect -897 -323 -831 -289
rect -897 -357 -881 -323
rect -847 -357 -831 -323
rect -897 -391 -831 -357
rect -897 -425 -881 -391
rect -847 -425 -831 -391
rect -897 -459 -831 -425
rect -897 -493 -881 -459
rect -847 -493 -831 -459
rect -897 -527 -831 -493
rect -897 -561 -881 -527
rect -847 -561 -831 -527
rect -897 -595 -831 -561
rect -897 -629 -881 -595
rect -847 -629 -831 -595
rect -897 -663 -831 -629
rect -897 -697 -881 -663
rect -847 -697 -831 -663
rect -897 -731 -831 -697
rect -897 -765 -881 -731
rect -847 -765 -831 -731
rect -897 -799 -831 -765
rect -897 -833 -881 -799
rect -847 -833 -831 -799
rect -897 -867 -831 -833
rect -897 -901 -881 -867
rect -847 -901 -831 -867
rect -897 -935 -831 -901
rect -897 -969 -881 -935
rect -847 -969 -831 -935
rect -897 -1000 -831 -969
rect -801 969 -735 1000
rect -801 935 -785 969
rect -751 935 -735 969
rect -801 901 -735 935
rect -801 867 -785 901
rect -751 867 -735 901
rect -801 833 -735 867
rect -801 799 -785 833
rect -751 799 -735 833
rect -801 765 -735 799
rect -801 731 -785 765
rect -751 731 -735 765
rect -801 697 -735 731
rect -801 663 -785 697
rect -751 663 -735 697
rect -801 629 -735 663
rect -801 595 -785 629
rect -751 595 -735 629
rect -801 561 -735 595
rect -801 527 -785 561
rect -751 527 -735 561
rect -801 493 -735 527
rect -801 459 -785 493
rect -751 459 -735 493
rect -801 425 -735 459
rect -801 391 -785 425
rect -751 391 -735 425
rect -801 357 -735 391
rect -801 323 -785 357
rect -751 323 -735 357
rect -801 289 -735 323
rect -801 255 -785 289
rect -751 255 -735 289
rect -801 221 -735 255
rect -801 187 -785 221
rect -751 187 -735 221
rect -801 153 -735 187
rect -801 119 -785 153
rect -751 119 -735 153
rect -801 85 -735 119
rect -801 51 -785 85
rect -751 51 -735 85
rect -801 17 -735 51
rect -801 -17 -785 17
rect -751 -17 -735 17
rect -801 -51 -735 -17
rect -801 -85 -785 -51
rect -751 -85 -735 -51
rect -801 -119 -735 -85
rect -801 -153 -785 -119
rect -751 -153 -735 -119
rect -801 -187 -735 -153
rect -801 -221 -785 -187
rect -751 -221 -735 -187
rect -801 -255 -735 -221
rect -801 -289 -785 -255
rect -751 -289 -735 -255
rect -801 -323 -735 -289
rect -801 -357 -785 -323
rect -751 -357 -735 -323
rect -801 -391 -735 -357
rect -801 -425 -785 -391
rect -751 -425 -735 -391
rect -801 -459 -735 -425
rect -801 -493 -785 -459
rect -751 -493 -735 -459
rect -801 -527 -735 -493
rect -801 -561 -785 -527
rect -751 -561 -735 -527
rect -801 -595 -735 -561
rect -801 -629 -785 -595
rect -751 -629 -735 -595
rect -801 -663 -735 -629
rect -801 -697 -785 -663
rect -751 -697 -735 -663
rect -801 -731 -735 -697
rect -801 -765 -785 -731
rect -751 -765 -735 -731
rect -801 -799 -735 -765
rect -801 -833 -785 -799
rect -751 -833 -735 -799
rect -801 -867 -735 -833
rect -801 -901 -785 -867
rect -751 -901 -735 -867
rect -801 -935 -735 -901
rect -801 -969 -785 -935
rect -751 -969 -735 -935
rect -801 -1000 -735 -969
rect -705 969 -639 1000
rect -705 935 -689 969
rect -655 935 -639 969
rect -705 901 -639 935
rect -705 867 -689 901
rect -655 867 -639 901
rect -705 833 -639 867
rect -705 799 -689 833
rect -655 799 -639 833
rect -705 765 -639 799
rect -705 731 -689 765
rect -655 731 -639 765
rect -705 697 -639 731
rect -705 663 -689 697
rect -655 663 -639 697
rect -705 629 -639 663
rect -705 595 -689 629
rect -655 595 -639 629
rect -705 561 -639 595
rect -705 527 -689 561
rect -655 527 -639 561
rect -705 493 -639 527
rect -705 459 -689 493
rect -655 459 -639 493
rect -705 425 -639 459
rect -705 391 -689 425
rect -655 391 -639 425
rect -705 357 -639 391
rect -705 323 -689 357
rect -655 323 -639 357
rect -705 289 -639 323
rect -705 255 -689 289
rect -655 255 -639 289
rect -705 221 -639 255
rect -705 187 -689 221
rect -655 187 -639 221
rect -705 153 -639 187
rect -705 119 -689 153
rect -655 119 -639 153
rect -705 85 -639 119
rect -705 51 -689 85
rect -655 51 -639 85
rect -705 17 -639 51
rect -705 -17 -689 17
rect -655 -17 -639 17
rect -705 -51 -639 -17
rect -705 -85 -689 -51
rect -655 -85 -639 -51
rect -705 -119 -639 -85
rect -705 -153 -689 -119
rect -655 -153 -639 -119
rect -705 -187 -639 -153
rect -705 -221 -689 -187
rect -655 -221 -639 -187
rect -705 -255 -639 -221
rect -705 -289 -689 -255
rect -655 -289 -639 -255
rect -705 -323 -639 -289
rect -705 -357 -689 -323
rect -655 -357 -639 -323
rect -705 -391 -639 -357
rect -705 -425 -689 -391
rect -655 -425 -639 -391
rect -705 -459 -639 -425
rect -705 -493 -689 -459
rect -655 -493 -639 -459
rect -705 -527 -639 -493
rect -705 -561 -689 -527
rect -655 -561 -639 -527
rect -705 -595 -639 -561
rect -705 -629 -689 -595
rect -655 -629 -639 -595
rect -705 -663 -639 -629
rect -705 -697 -689 -663
rect -655 -697 -639 -663
rect -705 -731 -639 -697
rect -705 -765 -689 -731
rect -655 -765 -639 -731
rect -705 -799 -639 -765
rect -705 -833 -689 -799
rect -655 -833 -639 -799
rect -705 -867 -639 -833
rect -705 -901 -689 -867
rect -655 -901 -639 -867
rect -705 -935 -639 -901
rect -705 -969 -689 -935
rect -655 -969 -639 -935
rect -705 -1000 -639 -969
rect -609 969 -543 1000
rect -609 935 -593 969
rect -559 935 -543 969
rect -609 901 -543 935
rect -609 867 -593 901
rect -559 867 -543 901
rect -609 833 -543 867
rect -609 799 -593 833
rect -559 799 -543 833
rect -609 765 -543 799
rect -609 731 -593 765
rect -559 731 -543 765
rect -609 697 -543 731
rect -609 663 -593 697
rect -559 663 -543 697
rect -609 629 -543 663
rect -609 595 -593 629
rect -559 595 -543 629
rect -609 561 -543 595
rect -609 527 -593 561
rect -559 527 -543 561
rect -609 493 -543 527
rect -609 459 -593 493
rect -559 459 -543 493
rect -609 425 -543 459
rect -609 391 -593 425
rect -559 391 -543 425
rect -609 357 -543 391
rect -609 323 -593 357
rect -559 323 -543 357
rect -609 289 -543 323
rect -609 255 -593 289
rect -559 255 -543 289
rect -609 221 -543 255
rect -609 187 -593 221
rect -559 187 -543 221
rect -609 153 -543 187
rect -609 119 -593 153
rect -559 119 -543 153
rect -609 85 -543 119
rect -609 51 -593 85
rect -559 51 -543 85
rect -609 17 -543 51
rect -609 -17 -593 17
rect -559 -17 -543 17
rect -609 -51 -543 -17
rect -609 -85 -593 -51
rect -559 -85 -543 -51
rect -609 -119 -543 -85
rect -609 -153 -593 -119
rect -559 -153 -543 -119
rect -609 -187 -543 -153
rect -609 -221 -593 -187
rect -559 -221 -543 -187
rect -609 -255 -543 -221
rect -609 -289 -593 -255
rect -559 -289 -543 -255
rect -609 -323 -543 -289
rect -609 -357 -593 -323
rect -559 -357 -543 -323
rect -609 -391 -543 -357
rect -609 -425 -593 -391
rect -559 -425 -543 -391
rect -609 -459 -543 -425
rect -609 -493 -593 -459
rect -559 -493 -543 -459
rect -609 -527 -543 -493
rect -609 -561 -593 -527
rect -559 -561 -543 -527
rect -609 -595 -543 -561
rect -609 -629 -593 -595
rect -559 -629 -543 -595
rect -609 -663 -543 -629
rect -609 -697 -593 -663
rect -559 -697 -543 -663
rect -609 -731 -543 -697
rect -609 -765 -593 -731
rect -559 -765 -543 -731
rect -609 -799 -543 -765
rect -609 -833 -593 -799
rect -559 -833 -543 -799
rect -609 -867 -543 -833
rect -609 -901 -593 -867
rect -559 -901 -543 -867
rect -609 -935 -543 -901
rect -609 -969 -593 -935
rect -559 -969 -543 -935
rect -609 -1000 -543 -969
rect -513 969 -447 1000
rect -513 935 -497 969
rect -463 935 -447 969
rect -513 901 -447 935
rect -513 867 -497 901
rect -463 867 -447 901
rect -513 833 -447 867
rect -513 799 -497 833
rect -463 799 -447 833
rect -513 765 -447 799
rect -513 731 -497 765
rect -463 731 -447 765
rect -513 697 -447 731
rect -513 663 -497 697
rect -463 663 -447 697
rect -513 629 -447 663
rect -513 595 -497 629
rect -463 595 -447 629
rect -513 561 -447 595
rect -513 527 -497 561
rect -463 527 -447 561
rect -513 493 -447 527
rect -513 459 -497 493
rect -463 459 -447 493
rect -513 425 -447 459
rect -513 391 -497 425
rect -463 391 -447 425
rect -513 357 -447 391
rect -513 323 -497 357
rect -463 323 -447 357
rect -513 289 -447 323
rect -513 255 -497 289
rect -463 255 -447 289
rect -513 221 -447 255
rect -513 187 -497 221
rect -463 187 -447 221
rect -513 153 -447 187
rect -513 119 -497 153
rect -463 119 -447 153
rect -513 85 -447 119
rect -513 51 -497 85
rect -463 51 -447 85
rect -513 17 -447 51
rect -513 -17 -497 17
rect -463 -17 -447 17
rect -513 -51 -447 -17
rect -513 -85 -497 -51
rect -463 -85 -447 -51
rect -513 -119 -447 -85
rect -513 -153 -497 -119
rect -463 -153 -447 -119
rect -513 -187 -447 -153
rect -513 -221 -497 -187
rect -463 -221 -447 -187
rect -513 -255 -447 -221
rect -513 -289 -497 -255
rect -463 -289 -447 -255
rect -513 -323 -447 -289
rect -513 -357 -497 -323
rect -463 -357 -447 -323
rect -513 -391 -447 -357
rect -513 -425 -497 -391
rect -463 -425 -447 -391
rect -513 -459 -447 -425
rect -513 -493 -497 -459
rect -463 -493 -447 -459
rect -513 -527 -447 -493
rect -513 -561 -497 -527
rect -463 -561 -447 -527
rect -513 -595 -447 -561
rect -513 -629 -497 -595
rect -463 -629 -447 -595
rect -513 -663 -447 -629
rect -513 -697 -497 -663
rect -463 -697 -447 -663
rect -513 -731 -447 -697
rect -513 -765 -497 -731
rect -463 -765 -447 -731
rect -513 -799 -447 -765
rect -513 -833 -497 -799
rect -463 -833 -447 -799
rect -513 -867 -447 -833
rect -513 -901 -497 -867
rect -463 -901 -447 -867
rect -513 -935 -447 -901
rect -513 -969 -497 -935
rect -463 -969 -447 -935
rect -513 -1000 -447 -969
rect -417 969 -351 1000
rect -417 935 -401 969
rect -367 935 -351 969
rect -417 901 -351 935
rect -417 867 -401 901
rect -367 867 -351 901
rect -417 833 -351 867
rect -417 799 -401 833
rect -367 799 -351 833
rect -417 765 -351 799
rect -417 731 -401 765
rect -367 731 -351 765
rect -417 697 -351 731
rect -417 663 -401 697
rect -367 663 -351 697
rect -417 629 -351 663
rect -417 595 -401 629
rect -367 595 -351 629
rect -417 561 -351 595
rect -417 527 -401 561
rect -367 527 -351 561
rect -417 493 -351 527
rect -417 459 -401 493
rect -367 459 -351 493
rect -417 425 -351 459
rect -417 391 -401 425
rect -367 391 -351 425
rect -417 357 -351 391
rect -417 323 -401 357
rect -367 323 -351 357
rect -417 289 -351 323
rect -417 255 -401 289
rect -367 255 -351 289
rect -417 221 -351 255
rect -417 187 -401 221
rect -367 187 -351 221
rect -417 153 -351 187
rect -417 119 -401 153
rect -367 119 -351 153
rect -417 85 -351 119
rect -417 51 -401 85
rect -367 51 -351 85
rect -417 17 -351 51
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -51 -351 -17
rect -417 -85 -401 -51
rect -367 -85 -351 -51
rect -417 -119 -351 -85
rect -417 -153 -401 -119
rect -367 -153 -351 -119
rect -417 -187 -351 -153
rect -417 -221 -401 -187
rect -367 -221 -351 -187
rect -417 -255 -351 -221
rect -417 -289 -401 -255
rect -367 -289 -351 -255
rect -417 -323 -351 -289
rect -417 -357 -401 -323
rect -367 -357 -351 -323
rect -417 -391 -351 -357
rect -417 -425 -401 -391
rect -367 -425 -351 -391
rect -417 -459 -351 -425
rect -417 -493 -401 -459
rect -367 -493 -351 -459
rect -417 -527 -351 -493
rect -417 -561 -401 -527
rect -367 -561 -351 -527
rect -417 -595 -351 -561
rect -417 -629 -401 -595
rect -367 -629 -351 -595
rect -417 -663 -351 -629
rect -417 -697 -401 -663
rect -367 -697 -351 -663
rect -417 -731 -351 -697
rect -417 -765 -401 -731
rect -367 -765 -351 -731
rect -417 -799 -351 -765
rect -417 -833 -401 -799
rect -367 -833 -351 -799
rect -417 -867 -351 -833
rect -417 -901 -401 -867
rect -367 -901 -351 -867
rect -417 -935 -351 -901
rect -417 -969 -401 -935
rect -367 -969 -351 -935
rect -417 -1000 -351 -969
rect -321 969 -255 1000
rect -321 935 -305 969
rect -271 935 -255 969
rect -321 901 -255 935
rect -321 867 -305 901
rect -271 867 -255 901
rect -321 833 -255 867
rect -321 799 -305 833
rect -271 799 -255 833
rect -321 765 -255 799
rect -321 731 -305 765
rect -271 731 -255 765
rect -321 697 -255 731
rect -321 663 -305 697
rect -271 663 -255 697
rect -321 629 -255 663
rect -321 595 -305 629
rect -271 595 -255 629
rect -321 561 -255 595
rect -321 527 -305 561
rect -271 527 -255 561
rect -321 493 -255 527
rect -321 459 -305 493
rect -271 459 -255 493
rect -321 425 -255 459
rect -321 391 -305 425
rect -271 391 -255 425
rect -321 357 -255 391
rect -321 323 -305 357
rect -271 323 -255 357
rect -321 289 -255 323
rect -321 255 -305 289
rect -271 255 -255 289
rect -321 221 -255 255
rect -321 187 -305 221
rect -271 187 -255 221
rect -321 153 -255 187
rect -321 119 -305 153
rect -271 119 -255 153
rect -321 85 -255 119
rect -321 51 -305 85
rect -271 51 -255 85
rect -321 17 -255 51
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -51 -255 -17
rect -321 -85 -305 -51
rect -271 -85 -255 -51
rect -321 -119 -255 -85
rect -321 -153 -305 -119
rect -271 -153 -255 -119
rect -321 -187 -255 -153
rect -321 -221 -305 -187
rect -271 -221 -255 -187
rect -321 -255 -255 -221
rect -321 -289 -305 -255
rect -271 -289 -255 -255
rect -321 -323 -255 -289
rect -321 -357 -305 -323
rect -271 -357 -255 -323
rect -321 -391 -255 -357
rect -321 -425 -305 -391
rect -271 -425 -255 -391
rect -321 -459 -255 -425
rect -321 -493 -305 -459
rect -271 -493 -255 -459
rect -321 -527 -255 -493
rect -321 -561 -305 -527
rect -271 -561 -255 -527
rect -321 -595 -255 -561
rect -321 -629 -305 -595
rect -271 -629 -255 -595
rect -321 -663 -255 -629
rect -321 -697 -305 -663
rect -271 -697 -255 -663
rect -321 -731 -255 -697
rect -321 -765 -305 -731
rect -271 -765 -255 -731
rect -321 -799 -255 -765
rect -321 -833 -305 -799
rect -271 -833 -255 -799
rect -321 -867 -255 -833
rect -321 -901 -305 -867
rect -271 -901 -255 -867
rect -321 -935 -255 -901
rect -321 -969 -305 -935
rect -271 -969 -255 -935
rect -321 -1000 -255 -969
rect -225 969 -159 1000
rect -225 935 -209 969
rect -175 935 -159 969
rect -225 901 -159 935
rect -225 867 -209 901
rect -175 867 -159 901
rect -225 833 -159 867
rect -225 799 -209 833
rect -175 799 -159 833
rect -225 765 -159 799
rect -225 731 -209 765
rect -175 731 -159 765
rect -225 697 -159 731
rect -225 663 -209 697
rect -175 663 -159 697
rect -225 629 -159 663
rect -225 595 -209 629
rect -175 595 -159 629
rect -225 561 -159 595
rect -225 527 -209 561
rect -175 527 -159 561
rect -225 493 -159 527
rect -225 459 -209 493
rect -175 459 -159 493
rect -225 425 -159 459
rect -225 391 -209 425
rect -175 391 -159 425
rect -225 357 -159 391
rect -225 323 -209 357
rect -175 323 -159 357
rect -225 289 -159 323
rect -225 255 -209 289
rect -175 255 -159 289
rect -225 221 -159 255
rect -225 187 -209 221
rect -175 187 -159 221
rect -225 153 -159 187
rect -225 119 -209 153
rect -175 119 -159 153
rect -225 85 -159 119
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -119 -159 -85
rect -225 -153 -209 -119
rect -175 -153 -159 -119
rect -225 -187 -159 -153
rect -225 -221 -209 -187
rect -175 -221 -159 -187
rect -225 -255 -159 -221
rect -225 -289 -209 -255
rect -175 -289 -159 -255
rect -225 -323 -159 -289
rect -225 -357 -209 -323
rect -175 -357 -159 -323
rect -225 -391 -159 -357
rect -225 -425 -209 -391
rect -175 -425 -159 -391
rect -225 -459 -159 -425
rect -225 -493 -209 -459
rect -175 -493 -159 -459
rect -225 -527 -159 -493
rect -225 -561 -209 -527
rect -175 -561 -159 -527
rect -225 -595 -159 -561
rect -225 -629 -209 -595
rect -175 -629 -159 -595
rect -225 -663 -159 -629
rect -225 -697 -209 -663
rect -175 -697 -159 -663
rect -225 -731 -159 -697
rect -225 -765 -209 -731
rect -175 -765 -159 -731
rect -225 -799 -159 -765
rect -225 -833 -209 -799
rect -175 -833 -159 -799
rect -225 -867 -159 -833
rect -225 -901 -209 -867
rect -175 -901 -159 -867
rect -225 -935 -159 -901
rect -225 -969 -209 -935
rect -175 -969 -159 -935
rect -225 -1000 -159 -969
rect -129 969 -63 1000
rect -129 935 -113 969
rect -79 935 -63 969
rect -129 901 -63 935
rect -129 867 -113 901
rect -79 867 -63 901
rect -129 833 -63 867
rect -129 799 -113 833
rect -79 799 -63 833
rect -129 765 -63 799
rect -129 731 -113 765
rect -79 731 -63 765
rect -129 697 -63 731
rect -129 663 -113 697
rect -79 663 -63 697
rect -129 629 -63 663
rect -129 595 -113 629
rect -79 595 -63 629
rect -129 561 -63 595
rect -129 527 -113 561
rect -79 527 -63 561
rect -129 493 -63 527
rect -129 459 -113 493
rect -79 459 -63 493
rect -129 425 -63 459
rect -129 391 -113 425
rect -79 391 -63 425
rect -129 357 -63 391
rect -129 323 -113 357
rect -79 323 -63 357
rect -129 289 -63 323
rect -129 255 -113 289
rect -79 255 -63 289
rect -129 221 -63 255
rect -129 187 -113 221
rect -79 187 -63 221
rect -129 153 -63 187
rect -129 119 -113 153
rect -79 119 -63 153
rect -129 85 -63 119
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -119 -63 -85
rect -129 -153 -113 -119
rect -79 -153 -63 -119
rect -129 -187 -63 -153
rect -129 -221 -113 -187
rect -79 -221 -63 -187
rect -129 -255 -63 -221
rect -129 -289 -113 -255
rect -79 -289 -63 -255
rect -129 -323 -63 -289
rect -129 -357 -113 -323
rect -79 -357 -63 -323
rect -129 -391 -63 -357
rect -129 -425 -113 -391
rect -79 -425 -63 -391
rect -129 -459 -63 -425
rect -129 -493 -113 -459
rect -79 -493 -63 -459
rect -129 -527 -63 -493
rect -129 -561 -113 -527
rect -79 -561 -63 -527
rect -129 -595 -63 -561
rect -129 -629 -113 -595
rect -79 -629 -63 -595
rect -129 -663 -63 -629
rect -129 -697 -113 -663
rect -79 -697 -63 -663
rect -129 -731 -63 -697
rect -129 -765 -113 -731
rect -79 -765 -63 -731
rect -129 -799 -63 -765
rect -129 -833 -113 -799
rect -79 -833 -63 -799
rect -129 -867 -63 -833
rect -129 -901 -113 -867
rect -79 -901 -63 -867
rect -129 -935 -63 -901
rect -129 -969 -113 -935
rect -79 -969 -63 -935
rect -129 -1000 -63 -969
rect -33 969 33 1000
rect -33 935 -17 969
rect 17 935 33 969
rect -33 901 33 935
rect -33 867 -17 901
rect 17 867 33 901
rect -33 833 33 867
rect -33 799 -17 833
rect 17 799 33 833
rect -33 765 33 799
rect -33 731 -17 765
rect 17 731 33 765
rect -33 697 33 731
rect -33 663 -17 697
rect 17 663 33 697
rect -33 629 33 663
rect -33 595 -17 629
rect 17 595 33 629
rect -33 561 33 595
rect -33 527 -17 561
rect 17 527 33 561
rect -33 493 33 527
rect -33 459 -17 493
rect 17 459 33 493
rect -33 425 33 459
rect -33 391 -17 425
rect 17 391 33 425
rect -33 357 33 391
rect -33 323 -17 357
rect 17 323 33 357
rect -33 289 33 323
rect -33 255 -17 289
rect 17 255 33 289
rect -33 221 33 255
rect -33 187 -17 221
rect 17 187 33 221
rect -33 153 33 187
rect -33 119 -17 153
rect 17 119 33 153
rect -33 85 33 119
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -119 33 -85
rect -33 -153 -17 -119
rect 17 -153 33 -119
rect -33 -187 33 -153
rect -33 -221 -17 -187
rect 17 -221 33 -187
rect -33 -255 33 -221
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -33 -323 33 -289
rect -33 -357 -17 -323
rect 17 -357 33 -323
rect -33 -391 33 -357
rect -33 -425 -17 -391
rect 17 -425 33 -391
rect -33 -459 33 -425
rect -33 -493 -17 -459
rect 17 -493 33 -459
rect -33 -527 33 -493
rect -33 -561 -17 -527
rect 17 -561 33 -527
rect -33 -595 33 -561
rect -33 -629 -17 -595
rect 17 -629 33 -595
rect -33 -663 33 -629
rect -33 -697 -17 -663
rect 17 -697 33 -663
rect -33 -731 33 -697
rect -33 -765 -17 -731
rect 17 -765 33 -731
rect -33 -799 33 -765
rect -33 -833 -17 -799
rect 17 -833 33 -799
rect -33 -867 33 -833
rect -33 -901 -17 -867
rect 17 -901 33 -867
rect -33 -935 33 -901
rect -33 -969 -17 -935
rect 17 -969 33 -935
rect -33 -1000 33 -969
rect 63 969 129 1000
rect 63 935 79 969
rect 113 935 129 969
rect 63 901 129 935
rect 63 867 79 901
rect 113 867 129 901
rect 63 833 129 867
rect 63 799 79 833
rect 113 799 129 833
rect 63 765 129 799
rect 63 731 79 765
rect 113 731 129 765
rect 63 697 129 731
rect 63 663 79 697
rect 113 663 129 697
rect 63 629 129 663
rect 63 595 79 629
rect 113 595 129 629
rect 63 561 129 595
rect 63 527 79 561
rect 113 527 129 561
rect 63 493 129 527
rect 63 459 79 493
rect 113 459 129 493
rect 63 425 129 459
rect 63 391 79 425
rect 113 391 129 425
rect 63 357 129 391
rect 63 323 79 357
rect 113 323 129 357
rect 63 289 129 323
rect 63 255 79 289
rect 113 255 129 289
rect 63 221 129 255
rect 63 187 79 221
rect 113 187 129 221
rect 63 153 129 187
rect 63 119 79 153
rect 113 119 129 153
rect 63 85 129 119
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -119 129 -85
rect 63 -153 79 -119
rect 113 -153 129 -119
rect 63 -187 129 -153
rect 63 -221 79 -187
rect 113 -221 129 -187
rect 63 -255 129 -221
rect 63 -289 79 -255
rect 113 -289 129 -255
rect 63 -323 129 -289
rect 63 -357 79 -323
rect 113 -357 129 -323
rect 63 -391 129 -357
rect 63 -425 79 -391
rect 113 -425 129 -391
rect 63 -459 129 -425
rect 63 -493 79 -459
rect 113 -493 129 -459
rect 63 -527 129 -493
rect 63 -561 79 -527
rect 113 -561 129 -527
rect 63 -595 129 -561
rect 63 -629 79 -595
rect 113 -629 129 -595
rect 63 -663 129 -629
rect 63 -697 79 -663
rect 113 -697 129 -663
rect 63 -731 129 -697
rect 63 -765 79 -731
rect 113 -765 129 -731
rect 63 -799 129 -765
rect 63 -833 79 -799
rect 113 -833 129 -799
rect 63 -867 129 -833
rect 63 -901 79 -867
rect 113 -901 129 -867
rect 63 -935 129 -901
rect 63 -969 79 -935
rect 113 -969 129 -935
rect 63 -1000 129 -969
rect 159 969 225 1000
rect 159 935 175 969
rect 209 935 225 969
rect 159 901 225 935
rect 159 867 175 901
rect 209 867 225 901
rect 159 833 225 867
rect 159 799 175 833
rect 209 799 225 833
rect 159 765 225 799
rect 159 731 175 765
rect 209 731 225 765
rect 159 697 225 731
rect 159 663 175 697
rect 209 663 225 697
rect 159 629 225 663
rect 159 595 175 629
rect 209 595 225 629
rect 159 561 225 595
rect 159 527 175 561
rect 209 527 225 561
rect 159 493 225 527
rect 159 459 175 493
rect 209 459 225 493
rect 159 425 225 459
rect 159 391 175 425
rect 209 391 225 425
rect 159 357 225 391
rect 159 323 175 357
rect 209 323 225 357
rect 159 289 225 323
rect 159 255 175 289
rect 209 255 225 289
rect 159 221 225 255
rect 159 187 175 221
rect 209 187 225 221
rect 159 153 225 187
rect 159 119 175 153
rect 209 119 225 153
rect 159 85 225 119
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -119 225 -85
rect 159 -153 175 -119
rect 209 -153 225 -119
rect 159 -187 225 -153
rect 159 -221 175 -187
rect 209 -221 225 -187
rect 159 -255 225 -221
rect 159 -289 175 -255
rect 209 -289 225 -255
rect 159 -323 225 -289
rect 159 -357 175 -323
rect 209 -357 225 -323
rect 159 -391 225 -357
rect 159 -425 175 -391
rect 209 -425 225 -391
rect 159 -459 225 -425
rect 159 -493 175 -459
rect 209 -493 225 -459
rect 159 -527 225 -493
rect 159 -561 175 -527
rect 209 -561 225 -527
rect 159 -595 225 -561
rect 159 -629 175 -595
rect 209 -629 225 -595
rect 159 -663 225 -629
rect 159 -697 175 -663
rect 209 -697 225 -663
rect 159 -731 225 -697
rect 159 -765 175 -731
rect 209 -765 225 -731
rect 159 -799 225 -765
rect 159 -833 175 -799
rect 209 -833 225 -799
rect 159 -867 225 -833
rect 159 -901 175 -867
rect 209 -901 225 -867
rect 159 -935 225 -901
rect 159 -969 175 -935
rect 209 -969 225 -935
rect 159 -1000 225 -969
rect 255 969 321 1000
rect 255 935 271 969
rect 305 935 321 969
rect 255 901 321 935
rect 255 867 271 901
rect 305 867 321 901
rect 255 833 321 867
rect 255 799 271 833
rect 305 799 321 833
rect 255 765 321 799
rect 255 731 271 765
rect 305 731 321 765
rect 255 697 321 731
rect 255 663 271 697
rect 305 663 321 697
rect 255 629 321 663
rect 255 595 271 629
rect 305 595 321 629
rect 255 561 321 595
rect 255 527 271 561
rect 305 527 321 561
rect 255 493 321 527
rect 255 459 271 493
rect 305 459 321 493
rect 255 425 321 459
rect 255 391 271 425
rect 305 391 321 425
rect 255 357 321 391
rect 255 323 271 357
rect 305 323 321 357
rect 255 289 321 323
rect 255 255 271 289
rect 305 255 321 289
rect 255 221 321 255
rect 255 187 271 221
rect 305 187 321 221
rect 255 153 321 187
rect 255 119 271 153
rect 305 119 321 153
rect 255 85 321 119
rect 255 51 271 85
rect 305 51 321 85
rect 255 17 321 51
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -51 321 -17
rect 255 -85 271 -51
rect 305 -85 321 -51
rect 255 -119 321 -85
rect 255 -153 271 -119
rect 305 -153 321 -119
rect 255 -187 321 -153
rect 255 -221 271 -187
rect 305 -221 321 -187
rect 255 -255 321 -221
rect 255 -289 271 -255
rect 305 -289 321 -255
rect 255 -323 321 -289
rect 255 -357 271 -323
rect 305 -357 321 -323
rect 255 -391 321 -357
rect 255 -425 271 -391
rect 305 -425 321 -391
rect 255 -459 321 -425
rect 255 -493 271 -459
rect 305 -493 321 -459
rect 255 -527 321 -493
rect 255 -561 271 -527
rect 305 -561 321 -527
rect 255 -595 321 -561
rect 255 -629 271 -595
rect 305 -629 321 -595
rect 255 -663 321 -629
rect 255 -697 271 -663
rect 305 -697 321 -663
rect 255 -731 321 -697
rect 255 -765 271 -731
rect 305 -765 321 -731
rect 255 -799 321 -765
rect 255 -833 271 -799
rect 305 -833 321 -799
rect 255 -867 321 -833
rect 255 -901 271 -867
rect 305 -901 321 -867
rect 255 -935 321 -901
rect 255 -969 271 -935
rect 305 -969 321 -935
rect 255 -1000 321 -969
rect 351 969 417 1000
rect 351 935 367 969
rect 401 935 417 969
rect 351 901 417 935
rect 351 867 367 901
rect 401 867 417 901
rect 351 833 417 867
rect 351 799 367 833
rect 401 799 417 833
rect 351 765 417 799
rect 351 731 367 765
rect 401 731 417 765
rect 351 697 417 731
rect 351 663 367 697
rect 401 663 417 697
rect 351 629 417 663
rect 351 595 367 629
rect 401 595 417 629
rect 351 561 417 595
rect 351 527 367 561
rect 401 527 417 561
rect 351 493 417 527
rect 351 459 367 493
rect 401 459 417 493
rect 351 425 417 459
rect 351 391 367 425
rect 401 391 417 425
rect 351 357 417 391
rect 351 323 367 357
rect 401 323 417 357
rect 351 289 417 323
rect 351 255 367 289
rect 401 255 417 289
rect 351 221 417 255
rect 351 187 367 221
rect 401 187 417 221
rect 351 153 417 187
rect 351 119 367 153
rect 401 119 417 153
rect 351 85 417 119
rect 351 51 367 85
rect 401 51 417 85
rect 351 17 417 51
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -51 417 -17
rect 351 -85 367 -51
rect 401 -85 417 -51
rect 351 -119 417 -85
rect 351 -153 367 -119
rect 401 -153 417 -119
rect 351 -187 417 -153
rect 351 -221 367 -187
rect 401 -221 417 -187
rect 351 -255 417 -221
rect 351 -289 367 -255
rect 401 -289 417 -255
rect 351 -323 417 -289
rect 351 -357 367 -323
rect 401 -357 417 -323
rect 351 -391 417 -357
rect 351 -425 367 -391
rect 401 -425 417 -391
rect 351 -459 417 -425
rect 351 -493 367 -459
rect 401 -493 417 -459
rect 351 -527 417 -493
rect 351 -561 367 -527
rect 401 -561 417 -527
rect 351 -595 417 -561
rect 351 -629 367 -595
rect 401 -629 417 -595
rect 351 -663 417 -629
rect 351 -697 367 -663
rect 401 -697 417 -663
rect 351 -731 417 -697
rect 351 -765 367 -731
rect 401 -765 417 -731
rect 351 -799 417 -765
rect 351 -833 367 -799
rect 401 -833 417 -799
rect 351 -867 417 -833
rect 351 -901 367 -867
rect 401 -901 417 -867
rect 351 -935 417 -901
rect 351 -969 367 -935
rect 401 -969 417 -935
rect 351 -1000 417 -969
rect 447 969 513 1000
rect 447 935 463 969
rect 497 935 513 969
rect 447 901 513 935
rect 447 867 463 901
rect 497 867 513 901
rect 447 833 513 867
rect 447 799 463 833
rect 497 799 513 833
rect 447 765 513 799
rect 447 731 463 765
rect 497 731 513 765
rect 447 697 513 731
rect 447 663 463 697
rect 497 663 513 697
rect 447 629 513 663
rect 447 595 463 629
rect 497 595 513 629
rect 447 561 513 595
rect 447 527 463 561
rect 497 527 513 561
rect 447 493 513 527
rect 447 459 463 493
rect 497 459 513 493
rect 447 425 513 459
rect 447 391 463 425
rect 497 391 513 425
rect 447 357 513 391
rect 447 323 463 357
rect 497 323 513 357
rect 447 289 513 323
rect 447 255 463 289
rect 497 255 513 289
rect 447 221 513 255
rect 447 187 463 221
rect 497 187 513 221
rect 447 153 513 187
rect 447 119 463 153
rect 497 119 513 153
rect 447 85 513 119
rect 447 51 463 85
rect 497 51 513 85
rect 447 17 513 51
rect 447 -17 463 17
rect 497 -17 513 17
rect 447 -51 513 -17
rect 447 -85 463 -51
rect 497 -85 513 -51
rect 447 -119 513 -85
rect 447 -153 463 -119
rect 497 -153 513 -119
rect 447 -187 513 -153
rect 447 -221 463 -187
rect 497 -221 513 -187
rect 447 -255 513 -221
rect 447 -289 463 -255
rect 497 -289 513 -255
rect 447 -323 513 -289
rect 447 -357 463 -323
rect 497 -357 513 -323
rect 447 -391 513 -357
rect 447 -425 463 -391
rect 497 -425 513 -391
rect 447 -459 513 -425
rect 447 -493 463 -459
rect 497 -493 513 -459
rect 447 -527 513 -493
rect 447 -561 463 -527
rect 497 -561 513 -527
rect 447 -595 513 -561
rect 447 -629 463 -595
rect 497 -629 513 -595
rect 447 -663 513 -629
rect 447 -697 463 -663
rect 497 -697 513 -663
rect 447 -731 513 -697
rect 447 -765 463 -731
rect 497 -765 513 -731
rect 447 -799 513 -765
rect 447 -833 463 -799
rect 497 -833 513 -799
rect 447 -867 513 -833
rect 447 -901 463 -867
rect 497 -901 513 -867
rect 447 -935 513 -901
rect 447 -969 463 -935
rect 497 -969 513 -935
rect 447 -1000 513 -969
rect 543 969 609 1000
rect 543 935 559 969
rect 593 935 609 969
rect 543 901 609 935
rect 543 867 559 901
rect 593 867 609 901
rect 543 833 609 867
rect 543 799 559 833
rect 593 799 609 833
rect 543 765 609 799
rect 543 731 559 765
rect 593 731 609 765
rect 543 697 609 731
rect 543 663 559 697
rect 593 663 609 697
rect 543 629 609 663
rect 543 595 559 629
rect 593 595 609 629
rect 543 561 609 595
rect 543 527 559 561
rect 593 527 609 561
rect 543 493 609 527
rect 543 459 559 493
rect 593 459 609 493
rect 543 425 609 459
rect 543 391 559 425
rect 593 391 609 425
rect 543 357 609 391
rect 543 323 559 357
rect 593 323 609 357
rect 543 289 609 323
rect 543 255 559 289
rect 593 255 609 289
rect 543 221 609 255
rect 543 187 559 221
rect 593 187 609 221
rect 543 153 609 187
rect 543 119 559 153
rect 593 119 609 153
rect 543 85 609 119
rect 543 51 559 85
rect 593 51 609 85
rect 543 17 609 51
rect 543 -17 559 17
rect 593 -17 609 17
rect 543 -51 609 -17
rect 543 -85 559 -51
rect 593 -85 609 -51
rect 543 -119 609 -85
rect 543 -153 559 -119
rect 593 -153 609 -119
rect 543 -187 609 -153
rect 543 -221 559 -187
rect 593 -221 609 -187
rect 543 -255 609 -221
rect 543 -289 559 -255
rect 593 -289 609 -255
rect 543 -323 609 -289
rect 543 -357 559 -323
rect 593 -357 609 -323
rect 543 -391 609 -357
rect 543 -425 559 -391
rect 593 -425 609 -391
rect 543 -459 609 -425
rect 543 -493 559 -459
rect 593 -493 609 -459
rect 543 -527 609 -493
rect 543 -561 559 -527
rect 593 -561 609 -527
rect 543 -595 609 -561
rect 543 -629 559 -595
rect 593 -629 609 -595
rect 543 -663 609 -629
rect 543 -697 559 -663
rect 593 -697 609 -663
rect 543 -731 609 -697
rect 543 -765 559 -731
rect 593 -765 609 -731
rect 543 -799 609 -765
rect 543 -833 559 -799
rect 593 -833 609 -799
rect 543 -867 609 -833
rect 543 -901 559 -867
rect 593 -901 609 -867
rect 543 -935 609 -901
rect 543 -969 559 -935
rect 593 -969 609 -935
rect 543 -1000 609 -969
rect 639 969 705 1000
rect 639 935 655 969
rect 689 935 705 969
rect 639 901 705 935
rect 639 867 655 901
rect 689 867 705 901
rect 639 833 705 867
rect 639 799 655 833
rect 689 799 705 833
rect 639 765 705 799
rect 639 731 655 765
rect 689 731 705 765
rect 639 697 705 731
rect 639 663 655 697
rect 689 663 705 697
rect 639 629 705 663
rect 639 595 655 629
rect 689 595 705 629
rect 639 561 705 595
rect 639 527 655 561
rect 689 527 705 561
rect 639 493 705 527
rect 639 459 655 493
rect 689 459 705 493
rect 639 425 705 459
rect 639 391 655 425
rect 689 391 705 425
rect 639 357 705 391
rect 639 323 655 357
rect 689 323 705 357
rect 639 289 705 323
rect 639 255 655 289
rect 689 255 705 289
rect 639 221 705 255
rect 639 187 655 221
rect 689 187 705 221
rect 639 153 705 187
rect 639 119 655 153
rect 689 119 705 153
rect 639 85 705 119
rect 639 51 655 85
rect 689 51 705 85
rect 639 17 705 51
rect 639 -17 655 17
rect 689 -17 705 17
rect 639 -51 705 -17
rect 639 -85 655 -51
rect 689 -85 705 -51
rect 639 -119 705 -85
rect 639 -153 655 -119
rect 689 -153 705 -119
rect 639 -187 705 -153
rect 639 -221 655 -187
rect 689 -221 705 -187
rect 639 -255 705 -221
rect 639 -289 655 -255
rect 689 -289 705 -255
rect 639 -323 705 -289
rect 639 -357 655 -323
rect 689 -357 705 -323
rect 639 -391 705 -357
rect 639 -425 655 -391
rect 689 -425 705 -391
rect 639 -459 705 -425
rect 639 -493 655 -459
rect 689 -493 705 -459
rect 639 -527 705 -493
rect 639 -561 655 -527
rect 689 -561 705 -527
rect 639 -595 705 -561
rect 639 -629 655 -595
rect 689 -629 705 -595
rect 639 -663 705 -629
rect 639 -697 655 -663
rect 689 -697 705 -663
rect 639 -731 705 -697
rect 639 -765 655 -731
rect 689 -765 705 -731
rect 639 -799 705 -765
rect 639 -833 655 -799
rect 689 -833 705 -799
rect 639 -867 705 -833
rect 639 -901 655 -867
rect 689 -901 705 -867
rect 639 -935 705 -901
rect 639 -969 655 -935
rect 689 -969 705 -935
rect 639 -1000 705 -969
rect 735 969 801 1000
rect 735 935 751 969
rect 785 935 801 969
rect 735 901 801 935
rect 735 867 751 901
rect 785 867 801 901
rect 735 833 801 867
rect 735 799 751 833
rect 785 799 801 833
rect 735 765 801 799
rect 735 731 751 765
rect 785 731 801 765
rect 735 697 801 731
rect 735 663 751 697
rect 785 663 801 697
rect 735 629 801 663
rect 735 595 751 629
rect 785 595 801 629
rect 735 561 801 595
rect 735 527 751 561
rect 785 527 801 561
rect 735 493 801 527
rect 735 459 751 493
rect 785 459 801 493
rect 735 425 801 459
rect 735 391 751 425
rect 785 391 801 425
rect 735 357 801 391
rect 735 323 751 357
rect 785 323 801 357
rect 735 289 801 323
rect 735 255 751 289
rect 785 255 801 289
rect 735 221 801 255
rect 735 187 751 221
rect 785 187 801 221
rect 735 153 801 187
rect 735 119 751 153
rect 785 119 801 153
rect 735 85 801 119
rect 735 51 751 85
rect 785 51 801 85
rect 735 17 801 51
rect 735 -17 751 17
rect 785 -17 801 17
rect 735 -51 801 -17
rect 735 -85 751 -51
rect 785 -85 801 -51
rect 735 -119 801 -85
rect 735 -153 751 -119
rect 785 -153 801 -119
rect 735 -187 801 -153
rect 735 -221 751 -187
rect 785 -221 801 -187
rect 735 -255 801 -221
rect 735 -289 751 -255
rect 785 -289 801 -255
rect 735 -323 801 -289
rect 735 -357 751 -323
rect 785 -357 801 -323
rect 735 -391 801 -357
rect 735 -425 751 -391
rect 785 -425 801 -391
rect 735 -459 801 -425
rect 735 -493 751 -459
rect 785 -493 801 -459
rect 735 -527 801 -493
rect 735 -561 751 -527
rect 785 -561 801 -527
rect 735 -595 801 -561
rect 735 -629 751 -595
rect 785 -629 801 -595
rect 735 -663 801 -629
rect 735 -697 751 -663
rect 785 -697 801 -663
rect 735 -731 801 -697
rect 735 -765 751 -731
rect 785 -765 801 -731
rect 735 -799 801 -765
rect 735 -833 751 -799
rect 785 -833 801 -799
rect 735 -867 801 -833
rect 735 -901 751 -867
rect 785 -901 801 -867
rect 735 -935 801 -901
rect 735 -969 751 -935
rect 785 -969 801 -935
rect 735 -1000 801 -969
rect 831 969 897 1000
rect 831 935 847 969
rect 881 935 897 969
rect 831 901 897 935
rect 831 867 847 901
rect 881 867 897 901
rect 831 833 897 867
rect 831 799 847 833
rect 881 799 897 833
rect 831 765 897 799
rect 831 731 847 765
rect 881 731 897 765
rect 831 697 897 731
rect 831 663 847 697
rect 881 663 897 697
rect 831 629 897 663
rect 831 595 847 629
rect 881 595 897 629
rect 831 561 897 595
rect 831 527 847 561
rect 881 527 897 561
rect 831 493 897 527
rect 831 459 847 493
rect 881 459 897 493
rect 831 425 897 459
rect 831 391 847 425
rect 881 391 897 425
rect 831 357 897 391
rect 831 323 847 357
rect 881 323 897 357
rect 831 289 897 323
rect 831 255 847 289
rect 881 255 897 289
rect 831 221 897 255
rect 831 187 847 221
rect 881 187 897 221
rect 831 153 897 187
rect 831 119 847 153
rect 881 119 897 153
rect 831 85 897 119
rect 831 51 847 85
rect 881 51 897 85
rect 831 17 897 51
rect 831 -17 847 17
rect 881 -17 897 17
rect 831 -51 897 -17
rect 831 -85 847 -51
rect 881 -85 897 -51
rect 831 -119 897 -85
rect 831 -153 847 -119
rect 881 -153 897 -119
rect 831 -187 897 -153
rect 831 -221 847 -187
rect 881 -221 897 -187
rect 831 -255 897 -221
rect 831 -289 847 -255
rect 881 -289 897 -255
rect 831 -323 897 -289
rect 831 -357 847 -323
rect 881 -357 897 -323
rect 831 -391 897 -357
rect 831 -425 847 -391
rect 881 -425 897 -391
rect 831 -459 897 -425
rect 831 -493 847 -459
rect 881 -493 897 -459
rect 831 -527 897 -493
rect 831 -561 847 -527
rect 881 -561 897 -527
rect 831 -595 897 -561
rect 831 -629 847 -595
rect 881 -629 897 -595
rect 831 -663 897 -629
rect 831 -697 847 -663
rect 881 -697 897 -663
rect 831 -731 897 -697
rect 831 -765 847 -731
rect 881 -765 897 -731
rect 831 -799 897 -765
rect 831 -833 847 -799
rect 881 -833 897 -799
rect 831 -867 897 -833
rect 831 -901 847 -867
rect 881 -901 897 -867
rect 831 -935 897 -901
rect 831 -969 847 -935
rect 881 -969 897 -935
rect 831 -1000 897 -969
rect 927 969 993 1000
rect 927 935 943 969
rect 977 935 993 969
rect 927 901 993 935
rect 927 867 943 901
rect 977 867 993 901
rect 927 833 993 867
rect 927 799 943 833
rect 977 799 993 833
rect 927 765 993 799
rect 927 731 943 765
rect 977 731 993 765
rect 927 697 993 731
rect 927 663 943 697
rect 977 663 993 697
rect 927 629 993 663
rect 927 595 943 629
rect 977 595 993 629
rect 927 561 993 595
rect 927 527 943 561
rect 977 527 993 561
rect 927 493 993 527
rect 927 459 943 493
rect 977 459 993 493
rect 927 425 993 459
rect 927 391 943 425
rect 977 391 993 425
rect 927 357 993 391
rect 927 323 943 357
rect 977 323 993 357
rect 927 289 993 323
rect 927 255 943 289
rect 977 255 993 289
rect 927 221 993 255
rect 927 187 943 221
rect 977 187 993 221
rect 927 153 993 187
rect 927 119 943 153
rect 977 119 993 153
rect 927 85 993 119
rect 927 51 943 85
rect 977 51 993 85
rect 927 17 993 51
rect 927 -17 943 17
rect 977 -17 993 17
rect 927 -51 993 -17
rect 927 -85 943 -51
rect 977 -85 993 -51
rect 927 -119 993 -85
rect 927 -153 943 -119
rect 977 -153 993 -119
rect 927 -187 993 -153
rect 927 -221 943 -187
rect 977 -221 993 -187
rect 927 -255 993 -221
rect 927 -289 943 -255
rect 977 -289 993 -255
rect 927 -323 993 -289
rect 927 -357 943 -323
rect 977 -357 993 -323
rect 927 -391 993 -357
rect 927 -425 943 -391
rect 977 -425 993 -391
rect 927 -459 993 -425
rect 927 -493 943 -459
rect 977 -493 993 -459
rect 927 -527 993 -493
rect 927 -561 943 -527
rect 977 -561 993 -527
rect 927 -595 993 -561
rect 927 -629 943 -595
rect 977 -629 993 -595
rect 927 -663 993 -629
rect 927 -697 943 -663
rect 977 -697 993 -663
rect 927 -731 993 -697
rect 927 -765 943 -731
rect 977 -765 993 -731
rect 927 -799 993 -765
rect 927 -833 943 -799
rect 977 -833 993 -799
rect 927 -867 993 -833
rect 927 -901 943 -867
rect 977 -901 993 -867
rect 927 -935 993 -901
rect 927 -969 943 -935
rect 977 -969 993 -935
rect 927 -1000 993 -969
rect 1023 969 1089 1000
rect 1023 935 1039 969
rect 1073 935 1089 969
rect 1023 901 1089 935
rect 1023 867 1039 901
rect 1073 867 1089 901
rect 1023 833 1089 867
rect 1023 799 1039 833
rect 1073 799 1089 833
rect 1023 765 1089 799
rect 1023 731 1039 765
rect 1073 731 1089 765
rect 1023 697 1089 731
rect 1023 663 1039 697
rect 1073 663 1089 697
rect 1023 629 1089 663
rect 1023 595 1039 629
rect 1073 595 1089 629
rect 1023 561 1089 595
rect 1023 527 1039 561
rect 1073 527 1089 561
rect 1023 493 1089 527
rect 1023 459 1039 493
rect 1073 459 1089 493
rect 1023 425 1089 459
rect 1023 391 1039 425
rect 1073 391 1089 425
rect 1023 357 1089 391
rect 1023 323 1039 357
rect 1073 323 1089 357
rect 1023 289 1089 323
rect 1023 255 1039 289
rect 1073 255 1089 289
rect 1023 221 1089 255
rect 1023 187 1039 221
rect 1073 187 1089 221
rect 1023 153 1089 187
rect 1023 119 1039 153
rect 1073 119 1089 153
rect 1023 85 1089 119
rect 1023 51 1039 85
rect 1073 51 1089 85
rect 1023 17 1089 51
rect 1023 -17 1039 17
rect 1073 -17 1089 17
rect 1023 -51 1089 -17
rect 1023 -85 1039 -51
rect 1073 -85 1089 -51
rect 1023 -119 1089 -85
rect 1023 -153 1039 -119
rect 1073 -153 1089 -119
rect 1023 -187 1089 -153
rect 1023 -221 1039 -187
rect 1073 -221 1089 -187
rect 1023 -255 1089 -221
rect 1023 -289 1039 -255
rect 1073 -289 1089 -255
rect 1023 -323 1089 -289
rect 1023 -357 1039 -323
rect 1073 -357 1089 -323
rect 1023 -391 1089 -357
rect 1023 -425 1039 -391
rect 1073 -425 1089 -391
rect 1023 -459 1089 -425
rect 1023 -493 1039 -459
rect 1073 -493 1089 -459
rect 1023 -527 1089 -493
rect 1023 -561 1039 -527
rect 1073 -561 1089 -527
rect 1023 -595 1089 -561
rect 1023 -629 1039 -595
rect 1073 -629 1089 -595
rect 1023 -663 1089 -629
rect 1023 -697 1039 -663
rect 1073 -697 1089 -663
rect 1023 -731 1089 -697
rect 1023 -765 1039 -731
rect 1073 -765 1089 -731
rect 1023 -799 1089 -765
rect 1023 -833 1039 -799
rect 1073 -833 1089 -799
rect 1023 -867 1089 -833
rect 1023 -901 1039 -867
rect 1073 -901 1089 -867
rect 1023 -935 1089 -901
rect 1023 -969 1039 -935
rect 1073 -969 1089 -935
rect 1023 -1000 1089 -969
rect 1119 969 1185 1000
rect 1119 935 1135 969
rect 1169 935 1185 969
rect 1119 901 1185 935
rect 1119 867 1135 901
rect 1169 867 1185 901
rect 1119 833 1185 867
rect 1119 799 1135 833
rect 1169 799 1185 833
rect 1119 765 1185 799
rect 1119 731 1135 765
rect 1169 731 1185 765
rect 1119 697 1185 731
rect 1119 663 1135 697
rect 1169 663 1185 697
rect 1119 629 1185 663
rect 1119 595 1135 629
rect 1169 595 1185 629
rect 1119 561 1185 595
rect 1119 527 1135 561
rect 1169 527 1185 561
rect 1119 493 1185 527
rect 1119 459 1135 493
rect 1169 459 1185 493
rect 1119 425 1185 459
rect 1119 391 1135 425
rect 1169 391 1185 425
rect 1119 357 1185 391
rect 1119 323 1135 357
rect 1169 323 1185 357
rect 1119 289 1185 323
rect 1119 255 1135 289
rect 1169 255 1185 289
rect 1119 221 1185 255
rect 1119 187 1135 221
rect 1169 187 1185 221
rect 1119 153 1185 187
rect 1119 119 1135 153
rect 1169 119 1185 153
rect 1119 85 1185 119
rect 1119 51 1135 85
rect 1169 51 1185 85
rect 1119 17 1185 51
rect 1119 -17 1135 17
rect 1169 -17 1185 17
rect 1119 -51 1185 -17
rect 1119 -85 1135 -51
rect 1169 -85 1185 -51
rect 1119 -119 1185 -85
rect 1119 -153 1135 -119
rect 1169 -153 1185 -119
rect 1119 -187 1185 -153
rect 1119 -221 1135 -187
rect 1169 -221 1185 -187
rect 1119 -255 1185 -221
rect 1119 -289 1135 -255
rect 1169 -289 1185 -255
rect 1119 -323 1185 -289
rect 1119 -357 1135 -323
rect 1169 -357 1185 -323
rect 1119 -391 1185 -357
rect 1119 -425 1135 -391
rect 1169 -425 1185 -391
rect 1119 -459 1185 -425
rect 1119 -493 1135 -459
rect 1169 -493 1185 -459
rect 1119 -527 1185 -493
rect 1119 -561 1135 -527
rect 1169 -561 1185 -527
rect 1119 -595 1185 -561
rect 1119 -629 1135 -595
rect 1169 -629 1185 -595
rect 1119 -663 1185 -629
rect 1119 -697 1135 -663
rect 1169 -697 1185 -663
rect 1119 -731 1185 -697
rect 1119 -765 1135 -731
rect 1169 -765 1185 -731
rect 1119 -799 1185 -765
rect 1119 -833 1135 -799
rect 1169 -833 1185 -799
rect 1119 -867 1185 -833
rect 1119 -901 1135 -867
rect 1169 -901 1185 -867
rect 1119 -935 1185 -901
rect 1119 -969 1135 -935
rect 1169 -969 1185 -935
rect 1119 -1000 1185 -969
rect 1215 969 1281 1000
rect 1215 935 1231 969
rect 1265 935 1281 969
rect 1215 901 1281 935
rect 1215 867 1231 901
rect 1265 867 1281 901
rect 1215 833 1281 867
rect 1215 799 1231 833
rect 1265 799 1281 833
rect 1215 765 1281 799
rect 1215 731 1231 765
rect 1265 731 1281 765
rect 1215 697 1281 731
rect 1215 663 1231 697
rect 1265 663 1281 697
rect 1215 629 1281 663
rect 1215 595 1231 629
rect 1265 595 1281 629
rect 1215 561 1281 595
rect 1215 527 1231 561
rect 1265 527 1281 561
rect 1215 493 1281 527
rect 1215 459 1231 493
rect 1265 459 1281 493
rect 1215 425 1281 459
rect 1215 391 1231 425
rect 1265 391 1281 425
rect 1215 357 1281 391
rect 1215 323 1231 357
rect 1265 323 1281 357
rect 1215 289 1281 323
rect 1215 255 1231 289
rect 1265 255 1281 289
rect 1215 221 1281 255
rect 1215 187 1231 221
rect 1265 187 1281 221
rect 1215 153 1281 187
rect 1215 119 1231 153
rect 1265 119 1281 153
rect 1215 85 1281 119
rect 1215 51 1231 85
rect 1265 51 1281 85
rect 1215 17 1281 51
rect 1215 -17 1231 17
rect 1265 -17 1281 17
rect 1215 -51 1281 -17
rect 1215 -85 1231 -51
rect 1265 -85 1281 -51
rect 1215 -119 1281 -85
rect 1215 -153 1231 -119
rect 1265 -153 1281 -119
rect 1215 -187 1281 -153
rect 1215 -221 1231 -187
rect 1265 -221 1281 -187
rect 1215 -255 1281 -221
rect 1215 -289 1231 -255
rect 1265 -289 1281 -255
rect 1215 -323 1281 -289
rect 1215 -357 1231 -323
rect 1265 -357 1281 -323
rect 1215 -391 1281 -357
rect 1215 -425 1231 -391
rect 1265 -425 1281 -391
rect 1215 -459 1281 -425
rect 1215 -493 1231 -459
rect 1265 -493 1281 -459
rect 1215 -527 1281 -493
rect 1215 -561 1231 -527
rect 1265 -561 1281 -527
rect 1215 -595 1281 -561
rect 1215 -629 1231 -595
rect 1265 -629 1281 -595
rect 1215 -663 1281 -629
rect 1215 -697 1231 -663
rect 1265 -697 1281 -663
rect 1215 -731 1281 -697
rect 1215 -765 1231 -731
rect 1265 -765 1281 -731
rect 1215 -799 1281 -765
rect 1215 -833 1231 -799
rect 1265 -833 1281 -799
rect 1215 -867 1281 -833
rect 1215 -901 1231 -867
rect 1265 -901 1281 -867
rect 1215 -935 1281 -901
rect 1215 -969 1231 -935
rect 1265 -969 1281 -935
rect 1215 -1000 1281 -969
rect 1311 969 1377 1000
rect 1311 935 1327 969
rect 1361 935 1377 969
rect 1311 901 1377 935
rect 1311 867 1327 901
rect 1361 867 1377 901
rect 1311 833 1377 867
rect 1311 799 1327 833
rect 1361 799 1377 833
rect 1311 765 1377 799
rect 1311 731 1327 765
rect 1361 731 1377 765
rect 1311 697 1377 731
rect 1311 663 1327 697
rect 1361 663 1377 697
rect 1311 629 1377 663
rect 1311 595 1327 629
rect 1361 595 1377 629
rect 1311 561 1377 595
rect 1311 527 1327 561
rect 1361 527 1377 561
rect 1311 493 1377 527
rect 1311 459 1327 493
rect 1361 459 1377 493
rect 1311 425 1377 459
rect 1311 391 1327 425
rect 1361 391 1377 425
rect 1311 357 1377 391
rect 1311 323 1327 357
rect 1361 323 1377 357
rect 1311 289 1377 323
rect 1311 255 1327 289
rect 1361 255 1377 289
rect 1311 221 1377 255
rect 1311 187 1327 221
rect 1361 187 1377 221
rect 1311 153 1377 187
rect 1311 119 1327 153
rect 1361 119 1377 153
rect 1311 85 1377 119
rect 1311 51 1327 85
rect 1361 51 1377 85
rect 1311 17 1377 51
rect 1311 -17 1327 17
rect 1361 -17 1377 17
rect 1311 -51 1377 -17
rect 1311 -85 1327 -51
rect 1361 -85 1377 -51
rect 1311 -119 1377 -85
rect 1311 -153 1327 -119
rect 1361 -153 1377 -119
rect 1311 -187 1377 -153
rect 1311 -221 1327 -187
rect 1361 -221 1377 -187
rect 1311 -255 1377 -221
rect 1311 -289 1327 -255
rect 1361 -289 1377 -255
rect 1311 -323 1377 -289
rect 1311 -357 1327 -323
rect 1361 -357 1377 -323
rect 1311 -391 1377 -357
rect 1311 -425 1327 -391
rect 1361 -425 1377 -391
rect 1311 -459 1377 -425
rect 1311 -493 1327 -459
rect 1361 -493 1377 -459
rect 1311 -527 1377 -493
rect 1311 -561 1327 -527
rect 1361 -561 1377 -527
rect 1311 -595 1377 -561
rect 1311 -629 1327 -595
rect 1361 -629 1377 -595
rect 1311 -663 1377 -629
rect 1311 -697 1327 -663
rect 1361 -697 1377 -663
rect 1311 -731 1377 -697
rect 1311 -765 1327 -731
rect 1361 -765 1377 -731
rect 1311 -799 1377 -765
rect 1311 -833 1327 -799
rect 1361 -833 1377 -799
rect 1311 -867 1377 -833
rect 1311 -901 1327 -867
rect 1361 -901 1377 -867
rect 1311 -935 1377 -901
rect 1311 -969 1327 -935
rect 1361 -969 1377 -935
rect 1311 -1000 1377 -969
rect 1407 969 1473 1000
rect 1407 935 1423 969
rect 1457 935 1473 969
rect 1407 901 1473 935
rect 1407 867 1423 901
rect 1457 867 1473 901
rect 1407 833 1473 867
rect 1407 799 1423 833
rect 1457 799 1473 833
rect 1407 765 1473 799
rect 1407 731 1423 765
rect 1457 731 1473 765
rect 1407 697 1473 731
rect 1407 663 1423 697
rect 1457 663 1473 697
rect 1407 629 1473 663
rect 1407 595 1423 629
rect 1457 595 1473 629
rect 1407 561 1473 595
rect 1407 527 1423 561
rect 1457 527 1473 561
rect 1407 493 1473 527
rect 1407 459 1423 493
rect 1457 459 1473 493
rect 1407 425 1473 459
rect 1407 391 1423 425
rect 1457 391 1473 425
rect 1407 357 1473 391
rect 1407 323 1423 357
rect 1457 323 1473 357
rect 1407 289 1473 323
rect 1407 255 1423 289
rect 1457 255 1473 289
rect 1407 221 1473 255
rect 1407 187 1423 221
rect 1457 187 1473 221
rect 1407 153 1473 187
rect 1407 119 1423 153
rect 1457 119 1473 153
rect 1407 85 1473 119
rect 1407 51 1423 85
rect 1457 51 1473 85
rect 1407 17 1473 51
rect 1407 -17 1423 17
rect 1457 -17 1473 17
rect 1407 -51 1473 -17
rect 1407 -85 1423 -51
rect 1457 -85 1473 -51
rect 1407 -119 1473 -85
rect 1407 -153 1423 -119
rect 1457 -153 1473 -119
rect 1407 -187 1473 -153
rect 1407 -221 1423 -187
rect 1457 -221 1473 -187
rect 1407 -255 1473 -221
rect 1407 -289 1423 -255
rect 1457 -289 1473 -255
rect 1407 -323 1473 -289
rect 1407 -357 1423 -323
rect 1457 -357 1473 -323
rect 1407 -391 1473 -357
rect 1407 -425 1423 -391
rect 1457 -425 1473 -391
rect 1407 -459 1473 -425
rect 1407 -493 1423 -459
rect 1457 -493 1473 -459
rect 1407 -527 1473 -493
rect 1407 -561 1423 -527
rect 1457 -561 1473 -527
rect 1407 -595 1473 -561
rect 1407 -629 1423 -595
rect 1457 -629 1473 -595
rect 1407 -663 1473 -629
rect 1407 -697 1423 -663
rect 1457 -697 1473 -663
rect 1407 -731 1473 -697
rect 1407 -765 1423 -731
rect 1457 -765 1473 -731
rect 1407 -799 1473 -765
rect 1407 -833 1423 -799
rect 1457 -833 1473 -799
rect 1407 -867 1473 -833
rect 1407 -901 1423 -867
rect 1457 -901 1473 -867
rect 1407 -935 1473 -901
rect 1407 -969 1423 -935
rect 1457 -969 1473 -935
rect 1407 -1000 1473 -969
rect 1503 969 1569 1000
rect 1503 935 1519 969
rect 1553 935 1569 969
rect 1503 901 1569 935
rect 1503 867 1519 901
rect 1553 867 1569 901
rect 1503 833 1569 867
rect 1503 799 1519 833
rect 1553 799 1569 833
rect 1503 765 1569 799
rect 1503 731 1519 765
rect 1553 731 1569 765
rect 1503 697 1569 731
rect 1503 663 1519 697
rect 1553 663 1569 697
rect 1503 629 1569 663
rect 1503 595 1519 629
rect 1553 595 1569 629
rect 1503 561 1569 595
rect 1503 527 1519 561
rect 1553 527 1569 561
rect 1503 493 1569 527
rect 1503 459 1519 493
rect 1553 459 1569 493
rect 1503 425 1569 459
rect 1503 391 1519 425
rect 1553 391 1569 425
rect 1503 357 1569 391
rect 1503 323 1519 357
rect 1553 323 1569 357
rect 1503 289 1569 323
rect 1503 255 1519 289
rect 1553 255 1569 289
rect 1503 221 1569 255
rect 1503 187 1519 221
rect 1553 187 1569 221
rect 1503 153 1569 187
rect 1503 119 1519 153
rect 1553 119 1569 153
rect 1503 85 1569 119
rect 1503 51 1519 85
rect 1553 51 1569 85
rect 1503 17 1569 51
rect 1503 -17 1519 17
rect 1553 -17 1569 17
rect 1503 -51 1569 -17
rect 1503 -85 1519 -51
rect 1553 -85 1569 -51
rect 1503 -119 1569 -85
rect 1503 -153 1519 -119
rect 1553 -153 1569 -119
rect 1503 -187 1569 -153
rect 1503 -221 1519 -187
rect 1553 -221 1569 -187
rect 1503 -255 1569 -221
rect 1503 -289 1519 -255
rect 1553 -289 1569 -255
rect 1503 -323 1569 -289
rect 1503 -357 1519 -323
rect 1553 -357 1569 -323
rect 1503 -391 1569 -357
rect 1503 -425 1519 -391
rect 1553 -425 1569 -391
rect 1503 -459 1569 -425
rect 1503 -493 1519 -459
rect 1553 -493 1569 -459
rect 1503 -527 1569 -493
rect 1503 -561 1519 -527
rect 1553 -561 1569 -527
rect 1503 -595 1569 -561
rect 1503 -629 1519 -595
rect 1553 -629 1569 -595
rect 1503 -663 1569 -629
rect 1503 -697 1519 -663
rect 1553 -697 1569 -663
rect 1503 -731 1569 -697
rect 1503 -765 1519 -731
rect 1553 -765 1569 -731
rect 1503 -799 1569 -765
rect 1503 -833 1519 -799
rect 1553 -833 1569 -799
rect 1503 -867 1569 -833
rect 1503 -901 1519 -867
rect 1553 -901 1569 -867
rect 1503 -935 1569 -901
rect 1503 -969 1519 -935
rect 1553 -969 1569 -935
rect 1503 -1000 1569 -969
rect 1599 969 1665 1000
rect 1599 935 1615 969
rect 1649 935 1665 969
rect 1599 901 1665 935
rect 1599 867 1615 901
rect 1649 867 1665 901
rect 1599 833 1665 867
rect 1599 799 1615 833
rect 1649 799 1665 833
rect 1599 765 1665 799
rect 1599 731 1615 765
rect 1649 731 1665 765
rect 1599 697 1665 731
rect 1599 663 1615 697
rect 1649 663 1665 697
rect 1599 629 1665 663
rect 1599 595 1615 629
rect 1649 595 1665 629
rect 1599 561 1665 595
rect 1599 527 1615 561
rect 1649 527 1665 561
rect 1599 493 1665 527
rect 1599 459 1615 493
rect 1649 459 1665 493
rect 1599 425 1665 459
rect 1599 391 1615 425
rect 1649 391 1665 425
rect 1599 357 1665 391
rect 1599 323 1615 357
rect 1649 323 1665 357
rect 1599 289 1665 323
rect 1599 255 1615 289
rect 1649 255 1665 289
rect 1599 221 1665 255
rect 1599 187 1615 221
rect 1649 187 1665 221
rect 1599 153 1665 187
rect 1599 119 1615 153
rect 1649 119 1665 153
rect 1599 85 1665 119
rect 1599 51 1615 85
rect 1649 51 1665 85
rect 1599 17 1665 51
rect 1599 -17 1615 17
rect 1649 -17 1665 17
rect 1599 -51 1665 -17
rect 1599 -85 1615 -51
rect 1649 -85 1665 -51
rect 1599 -119 1665 -85
rect 1599 -153 1615 -119
rect 1649 -153 1665 -119
rect 1599 -187 1665 -153
rect 1599 -221 1615 -187
rect 1649 -221 1665 -187
rect 1599 -255 1665 -221
rect 1599 -289 1615 -255
rect 1649 -289 1665 -255
rect 1599 -323 1665 -289
rect 1599 -357 1615 -323
rect 1649 -357 1665 -323
rect 1599 -391 1665 -357
rect 1599 -425 1615 -391
rect 1649 -425 1665 -391
rect 1599 -459 1665 -425
rect 1599 -493 1615 -459
rect 1649 -493 1665 -459
rect 1599 -527 1665 -493
rect 1599 -561 1615 -527
rect 1649 -561 1665 -527
rect 1599 -595 1665 -561
rect 1599 -629 1615 -595
rect 1649 -629 1665 -595
rect 1599 -663 1665 -629
rect 1599 -697 1615 -663
rect 1649 -697 1665 -663
rect 1599 -731 1665 -697
rect 1599 -765 1615 -731
rect 1649 -765 1665 -731
rect 1599 -799 1665 -765
rect 1599 -833 1615 -799
rect 1649 -833 1665 -799
rect 1599 -867 1665 -833
rect 1599 -901 1615 -867
rect 1649 -901 1665 -867
rect 1599 -935 1665 -901
rect 1599 -969 1615 -935
rect 1649 -969 1665 -935
rect 1599 -1000 1665 -969
rect 1695 969 1761 1000
rect 1695 935 1711 969
rect 1745 935 1761 969
rect 1695 901 1761 935
rect 1695 867 1711 901
rect 1745 867 1761 901
rect 1695 833 1761 867
rect 1695 799 1711 833
rect 1745 799 1761 833
rect 1695 765 1761 799
rect 1695 731 1711 765
rect 1745 731 1761 765
rect 1695 697 1761 731
rect 1695 663 1711 697
rect 1745 663 1761 697
rect 1695 629 1761 663
rect 1695 595 1711 629
rect 1745 595 1761 629
rect 1695 561 1761 595
rect 1695 527 1711 561
rect 1745 527 1761 561
rect 1695 493 1761 527
rect 1695 459 1711 493
rect 1745 459 1761 493
rect 1695 425 1761 459
rect 1695 391 1711 425
rect 1745 391 1761 425
rect 1695 357 1761 391
rect 1695 323 1711 357
rect 1745 323 1761 357
rect 1695 289 1761 323
rect 1695 255 1711 289
rect 1745 255 1761 289
rect 1695 221 1761 255
rect 1695 187 1711 221
rect 1745 187 1761 221
rect 1695 153 1761 187
rect 1695 119 1711 153
rect 1745 119 1761 153
rect 1695 85 1761 119
rect 1695 51 1711 85
rect 1745 51 1761 85
rect 1695 17 1761 51
rect 1695 -17 1711 17
rect 1745 -17 1761 17
rect 1695 -51 1761 -17
rect 1695 -85 1711 -51
rect 1745 -85 1761 -51
rect 1695 -119 1761 -85
rect 1695 -153 1711 -119
rect 1745 -153 1761 -119
rect 1695 -187 1761 -153
rect 1695 -221 1711 -187
rect 1745 -221 1761 -187
rect 1695 -255 1761 -221
rect 1695 -289 1711 -255
rect 1745 -289 1761 -255
rect 1695 -323 1761 -289
rect 1695 -357 1711 -323
rect 1745 -357 1761 -323
rect 1695 -391 1761 -357
rect 1695 -425 1711 -391
rect 1745 -425 1761 -391
rect 1695 -459 1761 -425
rect 1695 -493 1711 -459
rect 1745 -493 1761 -459
rect 1695 -527 1761 -493
rect 1695 -561 1711 -527
rect 1745 -561 1761 -527
rect 1695 -595 1761 -561
rect 1695 -629 1711 -595
rect 1745 -629 1761 -595
rect 1695 -663 1761 -629
rect 1695 -697 1711 -663
rect 1745 -697 1761 -663
rect 1695 -731 1761 -697
rect 1695 -765 1711 -731
rect 1745 -765 1761 -731
rect 1695 -799 1761 -765
rect 1695 -833 1711 -799
rect 1745 -833 1761 -799
rect 1695 -867 1761 -833
rect 1695 -901 1711 -867
rect 1745 -901 1761 -867
rect 1695 -935 1761 -901
rect 1695 -969 1711 -935
rect 1745 -969 1761 -935
rect 1695 -1000 1761 -969
rect 1791 969 1857 1000
rect 1791 935 1807 969
rect 1841 935 1857 969
rect 1791 901 1857 935
rect 1791 867 1807 901
rect 1841 867 1857 901
rect 1791 833 1857 867
rect 1791 799 1807 833
rect 1841 799 1857 833
rect 1791 765 1857 799
rect 1791 731 1807 765
rect 1841 731 1857 765
rect 1791 697 1857 731
rect 1791 663 1807 697
rect 1841 663 1857 697
rect 1791 629 1857 663
rect 1791 595 1807 629
rect 1841 595 1857 629
rect 1791 561 1857 595
rect 1791 527 1807 561
rect 1841 527 1857 561
rect 1791 493 1857 527
rect 1791 459 1807 493
rect 1841 459 1857 493
rect 1791 425 1857 459
rect 1791 391 1807 425
rect 1841 391 1857 425
rect 1791 357 1857 391
rect 1791 323 1807 357
rect 1841 323 1857 357
rect 1791 289 1857 323
rect 1791 255 1807 289
rect 1841 255 1857 289
rect 1791 221 1857 255
rect 1791 187 1807 221
rect 1841 187 1857 221
rect 1791 153 1857 187
rect 1791 119 1807 153
rect 1841 119 1857 153
rect 1791 85 1857 119
rect 1791 51 1807 85
rect 1841 51 1857 85
rect 1791 17 1857 51
rect 1791 -17 1807 17
rect 1841 -17 1857 17
rect 1791 -51 1857 -17
rect 1791 -85 1807 -51
rect 1841 -85 1857 -51
rect 1791 -119 1857 -85
rect 1791 -153 1807 -119
rect 1841 -153 1857 -119
rect 1791 -187 1857 -153
rect 1791 -221 1807 -187
rect 1841 -221 1857 -187
rect 1791 -255 1857 -221
rect 1791 -289 1807 -255
rect 1841 -289 1857 -255
rect 1791 -323 1857 -289
rect 1791 -357 1807 -323
rect 1841 -357 1857 -323
rect 1791 -391 1857 -357
rect 1791 -425 1807 -391
rect 1841 -425 1857 -391
rect 1791 -459 1857 -425
rect 1791 -493 1807 -459
rect 1841 -493 1857 -459
rect 1791 -527 1857 -493
rect 1791 -561 1807 -527
rect 1841 -561 1857 -527
rect 1791 -595 1857 -561
rect 1791 -629 1807 -595
rect 1841 -629 1857 -595
rect 1791 -663 1857 -629
rect 1791 -697 1807 -663
rect 1841 -697 1857 -663
rect 1791 -731 1857 -697
rect 1791 -765 1807 -731
rect 1841 -765 1857 -731
rect 1791 -799 1857 -765
rect 1791 -833 1807 -799
rect 1841 -833 1857 -799
rect 1791 -867 1857 -833
rect 1791 -901 1807 -867
rect 1841 -901 1857 -867
rect 1791 -935 1857 -901
rect 1791 -969 1807 -935
rect 1841 -969 1857 -935
rect 1791 -1000 1857 -969
rect 1887 969 1953 1000
rect 1887 935 1903 969
rect 1937 935 1953 969
rect 1887 901 1953 935
rect 1887 867 1903 901
rect 1937 867 1953 901
rect 1887 833 1953 867
rect 1887 799 1903 833
rect 1937 799 1953 833
rect 1887 765 1953 799
rect 1887 731 1903 765
rect 1937 731 1953 765
rect 1887 697 1953 731
rect 1887 663 1903 697
rect 1937 663 1953 697
rect 1887 629 1953 663
rect 1887 595 1903 629
rect 1937 595 1953 629
rect 1887 561 1953 595
rect 1887 527 1903 561
rect 1937 527 1953 561
rect 1887 493 1953 527
rect 1887 459 1903 493
rect 1937 459 1953 493
rect 1887 425 1953 459
rect 1887 391 1903 425
rect 1937 391 1953 425
rect 1887 357 1953 391
rect 1887 323 1903 357
rect 1937 323 1953 357
rect 1887 289 1953 323
rect 1887 255 1903 289
rect 1937 255 1953 289
rect 1887 221 1953 255
rect 1887 187 1903 221
rect 1937 187 1953 221
rect 1887 153 1953 187
rect 1887 119 1903 153
rect 1937 119 1953 153
rect 1887 85 1953 119
rect 1887 51 1903 85
rect 1937 51 1953 85
rect 1887 17 1953 51
rect 1887 -17 1903 17
rect 1937 -17 1953 17
rect 1887 -51 1953 -17
rect 1887 -85 1903 -51
rect 1937 -85 1953 -51
rect 1887 -119 1953 -85
rect 1887 -153 1903 -119
rect 1937 -153 1953 -119
rect 1887 -187 1953 -153
rect 1887 -221 1903 -187
rect 1937 -221 1953 -187
rect 1887 -255 1953 -221
rect 1887 -289 1903 -255
rect 1937 -289 1953 -255
rect 1887 -323 1953 -289
rect 1887 -357 1903 -323
rect 1937 -357 1953 -323
rect 1887 -391 1953 -357
rect 1887 -425 1903 -391
rect 1937 -425 1953 -391
rect 1887 -459 1953 -425
rect 1887 -493 1903 -459
rect 1937 -493 1953 -459
rect 1887 -527 1953 -493
rect 1887 -561 1903 -527
rect 1937 -561 1953 -527
rect 1887 -595 1953 -561
rect 1887 -629 1903 -595
rect 1937 -629 1953 -595
rect 1887 -663 1953 -629
rect 1887 -697 1903 -663
rect 1937 -697 1953 -663
rect 1887 -731 1953 -697
rect 1887 -765 1903 -731
rect 1937 -765 1953 -731
rect 1887 -799 1953 -765
rect 1887 -833 1903 -799
rect 1937 -833 1953 -799
rect 1887 -867 1953 -833
rect 1887 -901 1903 -867
rect 1937 -901 1953 -867
rect 1887 -935 1953 -901
rect 1887 -969 1903 -935
rect 1937 -969 1953 -935
rect 1887 -1000 1953 -969
rect 1983 969 2049 1000
rect 1983 935 1999 969
rect 2033 935 2049 969
rect 1983 901 2049 935
rect 1983 867 1999 901
rect 2033 867 2049 901
rect 1983 833 2049 867
rect 1983 799 1999 833
rect 2033 799 2049 833
rect 1983 765 2049 799
rect 1983 731 1999 765
rect 2033 731 2049 765
rect 1983 697 2049 731
rect 1983 663 1999 697
rect 2033 663 2049 697
rect 1983 629 2049 663
rect 1983 595 1999 629
rect 2033 595 2049 629
rect 1983 561 2049 595
rect 1983 527 1999 561
rect 2033 527 2049 561
rect 1983 493 2049 527
rect 1983 459 1999 493
rect 2033 459 2049 493
rect 1983 425 2049 459
rect 1983 391 1999 425
rect 2033 391 2049 425
rect 1983 357 2049 391
rect 1983 323 1999 357
rect 2033 323 2049 357
rect 1983 289 2049 323
rect 1983 255 1999 289
rect 2033 255 2049 289
rect 1983 221 2049 255
rect 1983 187 1999 221
rect 2033 187 2049 221
rect 1983 153 2049 187
rect 1983 119 1999 153
rect 2033 119 2049 153
rect 1983 85 2049 119
rect 1983 51 1999 85
rect 2033 51 2049 85
rect 1983 17 2049 51
rect 1983 -17 1999 17
rect 2033 -17 2049 17
rect 1983 -51 2049 -17
rect 1983 -85 1999 -51
rect 2033 -85 2049 -51
rect 1983 -119 2049 -85
rect 1983 -153 1999 -119
rect 2033 -153 2049 -119
rect 1983 -187 2049 -153
rect 1983 -221 1999 -187
rect 2033 -221 2049 -187
rect 1983 -255 2049 -221
rect 1983 -289 1999 -255
rect 2033 -289 2049 -255
rect 1983 -323 2049 -289
rect 1983 -357 1999 -323
rect 2033 -357 2049 -323
rect 1983 -391 2049 -357
rect 1983 -425 1999 -391
rect 2033 -425 2049 -391
rect 1983 -459 2049 -425
rect 1983 -493 1999 -459
rect 2033 -493 2049 -459
rect 1983 -527 2049 -493
rect 1983 -561 1999 -527
rect 2033 -561 2049 -527
rect 1983 -595 2049 -561
rect 1983 -629 1999 -595
rect 2033 -629 2049 -595
rect 1983 -663 2049 -629
rect 1983 -697 1999 -663
rect 2033 -697 2049 -663
rect 1983 -731 2049 -697
rect 1983 -765 1999 -731
rect 2033 -765 2049 -731
rect 1983 -799 2049 -765
rect 1983 -833 1999 -799
rect 2033 -833 2049 -799
rect 1983 -867 2049 -833
rect 1983 -901 1999 -867
rect 2033 -901 2049 -867
rect 1983 -935 2049 -901
rect 1983 -969 1999 -935
rect 2033 -969 2049 -935
rect 1983 -1000 2049 -969
rect 2079 969 2145 1000
rect 2079 935 2095 969
rect 2129 935 2145 969
rect 2079 901 2145 935
rect 2079 867 2095 901
rect 2129 867 2145 901
rect 2079 833 2145 867
rect 2079 799 2095 833
rect 2129 799 2145 833
rect 2079 765 2145 799
rect 2079 731 2095 765
rect 2129 731 2145 765
rect 2079 697 2145 731
rect 2079 663 2095 697
rect 2129 663 2145 697
rect 2079 629 2145 663
rect 2079 595 2095 629
rect 2129 595 2145 629
rect 2079 561 2145 595
rect 2079 527 2095 561
rect 2129 527 2145 561
rect 2079 493 2145 527
rect 2079 459 2095 493
rect 2129 459 2145 493
rect 2079 425 2145 459
rect 2079 391 2095 425
rect 2129 391 2145 425
rect 2079 357 2145 391
rect 2079 323 2095 357
rect 2129 323 2145 357
rect 2079 289 2145 323
rect 2079 255 2095 289
rect 2129 255 2145 289
rect 2079 221 2145 255
rect 2079 187 2095 221
rect 2129 187 2145 221
rect 2079 153 2145 187
rect 2079 119 2095 153
rect 2129 119 2145 153
rect 2079 85 2145 119
rect 2079 51 2095 85
rect 2129 51 2145 85
rect 2079 17 2145 51
rect 2079 -17 2095 17
rect 2129 -17 2145 17
rect 2079 -51 2145 -17
rect 2079 -85 2095 -51
rect 2129 -85 2145 -51
rect 2079 -119 2145 -85
rect 2079 -153 2095 -119
rect 2129 -153 2145 -119
rect 2079 -187 2145 -153
rect 2079 -221 2095 -187
rect 2129 -221 2145 -187
rect 2079 -255 2145 -221
rect 2079 -289 2095 -255
rect 2129 -289 2145 -255
rect 2079 -323 2145 -289
rect 2079 -357 2095 -323
rect 2129 -357 2145 -323
rect 2079 -391 2145 -357
rect 2079 -425 2095 -391
rect 2129 -425 2145 -391
rect 2079 -459 2145 -425
rect 2079 -493 2095 -459
rect 2129 -493 2145 -459
rect 2079 -527 2145 -493
rect 2079 -561 2095 -527
rect 2129 -561 2145 -527
rect 2079 -595 2145 -561
rect 2079 -629 2095 -595
rect 2129 -629 2145 -595
rect 2079 -663 2145 -629
rect 2079 -697 2095 -663
rect 2129 -697 2145 -663
rect 2079 -731 2145 -697
rect 2079 -765 2095 -731
rect 2129 -765 2145 -731
rect 2079 -799 2145 -765
rect 2079 -833 2095 -799
rect 2129 -833 2145 -799
rect 2079 -867 2145 -833
rect 2079 -901 2095 -867
rect 2129 -901 2145 -867
rect 2079 -935 2145 -901
rect 2079 -969 2095 -935
rect 2129 -969 2145 -935
rect 2079 -1000 2145 -969
rect 2175 969 2241 1000
rect 2175 935 2191 969
rect 2225 935 2241 969
rect 2175 901 2241 935
rect 2175 867 2191 901
rect 2225 867 2241 901
rect 2175 833 2241 867
rect 2175 799 2191 833
rect 2225 799 2241 833
rect 2175 765 2241 799
rect 2175 731 2191 765
rect 2225 731 2241 765
rect 2175 697 2241 731
rect 2175 663 2191 697
rect 2225 663 2241 697
rect 2175 629 2241 663
rect 2175 595 2191 629
rect 2225 595 2241 629
rect 2175 561 2241 595
rect 2175 527 2191 561
rect 2225 527 2241 561
rect 2175 493 2241 527
rect 2175 459 2191 493
rect 2225 459 2241 493
rect 2175 425 2241 459
rect 2175 391 2191 425
rect 2225 391 2241 425
rect 2175 357 2241 391
rect 2175 323 2191 357
rect 2225 323 2241 357
rect 2175 289 2241 323
rect 2175 255 2191 289
rect 2225 255 2241 289
rect 2175 221 2241 255
rect 2175 187 2191 221
rect 2225 187 2241 221
rect 2175 153 2241 187
rect 2175 119 2191 153
rect 2225 119 2241 153
rect 2175 85 2241 119
rect 2175 51 2191 85
rect 2225 51 2241 85
rect 2175 17 2241 51
rect 2175 -17 2191 17
rect 2225 -17 2241 17
rect 2175 -51 2241 -17
rect 2175 -85 2191 -51
rect 2225 -85 2241 -51
rect 2175 -119 2241 -85
rect 2175 -153 2191 -119
rect 2225 -153 2241 -119
rect 2175 -187 2241 -153
rect 2175 -221 2191 -187
rect 2225 -221 2241 -187
rect 2175 -255 2241 -221
rect 2175 -289 2191 -255
rect 2225 -289 2241 -255
rect 2175 -323 2241 -289
rect 2175 -357 2191 -323
rect 2225 -357 2241 -323
rect 2175 -391 2241 -357
rect 2175 -425 2191 -391
rect 2225 -425 2241 -391
rect 2175 -459 2241 -425
rect 2175 -493 2191 -459
rect 2225 -493 2241 -459
rect 2175 -527 2241 -493
rect 2175 -561 2191 -527
rect 2225 -561 2241 -527
rect 2175 -595 2241 -561
rect 2175 -629 2191 -595
rect 2225 -629 2241 -595
rect 2175 -663 2241 -629
rect 2175 -697 2191 -663
rect 2225 -697 2241 -663
rect 2175 -731 2241 -697
rect 2175 -765 2191 -731
rect 2225 -765 2241 -731
rect 2175 -799 2241 -765
rect 2175 -833 2191 -799
rect 2225 -833 2241 -799
rect 2175 -867 2241 -833
rect 2175 -901 2191 -867
rect 2225 -901 2241 -867
rect 2175 -935 2241 -901
rect 2175 -969 2191 -935
rect 2225 -969 2241 -935
rect 2175 -1000 2241 -969
rect 2271 969 2337 1000
rect 2271 935 2287 969
rect 2321 935 2337 969
rect 2271 901 2337 935
rect 2271 867 2287 901
rect 2321 867 2337 901
rect 2271 833 2337 867
rect 2271 799 2287 833
rect 2321 799 2337 833
rect 2271 765 2337 799
rect 2271 731 2287 765
rect 2321 731 2337 765
rect 2271 697 2337 731
rect 2271 663 2287 697
rect 2321 663 2337 697
rect 2271 629 2337 663
rect 2271 595 2287 629
rect 2321 595 2337 629
rect 2271 561 2337 595
rect 2271 527 2287 561
rect 2321 527 2337 561
rect 2271 493 2337 527
rect 2271 459 2287 493
rect 2321 459 2337 493
rect 2271 425 2337 459
rect 2271 391 2287 425
rect 2321 391 2337 425
rect 2271 357 2337 391
rect 2271 323 2287 357
rect 2321 323 2337 357
rect 2271 289 2337 323
rect 2271 255 2287 289
rect 2321 255 2337 289
rect 2271 221 2337 255
rect 2271 187 2287 221
rect 2321 187 2337 221
rect 2271 153 2337 187
rect 2271 119 2287 153
rect 2321 119 2337 153
rect 2271 85 2337 119
rect 2271 51 2287 85
rect 2321 51 2337 85
rect 2271 17 2337 51
rect 2271 -17 2287 17
rect 2321 -17 2337 17
rect 2271 -51 2337 -17
rect 2271 -85 2287 -51
rect 2321 -85 2337 -51
rect 2271 -119 2337 -85
rect 2271 -153 2287 -119
rect 2321 -153 2337 -119
rect 2271 -187 2337 -153
rect 2271 -221 2287 -187
rect 2321 -221 2337 -187
rect 2271 -255 2337 -221
rect 2271 -289 2287 -255
rect 2321 -289 2337 -255
rect 2271 -323 2337 -289
rect 2271 -357 2287 -323
rect 2321 -357 2337 -323
rect 2271 -391 2337 -357
rect 2271 -425 2287 -391
rect 2321 -425 2337 -391
rect 2271 -459 2337 -425
rect 2271 -493 2287 -459
rect 2321 -493 2337 -459
rect 2271 -527 2337 -493
rect 2271 -561 2287 -527
rect 2321 -561 2337 -527
rect 2271 -595 2337 -561
rect 2271 -629 2287 -595
rect 2321 -629 2337 -595
rect 2271 -663 2337 -629
rect 2271 -697 2287 -663
rect 2321 -697 2337 -663
rect 2271 -731 2337 -697
rect 2271 -765 2287 -731
rect 2321 -765 2337 -731
rect 2271 -799 2337 -765
rect 2271 -833 2287 -799
rect 2321 -833 2337 -799
rect 2271 -867 2337 -833
rect 2271 -901 2287 -867
rect 2321 -901 2337 -867
rect 2271 -935 2337 -901
rect 2271 -969 2287 -935
rect 2321 -969 2337 -935
rect 2271 -1000 2337 -969
rect 2367 969 2433 1000
rect 2367 935 2383 969
rect 2417 935 2433 969
rect 2367 901 2433 935
rect 2367 867 2383 901
rect 2417 867 2433 901
rect 2367 833 2433 867
rect 2367 799 2383 833
rect 2417 799 2433 833
rect 2367 765 2433 799
rect 2367 731 2383 765
rect 2417 731 2433 765
rect 2367 697 2433 731
rect 2367 663 2383 697
rect 2417 663 2433 697
rect 2367 629 2433 663
rect 2367 595 2383 629
rect 2417 595 2433 629
rect 2367 561 2433 595
rect 2367 527 2383 561
rect 2417 527 2433 561
rect 2367 493 2433 527
rect 2367 459 2383 493
rect 2417 459 2433 493
rect 2367 425 2433 459
rect 2367 391 2383 425
rect 2417 391 2433 425
rect 2367 357 2433 391
rect 2367 323 2383 357
rect 2417 323 2433 357
rect 2367 289 2433 323
rect 2367 255 2383 289
rect 2417 255 2433 289
rect 2367 221 2433 255
rect 2367 187 2383 221
rect 2417 187 2433 221
rect 2367 153 2433 187
rect 2367 119 2383 153
rect 2417 119 2433 153
rect 2367 85 2433 119
rect 2367 51 2383 85
rect 2417 51 2433 85
rect 2367 17 2433 51
rect 2367 -17 2383 17
rect 2417 -17 2433 17
rect 2367 -51 2433 -17
rect 2367 -85 2383 -51
rect 2417 -85 2433 -51
rect 2367 -119 2433 -85
rect 2367 -153 2383 -119
rect 2417 -153 2433 -119
rect 2367 -187 2433 -153
rect 2367 -221 2383 -187
rect 2417 -221 2433 -187
rect 2367 -255 2433 -221
rect 2367 -289 2383 -255
rect 2417 -289 2433 -255
rect 2367 -323 2433 -289
rect 2367 -357 2383 -323
rect 2417 -357 2433 -323
rect 2367 -391 2433 -357
rect 2367 -425 2383 -391
rect 2417 -425 2433 -391
rect 2367 -459 2433 -425
rect 2367 -493 2383 -459
rect 2417 -493 2433 -459
rect 2367 -527 2433 -493
rect 2367 -561 2383 -527
rect 2417 -561 2433 -527
rect 2367 -595 2433 -561
rect 2367 -629 2383 -595
rect 2417 -629 2433 -595
rect 2367 -663 2433 -629
rect 2367 -697 2383 -663
rect 2417 -697 2433 -663
rect 2367 -731 2433 -697
rect 2367 -765 2383 -731
rect 2417 -765 2433 -731
rect 2367 -799 2433 -765
rect 2367 -833 2383 -799
rect 2417 -833 2433 -799
rect 2367 -867 2433 -833
rect 2367 -901 2383 -867
rect 2417 -901 2433 -867
rect 2367 -935 2433 -901
rect 2367 -969 2383 -935
rect 2417 -969 2433 -935
rect 2367 -1000 2433 -969
rect 2463 969 2529 1000
rect 2463 935 2479 969
rect 2513 935 2529 969
rect 2463 901 2529 935
rect 2463 867 2479 901
rect 2513 867 2529 901
rect 2463 833 2529 867
rect 2463 799 2479 833
rect 2513 799 2529 833
rect 2463 765 2529 799
rect 2463 731 2479 765
rect 2513 731 2529 765
rect 2463 697 2529 731
rect 2463 663 2479 697
rect 2513 663 2529 697
rect 2463 629 2529 663
rect 2463 595 2479 629
rect 2513 595 2529 629
rect 2463 561 2529 595
rect 2463 527 2479 561
rect 2513 527 2529 561
rect 2463 493 2529 527
rect 2463 459 2479 493
rect 2513 459 2529 493
rect 2463 425 2529 459
rect 2463 391 2479 425
rect 2513 391 2529 425
rect 2463 357 2529 391
rect 2463 323 2479 357
rect 2513 323 2529 357
rect 2463 289 2529 323
rect 2463 255 2479 289
rect 2513 255 2529 289
rect 2463 221 2529 255
rect 2463 187 2479 221
rect 2513 187 2529 221
rect 2463 153 2529 187
rect 2463 119 2479 153
rect 2513 119 2529 153
rect 2463 85 2529 119
rect 2463 51 2479 85
rect 2513 51 2529 85
rect 2463 17 2529 51
rect 2463 -17 2479 17
rect 2513 -17 2529 17
rect 2463 -51 2529 -17
rect 2463 -85 2479 -51
rect 2513 -85 2529 -51
rect 2463 -119 2529 -85
rect 2463 -153 2479 -119
rect 2513 -153 2529 -119
rect 2463 -187 2529 -153
rect 2463 -221 2479 -187
rect 2513 -221 2529 -187
rect 2463 -255 2529 -221
rect 2463 -289 2479 -255
rect 2513 -289 2529 -255
rect 2463 -323 2529 -289
rect 2463 -357 2479 -323
rect 2513 -357 2529 -323
rect 2463 -391 2529 -357
rect 2463 -425 2479 -391
rect 2513 -425 2529 -391
rect 2463 -459 2529 -425
rect 2463 -493 2479 -459
rect 2513 -493 2529 -459
rect 2463 -527 2529 -493
rect 2463 -561 2479 -527
rect 2513 -561 2529 -527
rect 2463 -595 2529 -561
rect 2463 -629 2479 -595
rect 2513 -629 2529 -595
rect 2463 -663 2529 -629
rect 2463 -697 2479 -663
rect 2513 -697 2529 -663
rect 2463 -731 2529 -697
rect 2463 -765 2479 -731
rect 2513 -765 2529 -731
rect 2463 -799 2529 -765
rect 2463 -833 2479 -799
rect 2513 -833 2529 -799
rect 2463 -867 2529 -833
rect 2463 -901 2479 -867
rect 2513 -901 2529 -867
rect 2463 -935 2529 -901
rect 2463 -969 2479 -935
rect 2513 -969 2529 -935
rect 2463 -1000 2529 -969
rect 2559 969 2625 1000
rect 2559 935 2575 969
rect 2609 935 2625 969
rect 2559 901 2625 935
rect 2559 867 2575 901
rect 2609 867 2625 901
rect 2559 833 2625 867
rect 2559 799 2575 833
rect 2609 799 2625 833
rect 2559 765 2625 799
rect 2559 731 2575 765
rect 2609 731 2625 765
rect 2559 697 2625 731
rect 2559 663 2575 697
rect 2609 663 2625 697
rect 2559 629 2625 663
rect 2559 595 2575 629
rect 2609 595 2625 629
rect 2559 561 2625 595
rect 2559 527 2575 561
rect 2609 527 2625 561
rect 2559 493 2625 527
rect 2559 459 2575 493
rect 2609 459 2625 493
rect 2559 425 2625 459
rect 2559 391 2575 425
rect 2609 391 2625 425
rect 2559 357 2625 391
rect 2559 323 2575 357
rect 2609 323 2625 357
rect 2559 289 2625 323
rect 2559 255 2575 289
rect 2609 255 2625 289
rect 2559 221 2625 255
rect 2559 187 2575 221
rect 2609 187 2625 221
rect 2559 153 2625 187
rect 2559 119 2575 153
rect 2609 119 2625 153
rect 2559 85 2625 119
rect 2559 51 2575 85
rect 2609 51 2625 85
rect 2559 17 2625 51
rect 2559 -17 2575 17
rect 2609 -17 2625 17
rect 2559 -51 2625 -17
rect 2559 -85 2575 -51
rect 2609 -85 2625 -51
rect 2559 -119 2625 -85
rect 2559 -153 2575 -119
rect 2609 -153 2625 -119
rect 2559 -187 2625 -153
rect 2559 -221 2575 -187
rect 2609 -221 2625 -187
rect 2559 -255 2625 -221
rect 2559 -289 2575 -255
rect 2609 -289 2625 -255
rect 2559 -323 2625 -289
rect 2559 -357 2575 -323
rect 2609 -357 2625 -323
rect 2559 -391 2625 -357
rect 2559 -425 2575 -391
rect 2609 -425 2625 -391
rect 2559 -459 2625 -425
rect 2559 -493 2575 -459
rect 2609 -493 2625 -459
rect 2559 -527 2625 -493
rect 2559 -561 2575 -527
rect 2609 -561 2625 -527
rect 2559 -595 2625 -561
rect 2559 -629 2575 -595
rect 2609 -629 2625 -595
rect 2559 -663 2625 -629
rect 2559 -697 2575 -663
rect 2609 -697 2625 -663
rect 2559 -731 2625 -697
rect 2559 -765 2575 -731
rect 2609 -765 2625 -731
rect 2559 -799 2625 -765
rect 2559 -833 2575 -799
rect 2609 -833 2625 -799
rect 2559 -867 2625 -833
rect 2559 -901 2575 -867
rect 2609 -901 2625 -867
rect 2559 -935 2625 -901
rect 2559 -969 2575 -935
rect 2609 -969 2625 -935
rect 2559 -1000 2625 -969
rect 2655 969 2721 1000
rect 2655 935 2671 969
rect 2705 935 2721 969
rect 2655 901 2721 935
rect 2655 867 2671 901
rect 2705 867 2721 901
rect 2655 833 2721 867
rect 2655 799 2671 833
rect 2705 799 2721 833
rect 2655 765 2721 799
rect 2655 731 2671 765
rect 2705 731 2721 765
rect 2655 697 2721 731
rect 2655 663 2671 697
rect 2705 663 2721 697
rect 2655 629 2721 663
rect 2655 595 2671 629
rect 2705 595 2721 629
rect 2655 561 2721 595
rect 2655 527 2671 561
rect 2705 527 2721 561
rect 2655 493 2721 527
rect 2655 459 2671 493
rect 2705 459 2721 493
rect 2655 425 2721 459
rect 2655 391 2671 425
rect 2705 391 2721 425
rect 2655 357 2721 391
rect 2655 323 2671 357
rect 2705 323 2721 357
rect 2655 289 2721 323
rect 2655 255 2671 289
rect 2705 255 2721 289
rect 2655 221 2721 255
rect 2655 187 2671 221
rect 2705 187 2721 221
rect 2655 153 2721 187
rect 2655 119 2671 153
rect 2705 119 2721 153
rect 2655 85 2721 119
rect 2655 51 2671 85
rect 2705 51 2721 85
rect 2655 17 2721 51
rect 2655 -17 2671 17
rect 2705 -17 2721 17
rect 2655 -51 2721 -17
rect 2655 -85 2671 -51
rect 2705 -85 2721 -51
rect 2655 -119 2721 -85
rect 2655 -153 2671 -119
rect 2705 -153 2721 -119
rect 2655 -187 2721 -153
rect 2655 -221 2671 -187
rect 2705 -221 2721 -187
rect 2655 -255 2721 -221
rect 2655 -289 2671 -255
rect 2705 -289 2721 -255
rect 2655 -323 2721 -289
rect 2655 -357 2671 -323
rect 2705 -357 2721 -323
rect 2655 -391 2721 -357
rect 2655 -425 2671 -391
rect 2705 -425 2721 -391
rect 2655 -459 2721 -425
rect 2655 -493 2671 -459
rect 2705 -493 2721 -459
rect 2655 -527 2721 -493
rect 2655 -561 2671 -527
rect 2705 -561 2721 -527
rect 2655 -595 2721 -561
rect 2655 -629 2671 -595
rect 2705 -629 2721 -595
rect 2655 -663 2721 -629
rect 2655 -697 2671 -663
rect 2705 -697 2721 -663
rect 2655 -731 2721 -697
rect 2655 -765 2671 -731
rect 2705 -765 2721 -731
rect 2655 -799 2721 -765
rect 2655 -833 2671 -799
rect 2705 -833 2721 -799
rect 2655 -867 2721 -833
rect 2655 -901 2671 -867
rect 2705 -901 2721 -867
rect 2655 -935 2721 -901
rect 2655 -969 2671 -935
rect 2705 -969 2721 -935
rect 2655 -1000 2721 -969
rect 2751 969 2817 1000
rect 2751 935 2767 969
rect 2801 935 2817 969
rect 2751 901 2817 935
rect 2751 867 2767 901
rect 2801 867 2817 901
rect 2751 833 2817 867
rect 2751 799 2767 833
rect 2801 799 2817 833
rect 2751 765 2817 799
rect 2751 731 2767 765
rect 2801 731 2817 765
rect 2751 697 2817 731
rect 2751 663 2767 697
rect 2801 663 2817 697
rect 2751 629 2817 663
rect 2751 595 2767 629
rect 2801 595 2817 629
rect 2751 561 2817 595
rect 2751 527 2767 561
rect 2801 527 2817 561
rect 2751 493 2817 527
rect 2751 459 2767 493
rect 2801 459 2817 493
rect 2751 425 2817 459
rect 2751 391 2767 425
rect 2801 391 2817 425
rect 2751 357 2817 391
rect 2751 323 2767 357
rect 2801 323 2817 357
rect 2751 289 2817 323
rect 2751 255 2767 289
rect 2801 255 2817 289
rect 2751 221 2817 255
rect 2751 187 2767 221
rect 2801 187 2817 221
rect 2751 153 2817 187
rect 2751 119 2767 153
rect 2801 119 2817 153
rect 2751 85 2817 119
rect 2751 51 2767 85
rect 2801 51 2817 85
rect 2751 17 2817 51
rect 2751 -17 2767 17
rect 2801 -17 2817 17
rect 2751 -51 2817 -17
rect 2751 -85 2767 -51
rect 2801 -85 2817 -51
rect 2751 -119 2817 -85
rect 2751 -153 2767 -119
rect 2801 -153 2817 -119
rect 2751 -187 2817 -153
rect 2751 -221 2767 -187
rect 2801 -221 2817 -187
rect 2751 -255 2817 -221
rect 2751 -289 2767 -255
rect 2801 -289 2817 -255
rect 2751 -323 2817 -289
rect 2751 -357 2767 -323
rect 2801 -357 2817 -323
rect 2751 -391 2817 -357
rect 2751 -425 2767 -391
rect 2801 -425 2817 -391
rect 2751 -459 2817 -425
rect 2751 -493 2767 -459
rect 2801 -493 2817 -459
rect 2751 -527 2817 -493
rect 2751 -561 2767 -527
rect 2801 -561 2817 -527
rect 2751 -595 2817 -561
rect 2751 -629 2767 -595
rect 2801 -629 2817 -595
rect 2751 -663 2817 -629
rect 2751 -697 2767 -663
rect 2801 -697 2817 -663
rect 2751 -731 2817 -697
rect 2751 -765 2767 -731
rect 2801 -765 2817 -731
rect 2751 -799 2817 -765
rect 2751 -833 2767 -799
rect 2801 -833 2817 -799
rect 2751 -867 2817 -833
rect 2751 -901 2767 -867
rect 2801 -901 2817 -867
rect 2751 -935 2817 -901
rect 2751 -969 2767 -935
rect 2801 -969 2817 -935
rect 2751 -1000 2817 -969
rect 2847 969 2913 1000
rect 2847 935 2863 969
rect 2897 935 2913 969
rect 2847 901 2913 935
rect 2847 867 2863 901
rect 2897 867 2913 901
rect 2847 833 2913 867
rect 2847 799 2863 833
rect 2897 799 2913 833
rect 2847 765 2913 799
rect 2847 731 2863 765
rect 2897 731 2913 765
rect 2847 697 2913 731
rect 2847 663 2863 697
rect 2897 663 2913 697
rect 2847 629 2913 663
rect 2847 595 2863 629
rect 2897 595 2913 629
rect 2847 561 2913 595
rect 2847 527 2863 561
rect 2897 527 2913 561
rect 2847 493 2913 527
rect 2847 459 2863 493
rect 2897 459 2913 493
rect 2847 425 2913 459
rect 2847 391 2863 425
rect 2897 391 2913 425
rect 2847 357 2913 391
rect 2847 323 2863 357
rect 2897 323 2913 357
rect 2847 289 2913 323
rect 2847 255 2863 289
rect 2897 255 2913 289
rect 2847 221 2913 255
rect 2847 187 2863 221
rect 2897 187 2913 221
rect 2847 153 2913 187
rect 2847 119 2863 153
rect 2897 119 2913 153
rect 2847 85 2913 119
rect 2847 51 2863 85
rect 2897 51 2913 85
rect 2847 17 2913 51
rect 2847 -17 2863 17
rect 2897 -17 2913 17
rect 2847 -51 2913 -17
rect 2847 -85 2863 -51
rect 2897 -85 2913 -51
rect 2847 -119 2913 -85
rect 2847 -153 2863 -119
rect 2897 -153 2913 -119
rect 2847 -187 2913 -153
rect 2847 -221 2863 -187
rect 2897 -221 2913 -187
rect 2847 -255 2913 -221
rect 2847 -289 2863 -255
rect 2897 -289 2913 -255
rect 2847 -323 2913 -289
rect 2847 -357 2863 -323
rect 2897 -357 2913 -323
rect 2847 -391 2913 -357
rect 2847 -425 2863 -391
rect 2897 -425 2913 -391
rect 2847 -459 2913 -425
rect 2847 -493 2863 -459
rect 2897 -493 2913 -459
rect 2847 -527 2913 -493
rect 2847 -561 2863 -527
rect 2897 -561 2913 -527
rect 2847 -595 2913 -561
rect 2847 -629 2863 -595
rect 2897 -629 2913 -595
rect 2847 -663 2913 -629
rect 2847 -697 2863 -663
rect 2897 -697 2913 -663
rect 2847 -731 2913 -697
rect 2847 -765 2863 -731
rect 2897 -765 2913 -731
rect 2847 -799 2913 -765
rect 2847 -833 2863 -799
rect 2897 -833 2913 -799
rect 2847 -867 2913 -833
rect 2847 -901 2863 -867
rect 2897 -901 2913 -867
rect 2847 -935 2913 -901
rect 2847 -969 2863 -935
rect 2897 -969 2913 -935
rect 2847 -1000 2913 -969
rect 2943 969 3009 1000
rect 2943 935 2959 969
rect 2993 935 3009 969
rect 2943 901 3009 935
rect 2943 867 2959 901
rect 2993 867 3009 901
rect 2943 833 3009 867
rect 2943 799 2959 833
rect 2993 799 3009 833
rect 2943 765 3009 799
rect 2943 731 2959 765
rect 2993 731 3009 765
rect 2943 697 3009 731
rect 2943 663 2959 697
rect 2993 663 3009 697
rect 2943 629 3009 663
rect 2943 595 2959 629
rect 2993 595 3009 629
rect 2943 561 3009 595
rect 2943 527 2959 561
rect 2993 527 3009 561
rect 2943 493 3009 527
rect 2943 459 2959 493
rect 2993 459 3009 493
rect 2943 425 3009 459
rect 2943 391 2959 425
rect 2993 391 3009 425
rect 2943 357 3009 391
rect 2943 323 2959 357
rect 2993 323 3009 357
rect 2943 289 3009 323
rect 2943 255 2959 289
rect 2993 255 3009 289
rect 2943 221 3009 255
rect 2943 187 2959 221
rect 2993 187 3009 221
rect 2943 153 3009 187
rect 2943 119 2959 153
rect 2993 119 3009 153
rect 2943 85 3009 119
rect 2943 51 2959 85
rect 2993 51 3009 85
rect 2943 17 3009 51
rect 2943 -17 2959 17
rect 2993 -17 3009 17
rect 2943 -51 3009 -17
rect 2943 -85 2959 -51
rect 2993 -85 3009 -51
rect 2943 -119 3009 -85
rect 2943 -153 2959 -119
rect 2993 -153 3009 -119
rect 2943 -187 3009 -153
rect 2943 -221 2959 -187
rect 2993 -221 3009 -187
rect 2943 -255 3009 -221
rect 2943 -289 2959 -255
rect 2993 -289 3009 -255
rect 2943 -323 3009 -289
rect 2943 -357 2959 -323
rect 2993 -357 3009 -323
rect 2943 -391 3009 -357
rect 2943 -425 2959 -391
rect 2993 -425 3009 -391
rect 2943 -459 3009 -425
rect 2943 -493 2959 -459
rect 2993 -493 3009 -459
rect 2943 -527 3009 -493
rect 2943 -561 2959 -527
rect 2993 -561 3009 -527
rect 2943 -595 3009 -561
rect 2943 -629 2959 -595
rect 2993 -629 3009 -595
rect 2943 -663 3009 -629
rect 2943 -697 2959 -663
rect 2993 -697 3009 -663
rect 2943 -731 3009 -697
rect 2943 -765 2959 -731
rect 2993 -765 3009 -731
rect 2943 -799 3009 -765
rect 2943 -833 2959 -799
rect 2993 -833 3009 -799
rect 2943 -867 3009 -833
rect 2943 -901 2959 -867
rect 2993 -901 3009 -867
rect 2943 -935 3009 -901
rect 2943 -969 2959 -935
rect 2993 -969 3009 -935
rect 2943 -1000 3009 -969
rect 3039 969 3105 1000
rect 3039 935 3055 969
rect 3089 935 3105 969
rect 3039 901 3105 935
rect 3039 867 3055 901
rect 3089 867 3105 901
rect 3039 833 3105 867
rect 3039 799 3055 833
rect 3089 799 3105 833
rect 3039 765 3105 799
rect 3039 731 3055 765
rect 3089 731 3105 765
rect 3039 697 3105 731
rect 3039 663 3055 697
rect 3089 663 3105 697
rect 3039 629 3105 663
rect 3039 595 3055 629
rect 3089 595 3105 629
rect 3039 561 3105 595
rect 3039 527 3055 561
rect 3089 527 3105 561
rect 3039 493 3105 527
rect 3039 459 3055 493
rect 3089 459 3105 493
rect 3039 425 3105 459
rect 3039 391 3055 425
rect 3089 391 3105 425
rect 3039 357 3105 391
rect 3039 323 3055 357
rect 3089 323 3105 357
rect 3039 289 3105 323
rect 3039 255 3055 289
rect 3089 255 3105 289
rect 3039 221 3105 255
rect 3039 187 3055 221
rect 3089 187 3105 221
rect 3039 153 3105 187
rect 3039 119 3055 153
rect 3089 119 3105 153
rect 3039 85 3105 119
rect 3039 51 3055 85
rect 3089 51 3105 85
rect 3039 17 3105 51
rect 3039 -17 3055 17
rect 3089 -17 3105 17
rect 3039 -51 3105 -17
rect 3039 -85 3055 -51
rect 3089 -85 3105 -51
rect 3039 -119 3105 -85
rect 3039 -153 3055 -119
rect 3089 -153 3105 -119
rect 3039 -187 3105 -153
rect 3039 -221 3055 -187
rect 3089 -221 3105 -187
rect 3039 -255 3105 -221
rect 3039 -289 3055 -255
rect 3089 -289 3105 -255
rect 3039 -323 3105 -289
rect 3039 -357 3055 -323
rect 3089 -357 3105 -323
rect 3039 -391 3105 -357
rect 3039 -425 3055 -391
rect 3089 -425 3105 -391
rect 3039 -459 3105 -425
rect 3039 -493 3055 -459
rect 3089 -493 3105 -459
rect 3039 -527 3105 -493
rect 3039 -561 3055 -527
rect 3089 -561 3105 -527
rect 3039 -595 3105 -561
rect 3039 -629 3055 -595
rect 3089 -629 3105 -595
rect 3039 -663 3105 -629
rect 3039 -697 3055 -663
rect 3089 -697 3105 -663
rect 3039 -731 3105 -697
rect 3039 -765 3055 -731
rect 3089 -765 3105 -731
rect 3039 -799 3105 -765
rect 3039 -833 3055 -799
rect 3089 -833 3105 -799
rect 3039 -867 3105 -833
rect 3039 -901 3055 -867
rect 3089 -901 3105 -867
rect 3039 -935 3105 -901
rect 3039 -969 3055 -935
rect 3089 -969 3105 -935
rect 3039 -1000 3105 -969
rect 3135 969 3201 1000
rect 3135 935 3151 969
rect 3185 935 3201 969
rect 3135 901 3201 935
rect 3135 867 3151 901
rect 3185 867 3201 901
rect 3135 833 3201 867
rect 3135 799 3151 833
rect 3185 799 3201 833
rect 3135 765 3201 799
rect 3135 731 3151 765
rect 3185 731 3201 765
rect 3135 697 3201 731
rect 3135 663 3151 697
rect 3185 663 3201 697
rect 3135 629 3201 663
rect 3135 595 3151 629
rect 3185 595 3201 629
rect 3135 561 3201 595
rect 3135 527 3151 561
rect 3185 527 3201 561
rect 3135 493 3201 527
rect 3135 459 3151 493
rect 3185 459 3201 493
rect 3135 425 3201 459
rect 3135 391 3151 425
rect 3185 391 3201 425
rect 3135 357 3201 391
rect 3135 323 3151 357
rect 3185 323 3201 357
rect 3135 289 3201 323
rect 3135 255 3151 289
rect 3185 255 3201 289
rect 3135 221 3201 255
rect 3135 187 3151 221
rect 3185 187 3201 221
rect 3135 153 3201 187
rect 3135 119 3151 153
rect 3185 119 3201 153
rect 3135 85 3201 119
rect 3135 51 3151 85
rect 3185 51 3201 85
rect 3135 17 3201 51
rect 3135 -17 3151 17
rect 3185 -17 3201 17
rect 3135 -51 3201 -17
rect 3135 -85 3151 -51
rect 3185 -85 3201 -51
rect 3135 -119 3201 -85
rect 3135 -153 3151 -119
rect 3185 -153 3201 -119
rect 3135 -187 3201 -153
rect 3135 -221 3151 -187
rect 3185 -221 3201 -187
rect 3135 -255 3201 -221
rect 3135 -289 3151 -255
rect 3185 -289 3201 -255
rect 3135 -323 3201 -289
rect 3135 -357 3151 -323
rect 3185 -357 3201 -323
rect 3135 -391 3201 -357
rect 3135 -425 3151 -391
rect 3185 -425 3201 -391
rect 3135 -459 3201 -425
rect 3135 -493 3151 -459
rect 3185 -493 3201 -459
rect 3135 -527 3201 -493
rect 3135 -561 3151 -527
rect 3185 -561 3201 -527
rect 3135 -595 3201 -561
rect 3135 -629 3151 -595
rect 3185 -629 3201 -595
rect 3135 -663 3201 -629
rect 3135 -697 3151 -663
rect 3185 -697 3201 -663
rect 3135 -731 3201 -697
rect 3135 -765 3151 -731
rect 3185 -765 3201 -731
rect 3135 -799 3201 -765
rect 3135 -833 3151 -799
rect 3185 -833 3201 -799
rect 3135 -867 3201 -833
rect 3135 -901 3151 -867
rect 3185 -901 3201 -867
rect 3135 -935 3201 -901
rect 3135 -969 3151 -935
rect 3185 -969 3201 -935
rect 3135 -1000 3201 -969
rect 3231 969 3297 1000
rect 3231 935 3247 969
rect 3281 935 3297 969
rect 3231 901 3297 935
rect 3231 867 3247 901
rect 3281 867 3297 901
rect 3231 833 3297 867
rect 3231 799 3247 833
rect 3281 799 3297 833
rect 3231 765 3297 799
rect 3231 731 3247 765
rect 3281 731 3297 765
rect 3231 697 3297 731
rect 3231 663 3247 697
rect 3281 663 3297 697
rect 3231 629 3297 663
rect 3231 595 3247 629
rect 3281 595 3297 629
rect 3231 561 3297 595
rect 3231 527 3247 561
rect 3281 527 3297 561
rect 3231 493 3297 527
rect 3231 459 3247 493
rect 3281 459 3297 493
rect 3231 425 3297 459
rect 3231 391 3247 425
rect 3281 391 3297 425
rect 3231 357 3297 391
rect 3231 323 3247 357
rect 3281 323 3297 357
rect 3231 289 3297 323
rect 3231 255 3247 289
rect 3281 255 3297 289
rect 3231 221 3297 255
rect 3231 187 3247 221
rect 3281 187 3297 221
rect 3231 153 3297 187
rect 3231 119 3247 153
rect 3281 119 3297 153
rect 3231 85 3297 119
rect 3231 51 3247 85
rect 3281 51 3297 85
rect 3231 17 3297 51
rect 3231 -17 3247 17
rect 3281 -17 3297 17
rect 3231 -51 3297 -17
rect 3231 -85 3247 -51
rect 3281 -85 3297 -51
rect 3231 -119 3297 -85
rect 3231 -153 3247 -119
rect 3281 -153 3297 -119
rect 3231 -187 3297 -153
rect 3231 -221 3247 -187
rect 3281 -221 3297 -187
rect 3231 -255 3297 -221
rect 3231 -289 3247 -255
rect 3281 -289 3297 -255
rect 3231 -323 3297 -289
rect 3231 -357 3247 -323
rect 3281 -357 3297 -323
rect 3231 -391 3297 -357
rect 3231 -425 3247 -391
rect 3281 -425 3297 -391
rect 3231 -459 3297 -425
rect 3231 -493 3247 -459
rect 3281 -493 3297 -459
rect 3231 -527 3297 -493
rect 3231 -561 3247 -527
rect 3281 -561 3297 -527
rect 3231 -595 3297 -561
rect 3231 -629 3247 -595
rect 3281 -629 3297 -595
rect 3231 -663 3297 -629
rect 3231 -697 3247 -663
rect 3281 -697 3297 -663
rect 3231 -731 3297 -697
rect 3231 -765 3247 -731
rect 3281 -765 3297 -731
rect 3231 -799 3297 -765
rect 3231 -833 3247 -799
rect 3281 -833 3297 -799
rect 3231 -867 3297 -833
rect 3231 -901 3247 -867
rect 3281 -901 3297 -867
rect 3231 -935 3297 -901
rect 3231 -969 3247 -935
rect 3281 -969 3297 -935
rect 3231 -1000 3297 -969
rect 3327 969 3393 1000
rect 3327 935 3343 969
rect 3377 935 3393 969
rect 3327 901 3393 935
rect 3327 867 3343 901
rect 3377 867 3393 901
rect 3327 833 3393 867
rect 3327 799 3343 833
rect 3377 799 3393 833
rect 3327 765 3393 799
rect 3327 731 3343 765
rect 3377 731 3393 765
rect 3327 697 3393 731
rect 3327 663 3343 697
rect 3377 663 3393 697
rect 3327 629 3393 663
rect 3327 595 3343 629
rect 3377 595 3393 629
rect 3327 561 3393 595
rect 3327 527 3343 561
rect 3377 527 3393 561
rect 3327 493 3393 527
rect 3327 459 3343 493
rect 3377 459 3393 493
rect 3327 425 3393 459
rect 3327 391 3343 425
rect 3377 391 3393 425
rect 3327 357 3393 391
rect 3327 323 3343 357
rect 3377 323 3393 357
rect 3327 289 3393 323
rect 3327 255 3343 289
rect 3377 255 3393 289
rect 3327 221 3393 255
rect 3327 187 3343 221
rect 3377 187 3393 221
rect 3327 153 3393 187
rect 3327 119 3343 153
rect 3377 119 3393 153
rect 3327 85 3393 119
rect 3327 51 3343 85
rect 3377 51 3393 85
rect 3327 17 3393 51
rect 3327 -17 3343 17
rect 3377 -17 3393 17
rect 3327 -51 3393 -17
rect 3327 -85 3343 -51
rect 3377 -85 3393 -51
rect 3327 -119 3393 -85
rect 3327 -153 3343 -119
rect 3377 -153 3393 -119
rect 3327 -187 3393 -153
rect 3327 -221 3343 -187
rect 3377 -221 3393 -187
rect 3327 -255 3393 -221
rect 3327 -289 3343 -255
rect 3377 -289 3393 -255
rect 3327 -323 3393 -289
rect 3327 -357 3343 -323
rect 3377 -357 3393 -323
rect 3327 -391 3393 -357
rect 3327 -425 3343 -391
rect 3377 -425 3393 -391
rect 3327 -459 3393 -425
rect 3327 -493 3343 -459
rect 3377 -493 3393 -459
rect 3327 -527 3393 -493
rect 3327 -561 3343 -527
rect 3377 -561 3393 -527
rect 3327 -595 3393 -561
rect 3327 -629 3343 -595
rect 3377 -629 3393 -595
rect 3327 -663 3393 -629
rect 3327 -697 3343 -663
rect 3377 -697 3393 -663
rect 3327 -731 3393 -697
rect 3327 -765 3343 -731
rect 3377 -765 3393 -731
rect 3327 -799 3393 -765
rect 3327 -833 3343 -799
rect 3377 -833 3393 -799
rect 3327 -867 3393 -833
rect 3327 -901 3343 -867
rect 3377 -901 3393 -867
rect 3327 -935 3393 -901
rect 3327 -969 3343 -935
rect 3377 -969 3393 -935
rect 3327 -1000 3393 -969
rect 3423 969 3489 1000
rect 3423 935 3439 969
rect 3473 935 3489 969
rect 3423 901 3489 935
rect 3423 867 3439 901
rect 3473 867 3489 901
rect 3423 833 3489 867
rect 3423 799 3439 833
rect 3473 799 3489 833
rect 3423 765 3489 799
rect 3423 731 3439 765
rect 3473 731 3489 765
rect 3423 697 3489 731
rect 3423 663 3439 697
rect 3473 663 3489 697
rect 3423 629 3489 663
rect 3423 595 3439 629
rect 3473 595 3489 629
rect 3423 561 3489 595
rect 3423 527 3439 561
rect 3473 527 3489 561
rect 3423 493 3489 527
rect 3423 459 3439 493
rect 3473 459 3489 493
rect 3423 425 3489 459
rect 3423 391 3439 425
rect 3473 391 3489 425
rect 3423 357 3489 391
rect 3423 323 3439 357
rect 3473 323 3489 357
rect 3423 289 3489 323
rect 3423 255 3439 289
rect 3473 255 3489 289
rect 3423 221 3489 255
rect 3423 187 3439 221
rect 3473 187 3489 221
rect 3423 153 3489 187
rect 3423 119 3439 153
rect 3473 119 3489 153
rect 3423 85 3489 119
rect 3423 51 3439 85
rect 3473 51 3489 85
rect 3423 17 3489 51
rect 3423 -17 3439 17
rect 3473 -17 3489 17
rect 3423 -51 3489 -17
rect 3423 -85 3439 -51
rect 3473 -85 3489 -51
rect 3423 -119 3489 -85
rect 3423 -153 3439 -119
rect 3473 -153 3489 -119
rect 3423 -187 3489 -153
rect 3423 -221 3439 -187
rect 3473 -221 3489 -187
rect 3423 -255 3489 -221
rect 3423 -289 3439 -255
rect 3473 -289 3489 -255
rect 3423 -323 3489 -289
rect 3423 -357 3439 -323
rect 3473 -357 3489 -323
rect 3423 -391 3489 -357
rect 3423 -425 3439 -391
rect 3473 -425 3489 -391
rect 3423 -459 3489 -425
rect 3423 -493 3439 -459
rect 3473 -493 3489 -459
rect 3423 -527 3489 -493
rect 3423 -561 3439 -527
rect 3473 -561 3489 -527
rect 3423 -595 3489 -561
rect 3423 -629 3439 -595
rect 3473 -629 3489 -595
rect 3423 -663 3489 -629
rect 3423 -697 3439 -663
rect 3473 -697 3489 -663
rect 3423 -731 3489 -697
rect 3423 -765 3439 -731
rect 3473 -765 3489 -731
rect 3423 -799 3489 -765
rect 3423 -833 3439 -799
rect 3473 -833 3489 -799
rect 3423 -867 3489 -833
rect 3423 -901 3439 -867
rect 3473 -901 3489 -867
rect 3423 -935 3489 -901
rect 3423 -969 3439 -935
rect 3473 -969 3489 -935
rect 3423 -1000 3489 -969
rect 3519 969 3585 1000
rect 3519 935 3535 969
rect 3569 935 3585 969
rect 3519 901 3585 935
rect 3519 867 3535 901
rect 3569 867 3585 901
rect 3519 833 3585 867
rect 3519 799 3535 833
rect 3569 799 3585 833
rect 3519 765 3585 799
rect 3519 731 3535 765
rect 3569 731 3585 765
rect 3519 697 3585 731
rect 3519 663 3535 697
rect 3569 663 3585 697
rect 3519 629 3585 663
rect 3519 595 3535 629
rect 3569 595 3585 629
rect 3519 561 3585 595
rect 3519 527 3535 561
rect 3569 527 3585 561
rect 3519 493 3585 527
rect 3519 459 3535 493
rect 3569 459 3585 493
rect 3519 425 3585 459
rect 3519 391 3535 425
rect 3569 391 3585 425
rect 3519 357 3585 391
rect 3519 323 3535 357
rect 3569 323 3585 357
rect 3519 289 3585 323
rect 3519 255 3535 289
rect 3569 255 3585 289
rect 3519 221 3585 255
rect 3519 187 3535 221
rect 3569 187 3585 221
rect 3519 153 3585 187
rect 3519 119 3535 153
rect 3569 119 3585 153
rect 3519 85 3585 119
rect 3519 51 3535 85
rect 3569 51 3585 85
rect 3519 17 3585 51
rect 3519 -17 3535 17
rect 3569 -17 3585 17
rect 3519 -51 3585 -17
rect 3519 -85 3535 -51
rect 3569 -85 3585 -51
rect 3519 -119 3585 -85
rect 3519 -153 3535 -119
rect 3569 -153 3585 -119
rect 3519 -187 3585 -153
rect 3519 -221 3535 -187
rect 3569 -221 3585 -187
rect 3519 -255 3585 -221
rect 3519 -289 3535 -255
rect 3569 -289 3585 -255
rect 3519 -323 3585 -289
rect 3519 -357 3535 -323
rect 3569 -357 3585 -323
rect 3519 -391 3585 -357
rect 3519 -425 3535 -391
rect 3569 -425 3585 -391
rect 3519 -459 3585 -425
rect 3519 -493 3535 -459
rect 3569 -493 3585 -459
rect 3519 -527 3585 -493
rect 3519 -561 3535 -527
rect 3569 -561 3585 -527
rect 3519 -595 3585 -561
rect 3519 -629 3535 -595
rect 3569 -629 3585 -595
rect 3519 -663 3585 -629
rect 3519 -697 3535 -663
rect 3569 -697 3585 -663
rect 3519 -731 3585 -697
rect 3519 -765 3535 -731
rect 3569 -765 3585 -731
rect 3519 -799 3585 -765
rect 3519 -833 3535 -799
rect 3569 -833 3585 -799
rect 3519 -867 3585 -833
rect 3519 -901 3535 -867
rect 3569 -901 3585 -867
rect 3519 -935 3585 -901
rect 3519 -969 3535 -935
rect 3569 -969 3585 -935
rect 3519 -1000 3585 -969
rect 3615 969 3681 1000
rect 3615 935 3631 969
rect 3665 935 3681 969
rect 3615 901 3681 935
rect 3615 867 3631 901
rect 3665 867 3681 901
rect 3615 833 3681 867
rect 3615 799 3631 833
rect 3665 799 3681 833
rect 3615 765 3681 799
rect 3615 731 3631 765
rect 3665 731 3681 765
rect 3615 697 3681 731
rect 3615 663 3631 697
rect 3665 663 3681 697
rect 3615 629 3681 663
rect 3615 595 3631 629
rect 3665 595 3681 629
rect 3615 561 3681 595
rect 3615 527 3631 561
rect 3665 527 3681 561
rect 3615 493 3681 527
rect 3615 459 3631 493
rect 3665 459 3681 493
rect 3615 425 3681 459
rect 3615 391 3631 425
rect 3665 391 3681 425
rect 3615 357 3681 391
rect 3615 323 3631 357
rect 3665 323 3681 357
rect 3615 289 3681 323
rect 3615 255 3631 289
rect 3665 255 3681 289
rect 3615 221 3681 255
rect 3615 187 3631 221
rect 3665 187 3681 221
rect 3615 153 3681 187
rect 3615 119 3631 153
rect 3665 119 3681 153
rect 3615 85 3681 119
rect 3615 51 3631 85
rect 3665 51 3681 85
rect 3615 17 3681 51
rect 3615 -17 3631 17
rect 3665 -17 3681 17
rect 3615 -51 3681 -17
rect 3615 -85 3631 -51
rect 3665 -85 3681 -51
rect 3615 -119 3681 -85
rect 3615 -153 3631 -119
rect 3665 -153 3681 -119
rect 3615 -187 3681 -153
rect 3615 -221 3631 -187
rect 3665 -221 3681 -187
rect 3615 -255 3681 -221
rect 3615 -289 3631 -255
rect 3665 -289 3681 -255
rect 3615 -323 3681 -289
rect 3615 -357 3631 -323
rect 3665 -357 3681 -323
rect 3615 -391 3681 -357
rect 3615 -425 3631 -391
rect 3665 -425 3681 -391
rect 3615 -459 3681 -425
rect 3615 -493 3631 -459
rect 3665 -493 3681 -459
rect 3615 -527 3681 -493
rect 3615 -561 3631 -527
rect 3665 -561 3681 -527
rect 3615 -595 3681 -561
rect 3615 -629 3631 -595
rect 3665 -629 3681 -595
rect 3615 -663 3681 -629
rect 3615 -697 3631 -663
rect 3665 -697 3681 -663
rect 3615 -731 3681 -697
rect 3615 -765 3631 -731
rect 3665 -765 3681 -731
rect 3615 -799 3681 -765
rect 3615 -833 3631 -799
rect 3665 -833 3681 -799
rect 3615 -867 3681 -833
rect 3615 -901 3631 -867
rect 3665 -901 3681 -867
rect 3615 -935 3681 -901
rect 3615 -969 3631 -935
rect 3665 -969 3681 -935
rect 3615 -1000 3681 -969
rect 3711 969 3777 1000
rect 3711 935 3727 969
rect 3761 935 3777 969
rect 3711 901 3777 935
rect 3711 867 3727 901
rect 3761 867 3777 901
rect 3711 833 3777 867
rect 3711 799 3727 833
rect 3761 799 3777 833
rect 3711 765 3777 799
rect 3711 731 3727 765
rect 3761 731 3777 765
rect 3711 697 3777 731
rect 3711 663 3727 697
rect 3761 663 3777 697
rect 3711 629 3777 663
rect 3711 595 3727 629
rect 3761 595 3777 629
rect 3711 561 3777 595
rect 3711 527 3727 561
rect 3761 527 3777 561
rect 3711 493 3777 527
rect 3711 459 3727 493
rect 3761 459 3777 493
rect 3711 425 3777 459
rect 3711 391 3727 425
rect 3761 391 3777 425
rect 3711 357 3777 391
rect 3711 323 3727 357
rect 3761 323 3777 357
rect 3711 289 3777 323
rect 3711 255 3727 289
rect 3761 255 3777 289
rect 3711 221 3777 255
rect 3711 187 3727 221
rect 3761 187 3777 221
rect 3711 153 3777 187
rect 3711 119 3727 153
rect 3761 119 3777 153
rect 3711 85 3777 119
rect 3711 51 3727 85
rect 3761 51 3777 85
rect 3711 17 3777 51
rect 3711 -17 3727 17
rect 3761 -17 3777 17
rect 3711 -51 3777 -17
rect 3711 -85 3727 -51
rect 3761 -85 3777 -51
rect 3711 -119 3777 -85
rect 3711 -153 3727 -119
rect 3761 -153 3777 -119
rect 3711 -187 3777 -153
rect 3711 -221 3727 -187
rect 3761 -221 3777 -187
rect 3711 -255 3777 -221
rect 3711 -289 3727 -255
rect 3761 -289 3777 -255
rect 3711 -323 3777 -289
rect 3711 -357 3727 -323
rect 3761 -357 3777 -323
rect 3711 -391 3777 -357
rect 3711 -425 3727 -391
rect 3761 -425 3777 -391
rect 3711 -459 3777 -425
rect 3711 -493 3727 -459
rect 3761 -493 3777 -459
rect 3711 -527 3777 -493
rect 3711 -561 3727 -527
rect 3761 -561 3777 -527
rect 3711 -595 3777 -561
rect 3711 -629 3727 -595
rect 3761 -629 3777 -595
rect 3711 -663 3777 -629
rect 3711 -697 3727 -663
rect 3761 -697 3777 -663
rect 3711 -731 3777 -697
rect 3711 -765 3727 -731
rect 3761 -765 3777 -731
rect 3711 -799 3777 -765
rect 3711 -833 3727 -799
rect 3761 -833 3777 -799
rect 3711 -867 3777 -833
rect 3711 -901 3727 -867
rect 3761 -901 3777 -867
rect 3711 -935 3777 -901
rect 3711 -969 3727 -935
rect 3761 -969 3777 -935
rect 3711 -1000 3777 -969
rect 3807 969 3873 1000
rect 3807 935 3823 969
rect 3857 935 3873 969
rect 3807 901 3873 935
rect 3807 867 3823 901
rect 3857 867 3873 901
rect 3807 833 3873 867
rect 3807 799 3823 833
rect 3857 799 3873 833
rect 3807 765 3873 799
rect 3807 731 3823 765
rect 3857 731 3873 765
rect 3807 697 3873 731
rect 3807 663 3823 697
rect 3857 663 3873 697
rect 3807 629 3873 663
rect 3807 595 3823 629
rect 3857 595 3873 629
rect 3807 561 3873 595
rect 3807 527 3823 561
rect 3857 527 3873 561
rect 3807 493 3873 527
rect 3807 459 3823 493
rect 3857 459 3873 493
rect 3807 425 3873 459
rect 3807 391 3823 425
rect 3857 391 3873 425
rect 3807 357 3873 391
rect 3807 323 3823 357
rect 3857 323 3873 357
rect 3807 289 3873 323
rect 3807 255 3823 289
rect 3857 255 3873 289
rect 3807 221 3873 255
rect 3807 187 3823 221
rect 3857 187 3873 221
rect 3807 153 3873 187
rect 3807 119 3823 153
rect 3857 119 3873 153
rect 3807 85 3873 119
rect 3807 51 3823 85
rect 3857 51 3873 85
rect 3807 17 3873 51
rect 3807 -17 3823 17
rect 3857 -17 3873 17
rect 3807 -51 3873 -17
rect 3807 -85 3823 -51
rect 3857 -85 3873 -51
rect 3807 -119 3873 -85
rect 3807 -153 3823 -119
rect 3857 -153 3873 -119
rect 3807 -187 3873 -153
rect 3807 -221 3823 -187
rect 3857 -221 3873 -187
rect 3807 -255 3873 -221
rect 3807 -289 3823 -255
rect 3857 -289 3873 -255
rect 3807 -323 3873 -289
rect 3807 -357 3823 -323
rect 3857 -357 3873 -323
rect 3807 -391 3873 -357
rect 3807 -425 3823 -391
rect 3857 -425 3873 -391
rect 3807 -459 3873 -425
rect 3807 -493 3823 -459
rect 3857 -493 3873 -459
rect 3807 -527 3873 -493
rect 3807 -561 3823 -527
rect 3857 -561 3873 -527
rect 3807 -595 3873 -561
rect 3807 -629 3823 -595
rect 3857 -629 3873 -595
rect 3807 -663 3873 -629
rect 3807 -697 3823 -663
rect 3857 -697 3873 -663
rect 3807 -731 3873 -697
rect 3807 -765 3823 -731
rect 3857 -765 3873 -731
rect 3807 -799 3873 -765
rect 3807 -833 3823 -799
rect 3857 -833 3873 -799
rect 3807 -867 3873 -833
rect 3807 -901 3823 -867
rect 3857 -901 3873 -867
rect 3807 -935 3873 -901
rect 3807 -969 3823 -935
rect 3857 -969 3873 -935
rect 3807 -1000 3873 -969
rect 3903 969 3969 1000
rect 3903 935 3919 969
rect 3953 935 3969 969
rect 3903 901 3969 935
rect 3903 867 3919 901
rect 3953 867 3969 901
rect 3903 833 3969 867
rect 3903 799 3919 833
rect 3953 799 3969 833
rect 3903 765 3969 799
rect 3903 731 3919 765
rect 3953 731 3969 765
rect 3903 697 3969 731
rect 3903 663 3919 697
rect 3953 663 3969 697
rect 3903 629 3969 663
rect 3903 595 3919 629
rect 3953 595 3969 629
rect 3903 561 3969 595
rect 3903 527 3919 561
rect 3953 527 3969 561
rect 3903 493 3969 527
rect 3903 459 3919 493
rect 3953 459 3969 493
rect 3903 425 3969 459
rect 3903 391 3919 425
rect 3953 391 3969 425
rect 3903 357 3969 391
rect 3903 323 3919 357
rect 3953 323 3969 357
rect 3903 289 3969 323
rect 3903 255 3919 289
rect 3953 255 3969 289
rect 3903 221 3969 255
rect 3903 187 3919 221
rect 3953 187 3969 221
rect 3903 153 3969 187
rect 3903 119 3919 153
rect 3953 119 3969 153
rect 3903 85 3969 119
rect 3903 51 3919 85
rect 3953 51 3969 85
rect 3903 17 3969 51
rect 3903 -17 3919 17
rect 3953 -17 3969 17
rect 3903 -51 3969 -17
rect 3903 -85 3919 -51
rect 3953 -85 3969 -51
rect 3903 -119 3969 -85
rect 3903 -153 3919 -119
rect 3953 -153 3969 -119
rect 3903 -187 3969 -153
rect 3903 -221 3919 -187
rect 3953 -221 3969 -187
rect 3903 -255 3969 -221
rect 3903 -289 3919 -255
rect 3953 -289 3969 -255
rect 3903 -323 3969 -289
rect 3903 -357 3919 -323
rect 3953 -357 3969 -323
rect 3903 -391 3969 -357
rect 3903 -425 3919 -391
rect 3953 -425 3969 -391
rect 3903 -459 3969 -425
rect 3903 -493 3919 -459
rect 3953 -493 3969 -459
rect 3903 -527 3969 -493
rect 3903 -561 3919 -527
rect 3953 -561 3969 -527
rect 3903 -595 3969 -561
rect 3903 -629 3919 -595
rect 3953 -629 3969 -595
rect 3903 -663 3969 -629
rect 3903 -697 3919 -663
rect 3953 -697 3969 -663
rect 3903 -731 3969 -697
rect 3903 -765 3919 -731
rect 3953 -765 3969 -731
rect 3903 -799 3969 -765
rect 3903 -833 3919 -799
rect 3953 -833 3969 -799
rect 3903 -867 3969 -833
rect 3903 -901 3919 -867
rect 3953 -901 3969 -867
rect 3903 -935 3969 -901
rect 3903 -969 3919 -935
rect 3953 -969 3969 -935
rect 3903 -1000 3969 -969
rect 3999 969 4065 1000
rect 3999 935 4015 969
rect 4049 935 4065 969
rect 3999 901 4065 935
rect 3999 867 4015 901
rect 4049 867 4065 901
rect 3999 833 4065 867
rect 3999 799 4015 833
rect 4049 799 4065 833
rect 3999 765 4065 799
rect 3999 731 4015 765
rect 4049 731 4065 765
rect 3999 697 4065 731
rect 3999 663 4015 697
rect 4049 663 4065 697
rect 3999 629 4065 663
rect 3999 595 4015 629
rect 4049 595 4065 629
rect 3999 561 4065 595
rect 3999 527 4015 561
rect 4049 527 4065 561
rect 3999 493 4065 527
rect 3999 459 4015 493
rect 4049 459 4065 493
rect 3999 425 4065 459
rect 3999 391 4015 425
rect 4049 391 4065 425
rect 3999 357 4065 391
rect 3999 323 4015 357
rect 4049 323 4065 357
rect 3999 289 4065 323
rect 3999 255 4015 289
rect 4049 255 4065 289
rect 3999 221 4065 255
rect 3999 187 4015 221
rect 4049 187 4065 221
rect 3999 153 4065 187
rect 3999 119 4015 153
rect 4049 119 4065 153
rect 3999 85 4065 119
rect 3999 51 4015 85
rect 4049 51 4065 85
rect 3999 17 4065 51
rect 3999 -17 4015 17
rect 4049 -17 4065 17
rect 3999 -51 4065 -17
rect 3999 -85 4015 -51
rect 4049 -85 4065 -51
rect 3999 -119 4065 -85
rect 3999 -153 4015 -119
rect 4049 -153 4065 -119
rect 3999 -187 4065 -153
rect 3999 -221 4015 -187
rect 4049 -221 4065 -187
rect 3999 -255 4065 -221
rect 3999 -289 4015 -255
rect 4049 -289 4065 -255
rect 3999 -323 4065 -289
rect 3999 -357 4015 -323
rect 4049 -357 4065 -323
rect 3999 -391 4065 -357
rect 3999 -425 4015 -391
rect 4049 -425 4065 -391
rect 3999 -459 4065 -425
rect 3999 -493 4015 -459
rect 4049 -493 4065 -459
rect 3999 -527 4065 -493
rect 3999 -561 4015 -527
rect 4049 -561 4065 -527
rect 3999 -595 4065 -561
rect 3999 -629 4015 -595
rect 4049 -629 4065 -595
rect 3999 -663 4065 -629
rect 3999 -697 4015 -663
rect 4049 -697 4065 -663
rect 3999 -731 4065 -697
rect 3999 -765 4015 -731
rect 4049 -765 4065 -731
rect 3999 -799 4065 -765
rect 3999 -833 4015 -799
rect 4049 -833 4065 -799
rect 3999 -867 4065 -833
rect 3999 -901 4015 -867
rect 4049 -901 4065 -867
rect 3999 -935 4065 -901
rect 3999 -969 4015 -935
rect 4049 -969 4065 -935
rect 3999 -1000 4065 -969
rect 4095 969 4161 1000
rect 4095 935 4111 969
rect 4145 935 4161 969
rect 4095 901 4161 935
rect 4095 867 4111 901
rect 4145 867 4161 901
rect 4095 833 4161 867
rect 4095 799 4111 833
rect 4145 799 4161 833
rect 4095 765 4161 799
rect 4095 731 4111 765
rect 4145 731 4161 765
rect 4095 697 4161 731
rect 4095 663 4111 697
rect 4145 663 4161 697
rect 4095 629 4161 663
rect 4095 595 4111 629
rect 4145 595 4161 629
rect 4095 561 4161 595
rect 4095 527 4111 561
rect 4145 527 4161 561
rect 4095 493 4161 527
rect 4095 459 4111 493
rect 4145 459 4161 493
rect 4095 425 4161 459
rect 4095 391 4111 425
rect 4145 391 4161 425
rect 4095 357 4161 391
rect 4095 323 4111 357
rect 4145 323 4161 357
rect 4095 289 4161 323
rect 4095 255 4111 289
rect 4145 255 4161 289
rect 4095 221 4161 255
rect 4095 187 4111 221
rect 4145 187 4161 221
rect 4095 153 4161 187
rect 4095 119 4111 153
rect 4145 119 4161 153
rect 4095 85 4161 119
rect 4095 51 4111 85
rect 4145 51 4161 85
rect 4095 17 4161 51
rect 4095 -17 4111 17
rect 4145 -17 4161 17
rect 4095 -51 4161 -17
rect 4095 -85 4111 -51
rect 4145 -85 4161 -51
rect 4095 -119 4161 -85
rect 4095 -153 4111 -119
rect 4145 -153 4161 -119
rect 4095 -187 4161 -153
rect 4095 -221 4111 -187
rect 4145 -221 4161 -187
rect 4095 -255 4161 -221
rect 4095 -289 4111 -255
rect 4145 -289 4161 -255
rect 4095 -323 4161 -289
rect 4095 -357 4111 -323
rect 4145 -357 4161 -323
rect 4095 -391 4161 -357
rect 4095 -425 4111 -391
rect 4145 -425 4161 -391
rect 4095 -459 4161 -425
rect 4095 -493 4111 -459
rect 4145 -493 4161 -459
rect 4095 -527 4161 -493
rect 4095 -561 4111 -527
rect 4145 -561 4161 -527
rect 4095 -595 4161 -561
rect 4095 -629 4111 -595
rect 4145 -629 4161 -595
rect 4095 -663 4161 -629
rect 4095 -697 4111 -663
rect 4145 -697 4161 -663
rect 4095 -731 4161 -697
rect 4095 -765 4111 -731
rect 4145 -765 4161 -731
rect 4095 -799 4161 -765
rect 4095 -833 4111 -799
rect 4145 -833 4161 -799
rect 4095 -867 4161 -833
rect 4095 -901 4111 -867
rect 4145 -901 4161 -867
rect 4095 -935 4161 -901
rect 4095 -969 4111 -935
rect 4145 -969 4161 -935
rect 4095 -1000 4161 -969
rect 4191 969 4257 1000
rect 4191 935 4207 969
rect 4241 935 4257 969
rect 4191 901 4257 935
rect 4191 867 4207 901
rect 4241 867 4257 901
rect 4191 833 4257 867
rect 4191 799 4207 833
rect 4241 799 4257 833
rect 4191 765 4257 799
rect 4191 731 4207 765
rect 4241 731 4257 765
rect 4191 697 4257 731
rect 4191 663 4207 697
rect 4241 663 4257 697
rect 4191 629 4257 663
rect 4191 595 4207 629
rect 4241 595 4257 629
rect 4191 561 4257 595
rect 4191 527 4207 561
rect 4241 527 4257 561
rect 4191 493 4257 527
rect 4191 459 4207 493
rect 4241 459 4257 493
rect 4191 425 4257 459
rect 4191 391 4207 425
rect 4241 391 4257 425
rect 4191 357 4257 391
rect 4191 323 4207 357
rect 4241 323 4257 357
rect 4191 289 4257 323
rect 4191 255 4207 289
rect 4241 255 4257 289
rect 4191 221 4257 255
rect 4191 187 4207 221
rect 4241 187 4257 221
rect 4191 153 4257 187
rect 4191 119 4207 153
rect 4241 119 4257 153
rect 4191 85 4257 119
rect 4191 51 4207 85
rect 4241 51 4257 85
rect 4191 17 4257 51
rect 4191 -17 4207 17
rect 4241 -17 4257 17
rect 4191 -51 4257 -17
rect 4191 -85 4207 -51
rect 4241 -85 4257 -51
rect 4191 -119 4257 -85
rect 4191 -153 4207 -119
rect 4241 -153 4257 -119
rect 4191 -187 4257 -153
rect 4191 -221 4207 -187
rect 4241 -221 4257 -187
rect 4191 -255 4257 -221
rect 4191 -289 4207 -255
rect 4241 -289 4257 -255
rect 4191 -323 4257 -289
rect 4191 -357 4207 -323
rect 4241 -357 4257 -323
rect 4191 -391 4257 -357
rect 4191 -425 4207 -391
rect 4241 -425 4257 -391
rect 4191 -459 4257 -425
rect 4191 -493 4207 -459
rect 4241 -493 4257 -459
rect 4191 -527 4257 -493
rect 4191 -561 4207 -527
rect 4241 -561 4257 -527
rect 4191 -595 4257 -561
rect 4191 -629 4207 -595
rect 4241 -629 4257 -595
rect 4191 -663 4257 -629
rect 4191 -697 4207 -663
rect 4241 -697 4257 -663
rect 4191 -731 4257 -697
rect 4191 -765 4207 -731
rect 4241 -765 4257 -731
rect 4191 -799 4257 -765
rect 4191 -833 4207 -799
rect 4241 -833 4257 -799
rect 4191 -867 4257 -833
rect 4191 -901 4207 -867
rect 4241 -901 4257 -867
rect 4191 -935 4257 -901
rect 4191 -969 4207 -935
rect 4241 -969 4257 -935
rect 4191 -1000 4257 -969
rect 4287 969 4353 1000
rect 4287 935 4303 969
rect 4337 935 4353 969
rect 4287 901 4353 935
rect 4287 867 4303 901
rect 4337 867 4353 901
rect 4287 833 4353 867
rect 4287 799 4303 833
rect 4337 799 4353 833
rect 4287 765 4353 799
rect 4287 731 4303 765
rect 4337 731 4353 765
rect 4287 697 4353 731
rect 4287 663 4303 697
rect 4337 663 4353 697
rect 4287 629 4353 663
rect 4287 595 4303 629
rect 4337 595 4353 629
rect 4287 561 4353 595
rect 4287 527 4303 561
rect 4337 527 4353 561
rect 4287 493 4353 527
rect 4287 459 4303 493
rect 4337 459 4353 493
rect 4287 425 4353 459
rect 4287 391 4303 425
rect 4337 391 4353 425
rect 4287 357 4353 391
rect 4287 323 4303 357
rect 4337 323 4353 357
rect 4287 289 4353 323
rect 4287 255 4303 289
rect 4337 255 4353 289
rect 4287 221 4353 255
rect 4287 187 4303 221
rect 4337 187 4353 221
rect 4287 153 4353 187
rect 4287 119 4303 153
rect 4337 119 4353 153
rect 4287 85 4353 119
rect 4287 51 4303 85
rect 4337 51 4353 85
rect 4287 17 4353 51
rect 4287 -17 4303 17
rect 4337 -17 4353 17
rect 4287 -51 4353 -17
rect 4287 -85 4303 -51
rect 4337 -85 4353 -51
rect 4287 -119 4353 -85
rect 4287 -153 4303 -119
rect 4337 -153 4353 -119
rect 4287 -187 4353 -153
rect 4287 -221 4303 -187
rect 4337 -221 4353 -187
rect 4287 -255 4353 -221
rect 4287 -289 4303 -255
rect 4337 -289 4353 -255
rect 4287 -323 4353 -289
rect 4287 -357 4303 -323
rect 4337 -357 4353 -323
rect 4287 -391 4353 -357
rect 4287 -425 4303 -391
rect 4337 -425 4353 -391
rect 4287 -459 4353 -425
rect 4287 -493 4303 -459
rect 4337 -493 4353 -459
rect 4287 -527 4353 -493
rect 4287 -561 4303 -527
rect 4337 -561 4353 -527
rect 4287 -595 4353 -561
rect 4287 -629 4303 -595
rect 4337 -629 4353 -595
rect 4287 -663 4353 -629
rect 4287 -697 4303 -663
rect 4337 -697 4353 -663
rect 4287 -731 4353 -697
rect 4287 -765 4303 -731
rect 4337 -765 4353 -731
rect 4287 -799 4353 -765
rect 4287 -833 4303 -799
rect 4337 -833 4353 -799
rect 4287 -867 4353 -833
rect 4287 -901 4303 -867
rect 4337 -901 4353 -867
rect 4287 -935 4353 -901
rect 4287 -969 4303 -935
rect 4337 -969 4353 -935
rect 4287 -1000 4353 -969
rect 4383 969 4449 1000
rect 4383 935 4399 969
rect 4433 935 4449 969
rect 4383 901 4449 935
rect 4383 867 4399 901
rect 4433 867 4449 901
rect 4383 833 4449 867
rect 4383 799 4399 833
rect 4433 799 4449 833
rect 4383 765 4449 799
rect 4383 731 4399 765
rect 4433 731 4449 765
rect 4383 697 4449 731
rect 4383 663 4399 697
rect 4433 663 4449 697
rect 4383 629 4449 663
rect 4383 595 4399 629
rect 4433 595 4449 629
rect 4383 561 4449 595
rect 4383 527 4399 561
rect 4433 527 4449 561
rect 4383 493 4449 527
rect 4383 459 4399 493
rect 4433 459 4449 493
rect 4383 425 4449 459
rect 4383 391 4399 425
rect 4433 391 4449 425
rect 4383 357 4449 391
rect 4383 323 4399 357
rect 4433 323 4449 357
rect 4383 289 4449 323
rect 4383 255 4399 289
rect 4433 255 4449 289
rect 4383 221 4449 255
rect 4383 187 4399 221
rect 4433 187 4449 221
rect 4383 153 4449 187
rect 4383 119 4399 153
rect 4433 119 4449 153
rect 4383 85 4449 119
rect 4383 51 4399 85
rect 4433 51 4449 85
rect 4383 17 4449 51
rect 4383 -17 4399 17
rect 4433 -17 4449 17
rect 4383 -51 4449 -17
rect 4383 -85 4399 -51
rect 4433 -85 4449 -51
rect 4383 -119 4449 -85
rect 4383 -153 4399 -119
rect 4433 -153 4449 -119
rect 4383 -187 4449 -153
rect 4383 -221 4399 -187
rect 4433 -221 4449 -187
rect 4383 -255 4449 -221
rect 4383 -289 4399 -255
rect 4433 -289 4449 -255
rect 4383 -323 4449 -289
rect 4383 -357 4399 -323
rect 4433 -357 4449 -323
rect 4383 -391 4449 -357
rect 4383 -425 4399 -391
rect 4433 -425 4449 -391
rect 4383 -459 4449 -425
rect 4383 -493 4399 -459
rect 4433 -493 4449 -459
rect 4383 -527 4449 -493
rect 4383 -561 4399 -527
rect 4433 -561 4449 -527
rect 4383 -595 4449 -561
rect 4383 -629 4399 -595
rect 4433 -629 4449 -595
rect 4383 -663 4449 -629
rect 4383 -697 4399 -663
rect 4433 -697 4449 -663
rect 4383 -731 4449 -697
rect 4383 -765 4399 -731
rect 4433 -765 4449 -731
rect 4383 -799 4449 -765
rect 4383 -833 4399 -799
rect 4433 -833 4449 -799
rect 4383 -867 4449 -833
rect 4383 -901 4399 -867
rect 4433 -901 4449 -867
rect 4383 -935 4449 -901
rect 4383 -969 4399 -935
rect 4433 -969 4449 -935
rect 4383 -1000 4449 -969
rect 4479 969 4545 1000
rect 4479 935 4495 969
rect 4529 935 4545 969
rect 4479 901 4545 935
rect 4479 867 4495 901
rect 4529 867 4545 901
rect 4479 833 4545 867
rect 4479 799 4495 833
rect 4529 799 4545 833
rect 4479 765 4545 799
rect 4479 731 4495 765
rect 4529 731 4545 765
rect 4479 697 4545 731
rect 4479 663 4495 697
rect 4529 663 4545 697
rect 4479 629 4545 663
rect 4479 595 4495 629
rect 4529 595 4545 629
rect 4479 561 4545 595
rect 4479 527 4495 561
rect 4529 527 4545 561
rect 4479 493 4545 527
rect 4479 459 4495 493
rect 4529 459 4545 493
rect 4479 425 4545 459
rect 4479 391 4495 425
rect 4529 391 4545 425
rect 4479 357 4545 391
rect 4479 323 4495 357
rect 4529 323 4545 357
rect 4479 289 4545 323
rect 4479 255 4495 289
rect 4529 255 4545 289
rect 4479 221 4545 255
rect 4479 187 4495 221
rect 4529 187 4545 221
rect 4479 153 4545 187
rect 4479 119 4495 153
rect 4529 119 4545 153
rect 4479 85 4545 119
rect 4479 51 4495 85
rect 4529 51 4545 85
rect 4479 17 4545 51
rect 4479 -17 4495 17
rect 4529 -17 4545 17
rect 4479 -51 4545 -17
rect 4479 -85 4495 -51
rect 4529 -85 4545 -51
rect 4479 -119 4545 -85
rect 4479 -153 4495 -119
rect 4529 -153 4545 -119
rect 4479 -187 4545 -153
rect 4479 -221 4495 -187
rect 4529 -221 4545 -187
rect 4479 -255 4545 -221
rect 4479 -289 4495 -255
rect 4529 -289 4545 -255
rect 4479 -323 4545 -289
rect 4479 -357 4495 -323
rect 4529 -357 4545 -323
rect 4479 -391 4545 -357
rect 4479 -425 4495 -391
rect 4529 -425 4545 -391
rect 4479 -459 4545 -425
rect 4479 -493 4495 -459
rect 4529 -493 4545 -459
rect 4479 -527 4545 -493
rect 4479 -561 4495 -527
rect 4529 -561 4545 -527
rect 4479 -595 4545 -561
rect 4479 -629 4495 -595
rect 4529 -629 4545 -595
rect 4479 -663 4545 -629
rect 4479 -697 4495 -663
rect 4529 -697 4545 -663
rect 4479 -731 4545 -697
rect 4479 -765 4495 -731
rect 4529 -765 4545 -731
rect 4479 -799 4545 -765
rect 4479 -833 4495 -799
rect 4529 -833 4545 -799
rect 4479 -867 4545 -833
rect 4479 -901 4495 -867
rect 4529 -901 4545 -867
rect 4479 -935 4545 -901
rect 4479 -969 4495 -935
rect 4529 -969 4545 -935
rect 4479 -1000 4545 -969
rect 4575 969 4641 1000
rect 4575 935 4591 969
rect 4625 935 4641 969
rect 4575 901 4641 935
rect 4575 867 4591 901
rect 4625 867 4641 901
rect 4575 833 4641 867
rect 4575 799 4591 833
rect 4625 799 4641 833
rect 4575 765 4641 799
rect 4575 731 4591 765
rect 4625 731 4641 765
rect 4575 697 4641 731
rect 4575 663 4591 697
rect 4625 663 4641 697
rect 4575 629 4641 663
rect 4575 595 4591 629
rect 4625 595 4641 629
rect 4575 561 4641 595
rect 4575 527 4591 561
rect 4625 527 4641 561
rect 4575 493 4641 527
rect 4575 459 4591 493
rect 4625 459 4641 493
rect 4575 425 4641 459
rect 4575 391 4591 425
rect 4625 391 4641 425
rect 4575 357 4641 391
rect 4575 323 4591 357
rect 4625 323 4641 357
rect 4575 289 4641 323
rect 4575 255 4591 289
rect 4625 255 4641 289
rect 4575 221 4641 255
rect 4575 187 4591 221
rect 4625 187 4641 221
rect 4575 153 4641 187
rect 4575 119 4591 153
rect 4625 119 4641 153
rect 4575 85 4641 119
rect 4575 51 4591 85
rect 4625 51 4641 85
rect 4575 17 4641 51
rect 4575 -17 4591 17
rect 4625 -17 4641 17
rect 4575 -51 4641 -17
rect 4575 -85 4591 -51
rect 4625 -85 4641 -51
rect 4575 -119 4641 -85
rect 4575 -153 4591 -119
rect 4625 -153 4641 -119
rect 4575 -187 4641 -153
rect 4575 -221 4591 -187
rect 4625 -221 4641 -187
rect 4575 -255 4641 -221
rect 4575 -289 4591 -255
rect 4625 -289 4641 -255
rect 4575 -323 4641 -289
rect 4575 -357 4591 -323
rect 4625 -357 4641 -323
rect 4575 -391 4641 -357
rect 4575 -425 4591 -391
rect 4625 -425 4641 -391
rect 4575 -459 4641 -425
rect 4575 -493 4591 -459
rect 4625 -493 4641 -459
rect 4575 -527 4641 -493
rect 4575 -561 4591 -527
rect 4625 -561 4641 -527
rect 4575 -595 4641 -561
rect 4575 -629 4591 -595
rect 4625 -629 4641 -595
rect 4575 -663 4641 -629
rect 4575 -697 4591 -663
rect 4625 -697 4641 -663
rect 4575 -731 4641 -697
rect 4575 -765 4591 -731
rect 4625 -765 4641 -731
rect 4575 -799 4641 -765
rect 4575 -833 4591 -799
rect 4625 -833 4641 -799
rect 4575 -867 4641 -833
rect 4575 -901 4591 -867
rect 4625 -901 4641 -867
rect 4575 -935 4641 -901
rect 4575 -969 4591 -935
rect 4625 -969 4641 -935
rect 4575 -1000 4641 -969
rect 4671 969 4737 1000
rect 4671 935 4687 969
rect 4721 935 4737 969
rect 4671 901 4737 935
rect 4671 867 4687 901
rect 4721 867 4737 901
rect 4671 833 4737 867
rect 4671 799 4687 833
rect 4721 799 4737 833
rect 4671 765 4737 799
rect 4671 731 4687 765
rect 4721 731 4737 765
rect 4671 697 4737 731
rect 4671 663 4687 697
rect 4721 663 4737 697
rect 4671 629 4737 663
rect 4671 595 4687 629
rect 4721 595 4737 629
rect 4671 561 4737 595
rect 4671 527 4687 561
rect 4721 527 4737 561
rect 4671 493 4737 527
rect 4671 459 4687 493
rect 4721 459 4737 493
rect 4671 425 4737 459
rect 4671 391 4687 425
rect 4721 391 4737 425
rect 4671 357 4737 391
rect 4671 323 4687 357
rect 4721 323 4737 357
rect 4671 289 4737 323
rect 4671 255 4687 289
rect 4721 255 4737 289
rect 4671 221 4737 255
rect 4671 187 4687 221
rect 4721 187 4737 221
rect 4671 153 4737 187
rect 4671 119 4687 153
rect 4721 119 4737 153
rect 4671 85 4737 119
rect 4671 51 4687 85
rect 4721 51 4737 85
rect 4671 17 4737 51
rect 4671 -17 4687 17
rect 4721 -17 4737 17
rect 4671 -51 4737 -17
rect 4671 -85 4687 -51
rect 4721 -85 4737 -51
rect 4671 -119 4737 -85
rect 4671 -153 4687 -119
rect 4721 -153 4737 -119
rect 4671 -187 4737 -153
rect 4671 -221 4687 -187
rect 4721 -221 4737 -187
rect 4671 -255 4737 -221
rect 4671 -289 4687 -255
rect 4721 -289 4737 -255
rect 4671 -323 4737 -289
rect 4671 -357 4687 -323
rect 4721 -357 4737 -323
rect 4671 -391 4737 -357
rect 4671 -425 4687 -391
rect 4721 -425 4737 -391
rect 4671 -459 4737 -425
rect 4671 -493 4687 -459
rect 4721 -493 4737 -459
rect 4671 -527 4737 -493
rect 4671 -561 4687 -527
rect 4721 -561 4737 -527
rect 4671 -595 4737 -561
rect 4671 -629 4687 -595
rect 4721 -629 4737 -595
rect 4671 -663 4737 -629
rect 4671 -697 4687 -663
rect 4721 -697 4737 -663
rect 4671 -731 4737 -697
rect 4671 -765 4687 -731
rect 4721 -765 4737 -731
rect 4671 -799 4737 -765
rect 4671 -833 4687 -799
rect 4721 -833 4737 -799
rect 4671 -867 4737 -833
rect 4671 -901 4687 -867
rect 4721 -901 4737 -867
rect 4671 -935 4737 -901
rect 4671 -969 4687 -935
rect 4721 -969 4737 -935
rect 4671 -1000 4737 -969
rect 4767 969 4829 1000
rect 4767 935 4783 969
rect 4817 935 4829 969
rect 4767 901 4829 935
rect 4767 867 4783 901
rect 4817 867 4829 901
rect 4767 833 4829 867
rect 4767 799 4783 833
rect 4817 799 4829 833
rect 4767 765 4829 799
rect 4767 731 4783 765
rect 4817 731 4829 765
rect 4767 697 4829 731
rect 4767 663 4783 697
rect 4817 663 4829 697
rect 4767 629 4829 663
rect 4767 595 4783 629
rect 4817 595 4829 629
rect 4767 561 4829 595
rect 4767 527 4783 561
rect 4817 527 4829 561
rect 4767 493 4829 527
rect 4767 459 4783 493
rect 4817 459 4829 493
rect 4767 425 4829 459
rect 4767 391 4783 425
rect 4817 391 4829 425
rect 4767 357 4829 391
rect 4767 323 4783 357
rect 4817 323 4829 357
rect 4767 289 4829 323
rect 4767 255 4783 289
rect 4817 255 4829 289
rect 4767 221 4829 255
rect 4767 187 4783 221
rect 4817 187 4829 221
rect 4767 153 4829 187
rect 4767 119 4783 153
rect 4817 119 4829 153
rect 4767 85 4829 119
rect 4767 51 4783 85
rect 4817 51 4829 85
rect 4767 17 4829 51
rect 4767 -17 4783 17
rect 4817 -17 4829 17
rect 4767 -51 4829 -17
rect 4767 -85 4783 -51
rect 4817 -85 4829 -51
rect 4767 -119 4829 -85
rect 4767 -153 4783 -119
rect 4817 -153 4829 -119
rect 4767 -187 4829 -153
rect 4767 -221 4783 -187
rect 4817 -221 4829 -187
rect 4767 -255 4829 -221
rect 4767 -289 4783 -255
rect 4817 -289 4829 -255
rect 4767 -323 4829 -289
rect 4767 -357 4783 -323
rect 4817 -357 4829 -323
rect 4767 -391 4829 -357
rect 4767 -425 4783 -391
rect 4817 -425 4829 -391
rect 4767 -459 4829 -425
rect 4767 -493 4783 -459
rect 4817 -493 4829 -459
rect 4767 -527 4829 -493
rect 4767 -561 4783 -527
rect 4817 -561 4829 -527
rect 4767 -595 4829 -561
rect 4767 -629 4783 -595
rect 4817 -629 4829 -595
rect 4767 -663 4829 -629
rect 4767 -697 4783 -663
rect 4817 -697 4829 -663
rect 4767 -731 4829 -697
rect 4767 -765 4783 -731
rect 4817 -765 4829 -731
rect 4767 -799 4829 -765
rect 4767 -833 4783 -799
rect 4817 -833 4829 -799
rect 4767 -867 4829 -833
rect 4767 -901 4783 -867
rect 4817 -901 4829 -867
rect 4767 -935 4829 -901
rect 4767 -969 4783 -935
rect 4817 -969 4829 -935
rect 4767 -1000 4829 -969
<< ndiffc >>
rect -4817 935 -4783 969
rect -4817 867 -4783 901
rect -4817 799 -4783 833
rect -4817 731 -4783 765
rect -4817 663 -4783 697
rect -4817 595 -4783 629
rect -4817 527 -4783 561
rect -4817 459 -4783 493
rect -4817 391 -4783 425
rect -4817 323 -4783 357
rect -4817 255 -4783 289
rect -4817 187 -4783 221
rect -4817 119 -4783 153
rect -4817 51 -4783 85
rect -4817 -17 -4783 17
rect -4817 -85 -4783 -51
rect -4817 -153 -4783 -119
rect -4817 -221 -4783 -187
rect -4817 -289 -4783 -255
rect -4817 -357 -4783 -323
rect -4817 -425 -4783 -391
rect -4817 -493 -4783 -459
rect -4817 -561 -4783 -527
rect -4817 -629 -4783 -595
rect -4817 -697 -4783 -663
rect -4817 -765 -4783 -731
rect -4817 -833 -4783 -799
rect -4817 -901 -4783 -867
rect -4817 -969 -4783 -935
rect -4721 935 -4687 969
rect -4721 867 -4687 901
rect -4721 799 -4687 833
rect -4721 731 -4687 765
rect -4721 663 -4687 697
rect -4721 595 -4687 629
rect -4721 527 -4687 561
rect -4721 459 -4687 493
rect -4721 391 -4687 425
rect -4721 323 -4687 357
rect -4721 255 -4687 289
rect -4721 187 -4687 221
rect -4721 119 -4687 153
rect -4721 51 -4687 85
rect -4721 -17 -4687 17
rect -4721 -85 -4687 -51
rect -4721 -153 -4687 -119
rect -4721 -221 -4687 -187
rect -4721 -289 -4687 -255
rect -4721 -357 -4687 -323
rect -4721 -425 -4687 -391
rect -4721 -493 -4687 -459
rect -4721 -561 -4687 -527
rect -4721 -629 -4687 -595
rect -4721 -697 -4687 -663
rect -4721 -765 -4687 -731
rect -4721 -833 -4687 -799
rect -4721 -901 -4687 -867
rect -4721 -969 -4687 -935
rect -4625 935 -4591 969
rect -4625 867 -4591 901
rect -4625 799 -4591 833
rect -4625 731 -4591 765
rect -4625 663 -4591 697
rect -4625 595 -4591 629
rect -4625 527 -4591 561
rect -4625 459 -4591 493
rect -4625 391 -4591 425
rect -4625 323 -4591 357
rect -4625 255 -4591 289
rect -4625 187 -4591 221
rect -4625 119 -4591 153
rect -4625 51 -4591 85
rect -4625 -17 -4591 17
rect -4625 -85 -4591 -51
rect -4625 -153 -4591 -119
rect -4625 -221 -4591 -187
rect -4625 -289 -4591 -255
rect -4625 -357 -4591 -323
rect -4625 -425 -4591 -391
rect -4625 -493 -4591 -459
rect -4625 -561 -4591 -527
rect -4625 -629 -4591 -595
rect -4625 -697 -4591 -663
rect -4625 -765 -4591 -731
rect -4625 -833 -4591 -799
rect -4625 -901 -4591 -867
rect -4625 -969 -4591 -935
rect -4529 935 -4495 969
rect -4529 867 -4495 901
rect -4529 799 -4495 833
rect -4529 731 -4495 765
rect -4529 663 -4495 697
rect -4529 595 -4495 629
rect -4529 527 -4495 561
rect -4529 459 -4495 493
rect -4529 391 -4495 425
rect -4529 323 -4495 357
rect -4529 255 -4495 289
rect -4529 187 -4495 221
rect -4529 119 -4495 153
rect -4529 51 -4495 85
rect -4529 -17 -4495 17
rect -4529 -85 -4495 -51
rect -4529 -153 -4495 -119
rect -4529 -221 -4495 -187
rect -4529 -289 -4495 -255
rect -4529 -357 -4495 -323
rect -4529 -425 -4495 -391
rect -4529 -493 -4495 -459
rect -4529 -561 -4495 -527
rect -4529 -629 -4495 -595
rect -4529 -697 -4495 -663
rect -4529 -765 -4495 -731
rect -4529 -833 -4495 -799
rect -4529 -901 -4495 -867
rect -4529 -969 -4495 -935
rect -4433 935 -4399 969
rect -4433 867 -4399 901
rect -4433 799 -4399 833
rect -4433 731 -4399 765
rect -4433 663 -4399 697
rect -4433 595 -4399 629
rect -4433 527 -4399 561
rect -4433 459 -4399 493
rect -4433 391 -4399 425
rect -4433 323 -4399 357
rect -4433 255 -4399 289
rect -4433 187 -4399 221
rect -4433 119 -4399 153
rect -4433 51 -4399 85
rect -4433 -17 -4399 17
rect -4433 -85 -4399 -51
rect -4433 -153 -4399 -119
rect -4433 -221 -4399 -187
rect -4433 -289 -4399 -255
rect -4433 -357 -4399 -323
rect -4433 -425 -4399 -391
rect -4433 -493 -4399 -459
rect -4433 -561 -4399 -527
rect -4433 -629 -4399 -595
rect -4433 -697 -4399 -663
rect -4433 -765 -4399 -731
rect -4433 -833 -4399 -799
rect -4433 -901 -4399 -867
rect -4433 -969 -4399 -935
rect -4337 935 -4303 969
rect -4337 867 -4303 901
rect -4337 799 -4303 833
rect -4337 731 -4303 765
rect -4337 663 -4303 697
rect -4337 595 -4303 629
rect -4337 527 -4303 561
rect -4337 459 -4303 493
rect -4337 391 -4303 425
rect -4337 323 -4303 357
rect -4337 255 -4303 289
rect -4337 187 -4303 221
rect -4337 119 -4303 153
rect -4337 51 -4303 85
rect -4337 -17 -4303 17
rect -4337 -85 -4303 -51
rect -4337 -153 -4303 -119
rect -4337 -221 -4303 -187
rect -4337 -289 -4303 -255
rect -4337 -357 -4303 -323
rect -4337 -425 -4303 -391
rect -4337 -493 -4303 -459
rect -4337 -561 -4303 -527
rect -4337 -629 -4303 -595
rect -4337 -697 -4303 -663
rect -4337 -765 -4303 -731
rect -4337 -833 -4303 -799
rect -4337 -901 -4303 -867
rect -4337 -969 -4303 -935
rect -4241 935 -4207 969
rect -4241 867 -4207 901
rect -4241 799 -4207 833
rect -4241 731 -4207 765
rect -4241 663 -4207 697
rect -4241 595 -4207 629
rect -4241 527 -4207 561
rect -4241 459 -4207 493
rect -4241 391 -4207 425
rect -4241 323 -4207 357
rect -4241 255 -4207 289
rect -4241 187 -4207 221
rect -4241 119 -4207 153
rect -4241 51 -4207 85
rect -4241 -17 -4207 17
rect -4241 -85 -4207 -51
rect -4241 -153 -4207 -119
rect -4241 -221 -4207 -187
rect -4241 -289 -4207 -255
rect -4241 -357 -4207 -323
rect -4241 -425 -4207 -391
rect -4241 -493 -4207 -459
rect -4241 -561 -4207 -527
rect -4241 -629 -4207 -595
rect -4241 -697 -4207 -663
rect -4241 -765 -4207 -731
rect -4241 -833 -4207 -799
rect -4241 -901 -4207 -867
rect -4241 -969 -4207 -935
rect -4145 935 -4111 969
rect -4145 867 -4111 901
rect -4145 799 -4111 833
rect -4145 731 -4111 765
rect -4145 663 -4111 697
rect -4145 595 -4111 629
rect -4145 527 -4111 561
rect -4145 459 -4111 493
rect -4145 391 -4111 425
rect -4145 323 -4111 357
rect -4145 255 -4111 289
rect -4145 187 -4111 221
rect -4145 119 -4111 153
rect -4145 51 -4111 85
rect -4145 -17 -4111 17
rect -4145 -85 -4111 -51
rect -4145 -153 -4111 -119
rect -4145 -221 -4111 -187
rect -4145 -289 -4111 -255
rect -4145 -357 -4111 -323
rect -4145 -425 -4111 -391
rect -4145 -493 -4111 -459
rect -4145 -561 -4111 -527
rect -4145 -629 -4111 -595
rect -4145 -697 -4111 -663
rect -4145 -765 -4111 -731
rect -4145 -833 -4111 -799
rect -4145 -901 -4111 -867
rect -4145 -969 -4111 -935
rect -4049 935 -4015 969
rect -4049 867 -4015 901
rect -4049 799 -4015 833
rect -4049 731 -4015 765
rect -4049 663 -4015 697
rect -4049 595 -4015 629
rect -4049 527 -4015 561
rect -4049 459 -4015 493
rect -4049 391 -4015 425
rect -4049 323 -4015 357
rect -4049 255 -4015 289
rect -4049 187 -4015 221
rect -4049 119 -4015 153
rect -4049 51 -4015 85
rect -4049 -17 -4015 17
rect -4049 -85 -4015 -51
rect -4049 -153 -4015 -119
rect -4049 -221 -4015 -187
rect -4049 -289 -4015 -255
rect -4049 -357 -4015 -323
rect -4049 -425 -4015 -391
rect -4049 -493 -4015 -459
rect -4049 -561 -4015 -527
rect -4049 -629 -4015 -595
rect -4049 -697 -4015 -663
rect -4049 -765 -4015 -731
rect -4049 -833 -4015 -799
rect -4049 -901 -4015 -867
rect -4049 -969 -4015 -935
rect -3953 935 -3919 969
rect -3953 867 -3919 901
rect -3953 799 -3919 833
rect -3953 731 -3919 765
rect -3953 663 -3919 697
rect -3953 595 -3919 629
rect -3953 527 -3919 561
rect -3953 459 -3919 493
rect -3953 391 -3919 425
rect -3953 323 -3919 357
rect -3953 255 -3919 289
rect -3953 187 -3919 221
rect -3953 119 -3919 153
rect -3953 51 -3919 85
rect -3953 -17 -3919 17
rect -3953 -85 -3919 -51
rect -3953 -153 -3919 -119
rect -3953 -221 -3919 -187
rect -3953 -289 -3919 -255
rect -3953 -357 -3919 -323
rect -3953 -425 -3919 -391
rect -3953 -493 -3919 -459
rect -3953 -561 -3919 -527
rect -3953 -629 -3919 -595
rect -3953 -697 -3919 -663
rect -3953 -765 -3919 -731
rect -3953 -833 -3919 -799
rect -3953 -901 -3919 -867
rect -3953 -969 -3919 -935
rect -3857 935 -3823 969
rect -3857 867 -3823 901
rect -3857 799 -3823 833
rect -3857 731 -3823 765
rect -3857 663 -3823 697
rect -3857 595 -3823 629
rect -3857 527 -3823 561
rect -3857 459 -3823 493
rect -3857 391 -3823 425
rect -3857 323 -3823 357
rect -3857 255 -3823 289
rect -3857 187 -3823 221
rect -3857 119 -3823 153
rect -3857 51 -3823 85
rect -3857 -17 -3823 17
rect -3857 -85 -3823 -51
rect -3857 -153 -3823 -119
rect -3857 -221 -3823 -187
rect -3857 -289 -3823 -255
rect -3857 -357 -3823 -323
rect -3857 -425 -3823 -391
rect -3857 -493 -3823 -459
rect -3857 -561 -3823 -527
rect -3857 -629 -3823 -595
rect -3857 -697 -3823 -663
rect -3857 -765 -3823 -731
rect -3857 -833 -3823 -799
rect -3857 -901 -3823 -867
rect -3857 -969 -3823 -935
rect -3761 935 -3727 969
rect -3761 867 -3727 901
rect -3761 799 -3727 833
rect -3761 731 -3727 765
rect -3761 663 -3727 697
rect -3761 595 -3727 629
rect -3761 527 -3727 561
rect -3761 459 -3727 493
rect -3761 391 -3727 425
rect -3761 323 -3727 357
rect -3761 255 -3727 289
rect -3761 187 -3727 221
rect -3761 119 -3727 153
rect -3761 51 -3727 85
rect -3761 -17 -3727 17
rect -3761 -85 -3727 -51
rect -3761 -153 -3727 -119
rect -3761 -221 -3727 -187
rect -3761 -289 -3727 -255
rect -3761 -357 -3727 -323
rect -3761 -425 -3727 -391
rect -3761 -493 -3727 -459
rect -3761 -561 -3727 -527
rect -3761 -629 -3727 -595
rect -3761 -697 -3727 -663
rect -3761 -765 -3727 -731
rect -3761 -833 -3727 -799
rect -3761 -901 -3727 -867
rect -3761 -969 -3727 -935
rect -3665 935 -3631 969
rect -3665 867 -3631 901
rect -3665 799 -3631 833
rect -3665 731 -3631 765
rect -3665 663 -3631 697
rect -3665 595 -3631 629
rect -3665 527 -3631 561
rect -3665 459 -3631 493
rect -3665 391 -3631 425
rect -3665 323 -3631 357
rect -3665 255 -3631 289
rect -3665 187 -3631 221
rect -3665 119 -3631 153
rect -3665 51 -3631 85
rect -3665 -17 -3631 17
rect -3665 -85 -3631 -51
rect -3665 -153 -3631 -119
rect -3665 -221 -3631 -187
rect -3665 -289 -3631 -255
rect -3665 -357 -3631 -323
rect -3665 -425 -3631 -391
rect -3665 -493 -3631 -459
rect -3665 -561 -3631 -527
rect -3665 -629 -3631 -595
rect -3665 -697 -3631 -663
rect -3665 -765 -3631 -731
rect -3665 -833 -3631 -799
rect -3665 -901 -3631 -867
rect -3665 -969 -3631 -935
rect -3569 935 -3535 969
rect -3569 867 -3535 901
rect -3569 799 -3535 833
rect -3569 731 -3535 765
rect -3569 663 -3535 697
rect -3569 595 -3535 629
rect -3569 527 -3535 561
rect -3569 459 -3535 493
rect -3569 391 -3535 425
rect -3569 323 -3535 357
rect -3569 255 -3535 289
rect -3569 187 -3535 221
rect -3569 119 -3535 153
rect -3569 51 -3535 85
rect -3569 -17 -3535 17
rect -3569 -85 -3535 -51
rect -3569 -153 -3535 -119
rect -3569 -221 -3535 -187
rect -3569 -289 -3535 -255
rect -3569 -357 -3535 -323
rect -3569 -425 -3535 -391
rect -3569 -493 -3535 -459
rect -3569 -561 -3535 -527
rect -3569 -629 -3535 -595
rect -3569 -697 -3535 -663
rect -3569 -765 -3535 -731
rect -3569 -833 -3535 -799
rect -3569 -901 -3535 -867
rect -3569 -969 -3535 -935
rect -3473 935 -3439 969
rect -3473 867 -3439 901
rect -3473 799 -3439 833
rect -3473 731 -3439 765
rect -3473 663 -3439 697
rect -3473 595 -3439 629
rect -3473 527 -3439 561
rect -3473 459 -3439 493
rect -3473 391 -3439 425
rect -3473 323 -3439 357
rect -3473 255 -3439 289
rect -3473 187 -3439 221
rect -3473 119 -3439 153
rect -3473 51 -3439 85
rect -3473 -17 -3439 17
rect -3473 -85 -3439 -51
rect -3473 -153 -3439 -119
rect -3473 -221 -3439 -187
rect -3473 -289 -3439 -255
rect -3473 -357 -3439 -323
rect -3473 -425 -3439 -391
rect -3473 -493 -3439 -459
rect -3473 -561 -3439 -527
rect -3473 -629 -3439 -595
rect -3473 -697 -3439 -663
rect -3473 -765 -3439 -731
rect -3473 -833 -3439 -799
rect -3473 -901 -3439 -867
rect -3473 -969 -3439 -935
rect -3377 935 -3343 969
rect -3377 867 -3343 901
rect -3377 799 -3343 833
rect -3377 731 -3343 765
rect -3377 663 -3343 697
rect -3377 595 -3343 629
rect -3377 527 -3343 561
rect -3377 459 -3343 493
rect -3377 391 -3343 425
rect -3377 323 -3343 357
rect -3377 255 -3343 289
rect -3377 187 -3343 221
rect -3377 119 -3343 153
rect -3377 51 -3343 85
rect -3377 -17 -3343 17
rect -3377 -85 -3343 -51
rect -3377 -153 -3343 -119
rect -3377 -221 -3343 -187
rect -3377 -289 -3343 -255
rect -3377 -357 -3343 -323
rect -3377 -425 -3343 -391
rect -3377 -493 -3343 -459
rect -3377 -561 -3343 -527
rect -3377 -629 -3343 -595
rect -3377 -697 -3343 -663
rect -3377 -765 -3343 -731
rect -3377 -833 -3343 -799
rect -3377 -901 -3343 -867
rect -3377 -969 -3343 -935
rect -3281 935 -3247 969
rect -3281 867 -3247 901
rect -3281 799 -3247 833
rect -3281 731 -3247 765
rect -3281 663 -3247 697
rect -3281 595 -3247 629
rect -3281 527 -3247 561
rect -3281 459 -3247 493
rect -3281 391 -3247 425
rect -3281 323 -3247 357
rect -3281 255 -3247 289
rect -3281 187 -3247 221
rect -3281 119 -3247 153
rect -3281 51 -3247 85
rect -3281 -17 -3247 17
rect -3281 -85 -3247 -51
rect -3281 -153 -3247 -119
rect -3281 -221 -3247 -187
rect -3281 -289 -3247 -255
rect -3281 -357 -3247 -323
rect -3281 -425 -3247 -391
rect -3281 -493 -3247 -459
rect -3281 -561 -3247 -527
rect -3281 -629 -3247 -595
rect -3281 -697 -3247 -663
rect -3281 -765 -3247 -731
rect -3281 -833 -3247 -799
rect -3281 -901 -3247 -867
rect -3281 -969 -3247 -935
rect -3185 935 -3151 969
rect -3185 867 -3151 901
rect -3185 799 -3151 833
rect -3185 731 -3151 765
rect -3185 663 -3151 697
rect -3185 595 -3151 629
rect -3185 527 -3151 561
rect -3185 459 -3151 493
rect -3185 391 -3151 425
rect -3185 323 -3151 357
rect -3185 255 -3151 289
rect -3185 187 -3151 221
rect -3185 119 -3151 153
rect -3185 51 -3151 85
rect -3185 -17 -3151 17
rect -3185 -85 -3151 -51
rect -3185 -153 -3151 -119
rect -3185 -221 -3151 -187
rect -3185 -289 -3151 -255
rect -3185 -357 -3151 -323
rect -3185 -425 -3151 -391
rect -3185 -493 -3151 -459
rect -3185 -561 -3151 -527
rect -3185 -629 -3151 -595
rect -3185 -697 -3151 -663
rect -3185 -765 -3151 -731
rect -3185 -833 -3151 -799
rect -3185 -901 -3151 -867
rect -3185 -969 -3151 -935
rect -3089 935 -3055 969
rect -3089 867 -3055 901
rect -3089 799 -3055 833
rect -3089 731 -3055 765
rect -3089 663 -3055 697
rect -3089 595 -3055 629
rect -3089 527 -3055 561
rect -3089 459 -3055 493
rect -3089 391 -3055 425
rect -3089 323 -3055 357
rect -3089 255 -3055 289
rect -3089 187 -3055 221
rect -3089 119 -3055 153
rect -3089 51 -3055 85
rect -3089 -17 -3055 17
rect -3089 -85 -3055 -51
rect -3089 -153 -3055 -119
rect -3089 -221 -3055 -187
rect -3089 -289 -3055 -255
rect -3089 -357 -3055 -323
rect -3089 -425 -3055 -391
rect -3089 -493 -3055 -459
rect -3089 -561 -3055 -527
rect -3089 -629 -3055 -595
rect -3089 -697 -3055 -663
rect -3089 -765 -3055 -731
rect -3089 -833 -3055 -799
rect -3089 -901 -3055 -867
rect -3089 -969 -3055 -935
rect -2993 935 -2959 969
rect -2993 867 -2959 901
rect -2993 799 -2959 833
rect -2993 731 -2959 765
rect -2993 663 -2959 697
rect -2993 595 -2959 629
rect -2993 527 -2959 561
rect -2993 459 -2959 493
rect -2993 391 -2959 425
rect -2993 323 -2959 357
rect -2993 255 -2959 289
rect -2993 187 -2959 221
rect -2993 119 -2959 153
rect -2993 51 -2959 85
rect -2993 -17 -2959 17
rect -2993 -85 -2959 -51
rect -2993 -153 -2959 -119
rect -2993 -221 -2959 -187
rect -2993 -289 -2959 -255
rect -2993 -357 -2959 -323
rect -2993 -425 -2959 -391
rect -2993 -493 -2959 -459
rect -2993 -561 -2959 -527
rect -2993 -629 -2959 -595
rect -2993 -697 -2959 -663
rect -2993 -765 -2959 -731
rect -2993 -833 -2959 -799
rect -2993 -901 -2959 -867
rect -2993 -969 -2959 -935
rect -2897 935 -2863 969
rect -2897 867 -2863 901
rect -2897 799 -2863 833
rect -2897 731 -2863 765
rect -2897 663 -2863 697
rect -2897 595 -2863 629
rect -2897 527 -2863 561
rect -2897 459 -2863 493
rect -2897 391 -2863 425
rect -2897 323 -2863 357
rect -2897 255 -2863 289
rect -2897 187 -2863 221
rect -2897 119 -2863 153
rect -2897 51 -2863 85
rect -2897 -17 -2863 17
rect -2897 -85 -2863 -51
rect -2897 -153 -2863 -119
rect -2897 -221 -2863 -187
rect -2897 -289 -2863 -255
rect -2897 -357 -2863 -323
rect -2897 -425 -2863 -391
rect -2897 -493 -2863 -459
rect -2897 -561 -2863 -527
rect -2897 -629 -2863 -595
rect -2897 -697 -2863 -663
rect -2897 -765 -2863 -731
rect -2897 -833 -2863 -799
rect -2897 -901 -2863 -867
rect -2897 -969 -2863 -935
rect -2801 935 -2767 969
rect -2801 867 -2767 901
rect -2801 799 -2767 833
rect -2801 731 -2767 765
rect -2801 663 -2767 697
rect -2801 595 -2767 629
rect -2801 527 -2767 561
rect -2801 459 -2767 493
rect -2801 391 -2767 425
rect -2801 323 -2767 357
rect -2801 255 -2767 289
rect -2801 187 -2767 221
rect -2801 119 -2767 153
rect -2801 51 -2767 85
rect -2801 -17 -2767 17
rect -2801 -85 -2767 -51
rect -2801 -153 -2767 -119
rect -2801 -221 -2767 -187
rect -2801 -289 -2767 -255
rect -2801 -357 -2767 -323
rect -2801 -425 -2767 -391
rect -2801 -493 -2767 -459
rect -2801 -561 -2767 -527
rect -2801 -629 -2767 -595
rect -2801 -697 -2767 -663
rect -2801 -765 -2767 -731
rect -2801 -833 -2767 -799
rect -2801 -901 -2767 -867
rect -2801 -969 -2767 -935
rect -2705 935 -2671 969
rect -2705 867 -2671 901
rect -2705 799 -2671 833
rect -2705 731 -2671 765
rect -2705 663 -2671 697
rect -2705 595 -2671 629
rect -2705 527 -2671 561
rect -2705 459 -2671 493
rect -2705 391 -2671 425
rect -2705 323 -2671 357
rect -2705 255 -2671 289
rect -2705 187 -2671 221
rect -2705 119 -2671 153
rect -2705 51 -2671 85
rect -2705 -17 -2671 17
rect -2705 -85 -2671 -51
rect -2705 -153 -2671 -119
rect -2705 -221 -2671 -187
rect -2705 -289 -2671 -255
rect -2705 -357 -2671 -323
rect -2705 -425 -2671 -391
rect -2705 -493 -2671 -459
rect -2705 -561 -2671 -527
rect -2705 -629 -2671 -595
rect -2705 -697 -2671 -663
rect -2705 -765 -2671 -731
rect -2705 -833 -2671 -799
rect -2705 -901 -2671 -867
rect -2705 -969 -2671 -935
rect -2609 935 -2575 969
rect -2609 867 -2575 901
rect -2609 799 -2575 833
rect -2609 731 -2575 765
rect -2609 663 -2575 697
rect -2609 595 -2575 629
rect -2609 527 -2575 561
rect -2609 459 -2575 493
rect -2609 391 -2575 425
rect -2609 323 -2575 357
rect -2609 255 -2575 289
rect -2609 187 -2575 221
rect -2609 119 -2575 153
rect -2609 51 -2575 85
rect -2609 -17 -2575 17
rect -2609 -85 -2575 -51
rect -2609 -153 -2575 -119
rect -2609 -221 -2575 -187
rect -2609 -289 -2575 -255
rect -2609 -357 -2575 -323
rect -2609 -425 -2575 -391
rect -2609 -493 -2575 -459
rect -2609 -561 -2575 -527
rect -2609 -629 -2575 -595
rect -2609 -697 -2575 -663
rect -2609 -765 -2575 -731
rect -2609 -833 -2575 -799
rect -2609 -901 -2575 -867
rect -2609 -969 -2575 -935
rect -2513 935 -2479 969
rect -2513 867 -2479 901
rect -2513 799 -2479 833
rect -2513 731 -2479 765
rect -2513 663 -2479 697
rect -2513 595 -2479 629
rect -2513 527 -2479 561
rect -2513 459 -2479 493
rect -2513 391 -2479 425
rect -2513 323 -2479 357
rect -2513 255 -2479 289
rect -2513 187 -2479 221
rect -2513 119 -2479 153
rect -2513 51 -2479 85
rect -2513 -17 -2479 17
rect -2513 -85 -2479 -51
rect -2513 -153 -2479 -119
rect -2513 -221 -2479 -187
rect -2513 -289 -2479 -255
rect -2513 -357 -2479 -323
rect -2513 -425 -2479 -391
rect -2513 -493 -2479 -459
rect -2513 -561 -2479 -527
rect -2513 -629 -2479 -595
rect -2513 -697 -2479 -663
rect -2513 -765 -2479 -731
rect -2513 -833 -2479 -799
rect -2513 -901 -2479 -867
rect -2513 -969 -2479 -935
rect -2417 935 -2383 969
rect -2417 867 -2383 901
rect -2417 799 -2383 833
rect -2417 731 -2383 765
rect -2417 663 -2383 697
rect -2417 595 -2383 629
rect -2417 527 -2383 561
rect -2417 459 -2383 493
rect -2417 391 -2383 425
rect -2417 323 -2383 357
rect -2417 255 -2383 289
rect -2417 187 -2383 221
rect -2417 119 -2383 153
rect -2417 51 -2383 85
rect -2417 -17 -2383 17
rect -2417 -85 -2383 -51
rect -2417 -153 -2383 -119
rect -2417 -221 -2383 -187
rect -2417 -289 -2383 -255
rect -2417 -357 -2383 -323
rect -2417 -425 -2383 -391
rect -2417 -493 -2383 -459
rect -2417 -561 -2383 -527
rect -2417 -629 -2383 -595
rect -2417 -697 -2383 -663
rect -2417 -765 -2383 -731
rect -2417 -833 -2383 -799
rect -2417 -901 -2383 -867
rect -2417 -969 -2383 -935
rect -2321 935 -2287 969
rect -2321 867 -2287 901
rect -2321 799 -2287 833
rect -2321 731 -2287 765
rect -2321 663 -2287 697
rect -2321 595 -2287 629
rect -2321 527 -2287 561
rect -2321 459 -2287 493
rect -2321 391 -2287 425
rect -2321 323 -2287 357
rect -2321 255 -2287 289
rect -2321 187 -2287 221
rect -2321 119 -2287 153
rect -2321 51 -2287 85
rect -2321 -17 -2287 17
rect -2321 -85 -2287 -51
rect -2321 -153 -2287 -119
rect -2321 -221 -2287 -187
rect -2321 -289 -2287 -255
rect -2321 -357 -2287 -323
rect -2321 -425 -2287 -391
rect -2321 -493 -2287 -459
rect -2321 -561 -2287 -527
rect -2321 -629 -2287 -595
rect -2321 -697 -2287 -663
rect -2321 -765 -2287 -731
rect -2321 -833 -2287 -799
rect -2321 -901 -2287 -867
rect -2321 -969 -2287 -935
rect -2225 935 -2191 969
rect -2225 867 -2191 901
rect -2225 799 -2191 833
rect -2225 731 -2191 765
rect -2225 663 -2191 697
rect -2225 595 -2191 629
rect -2225 527 -2191 561
rect -2225 459 -2191 493
rect -2225 391 -2191 425
rect -2225 323 -2191 357
rect -2225 255 -2191 289
rect -2225 187 -2191 221
rect -2225 119 -2191 153
rect -2225 51 -2191 85
rect -2225 -17 -2191 17
rect -2225 -85 -2191 -51
rect -2225 -153 -2191 -119
rect -2225 -221 -2191 -187
rect -2225 -289 -2191 -255
rect -2225 -357 -2191 -323
rect -2225 -425 -2191 -391
rect -2225 -493 -2191 -459
rect -2225 -561 -2191 -527
rect -2225 -629 -2191 -595
rect -2225 -697 -2191 -663
rect -2225 -765 -2191 -731
rect -2225 -833 -2191 -799
rect -2225 -901 -2191 -867
rect -2225 -969 -2191 -935
rect -2129 935 -2095 969
rect -2129 867 -2095 901
rect -2129 799 -2095 833
rect -2129 731 -2095 765
rect -2129 663 -2095 697
rect -2129 595 -2095 629
rect -2129 527 -2095 561
rect -2129 459 -2095 493
rect -2129 391 -2095 425
rect -2129 323 -2095 357
rect -2129 255 -2095 289
rect -2129 187 -2095 221
rect -2129 119 -2095 153
rect -2129 51 -2095 85
rect -2129 -17 -2095 17
rect -2129 -85 -2095 -51
rect -2129 -153 -2095 -119
rect -2129 -221 -2095 -187
rect -2129 -289 -2095 -255
rect -2129 -357 -2095 -323
rect -2129 -425 -2095 -391
rect -2129 -493 -2095 -459
rect -2129 -561 -2095 -527
rect -2129 -629 -2095 -595
rect -2129 -697 -2095 -663
rect -2129 -765 -2095 -731
rect -2129 -833 -2095 -799
rect -2129 -901 -2095 -867
rect -2129 -969 -2095 -935
rect -2033 935 -1999 969
rect -2033 867 -1999 901
rect -2033 799 -1999 833
rect -2033 731 -1999 765
rect -2033 663 -1999 697
rect -2033 595 -1999 629
rect -2033 527 -1999 561
rect -2033 459 -1999 493
rect -2033 391 -1999 425
rect -2033 323 -1999 357
rect -2033 255 -1999 289
rect -2033 187 -1999 221
rect -2033 119 -1999 153
rect -2033 51 -1999 85
rect -2033 -17 -1999 17
rect -2033 -85 -1999 -51
rect -2033 -153 -1999 -119
rect -2033 -221 -1999 -187
rect -2033 -289 -1999 -255
rect -2033 -357 -1999 -323
rect -2033 -425 -1999 -391
rect -2033 -493 -1999 -459
rect -2033 -561 -1999 -527
rect -2033 -629 -1999 -595
rect -2033 -697 -1999 -663
rect -2033 -765 -1999 -731
rect -2033 -833 -1999 -799
rect -2033 -901 -1999 -867
rect -2033 -969 -1999 -935
rect -1937 935 -1903 969
rect -1937 867 -1903 901
rect -1937 799 -1903 833
rect -1937 731 -1903 765
rect -1937 663 -1903 697
rect -1937 595 -1903 629
rect -1937 527 -1903 561
rect -1937 459 -1903 493
rect -1937 391 -1903 425
rect -1937 323 -1903 357
rect -1937 255 -1903 289
rect -1937 187 -1903 221
rect -1937 119 -1903 153
rect -1937 51 -1903 85
rect -1937 -17 -1903 17
rect -1937 -85 -1903 -51
rect -1937 -153 -1903 -119
rect -1937 -221 -1903 -187
rect -1937 -289 -1903 -255
rect -1937 -357 -1903 -323
rect -1937 -425 -1903 -391
rect -1937 -493 -1903 -459
rect -1937 -561 -1903 -527
rect -1937 -629 -1903 -595
rect -1937 -697 -1903 -663
rect -1937 -765 -1903 -731
rect -1937 -833 -1903 -799
rect -1937 -901 -1903 -867
rect -1937 -969 -1903 -935
rect -1841 935 -1807 969
rect -1841 867 -1807 901
rect -1841 799 -1807 833
rect -1841 731 -1807 765
rect -1841 663 -1807 697
rect -1841 595 -1807 629
rect -1841 527 -1807 561
rect -1841 459 -1807 493
rect -1841 391 -1807 425
rect -1841 323 -1807 357
rect -1841 255 -1807 289
rect -1841 187 -1807 221
rect -1841 119 -1807 153
rect -1841 51 -1807 85
rect -1841 -17 -1807 17
rect -1841 -85 -1807 -51
rect -1841 -153 -1807 -119
rect -1841 -221 -1807 -187
rect -1841 -289 -1807 -255
rect -1841 -357 -1807 -323
rect -1841 -425 -1807 -391
rect -1841 -493 -1807 -459
rect -1841 -561 -1807 -527
rect -1841 -629 -1807 -595
rect -1841 -697 -1807 -663
rect -1841 -765 -1807 -731
rect -1841 -833 -1807 -799
rect -1841 -901 -1807 -867
rect -1841 -969 -1807 -935
rect -1745 935 -1711 969
rect -1745 867 -1711 901
rect -1745 799 -1711 833
rect -1745 731 -1711 765
rect -1745 663 -1711 697
rect -1745 595 -1711 629
rect -1745 527 -1711 561
rect -1745 459 -1711 493
rect -1745 391 -1711 425
rect -1745 323 -1711 357
rect -1745 255 -1711 289
rect -1745 187 -1711 221
rect -1745 119 -1711 153
rect -1745 51 -1711 85
rect -1745 -17 -1711 17
rect -1745 -85 -1711 -51
rect -1745 -153 -1711 -119
rect -1745 -221 -1711 -187
rect -1745 -289 -1711 -255
rect -1745 -357 -1711 -323
rect -1745 -425 -1711 -391
rect -1745 -493 -1711 -459
rect -1745 -561 -1711 -527
rect -1745 -629 -1711 -595
rect -1745 -697 -1711 -663
rect -1745 -765 -1711 -731
rect -1745 -833 -1711 -799
rect -1745 -901 -1711 -867
rect -1745 -969 -1711 -935
rect -1649 935 -1615 969
rect -1649 867 -1615 901
rect -1649 799 -1615 833
rect -1649 731 -1615 765
rect -1649 663 -1615 697
rect -1649 595 -1615 629
rect -1649 527 -1615 561
rect -1649 459 -1615 493
rect -1649 391 -1615 425
rect -1649 323 -1615 357
rect -1649 255 -1615 289
rect -1649 187 -1615 221
rect -1649 119 -1615 153
rect -1649 51 -1615 85
rect -1649 -17 -1615 17
rect -1649 -85 -1615 -51
rect -1649 -153 -1615 -119
rect -1649 -221 -1615 -187
rect -1649 -289 -1615 -255
rect -1649 -357 -1615 -323
rect -1649 -425 -1615 -391
rect -1649 -493 -1615 -459
rect -1649 -561 -1615 -527
rect -1649 -629 -1615 -595
rect -1649 -697 -1615 -663
rect -1649 -765 -1615 -731
rect -1649 -833 -1615 -799
rect -1649 -901 -1615 -867
rect -1649 -969 -1615 -935
rect -1553 935 -1519 969
rect -1553 867 -1519 901
rect -1553 799 -1519 833
rect -1553 731 -1519 765
rect -1553 663 -1519 697
rect -1553 595 -1519 629
rect -1553 527 -1519 561
rect -1553 459 -1519 493
rect -1553 391 -1519 425
rect -1553 323 -1519 357
rect -1553 255 -1519 289
rect -1553 187 -1519 221
rect -1553 119 -1519 153
rect -1553 51 -1519 85
rect -1553 -17 -1519 17
rect -1553 -85 -1519 -51
rect -1553 -153 -1519 -119
rect -1553 -221 -1519 -187
rect -1553 -289 -1519 -255
rect -1553 -357 -1519 -323
rect -1553 -425 -1519 -391
rect -1553 -493 -1519 -459
rect -1553 -561 -1519 -527
rect -1553 -629 -1519 -595
rect -1553 -697 -1519 -663
rect -1553 -765 -1519 -731
rect -1553 -833 -1519 -799
rect -1553 -901 -1519 -867
rect -1553 -969 -1519 -935
rect -1457 935 -1423 969
rect -1457 867 -1423 901
rect -1457 799 -1423 833
rect -1457 731 -1423 765
rect -1457 663 -1423 697
rect -1457 595 -1423 629
rect -1457 527 -1423 561
rect -1457 459 -1423 493
rect -1457 391 -1423 425
rect -1457 323 -1423 357
rect -1457 255 -1423 289
rect -1457 187 -1423 221
rect -1457 119 -1423 153
rect -1457 51 -1423 85
rect -1457 -17 -1423 17
rect -1457 -85 -1423 -51
rect -1457 -153 -1423 -119
rect -1457 -221 -1423 -187
rect -1457 -289 -1423 -255
rect -1457 -357 -1423 -323
rect -1457 -425 -1423 -391
rect -1457 -493 -1423 -459
rect -1457 -561 -1423 -527
rect -1457 -629 -1423 -595
rect -1457 -697 -1423 -663
rect -1457 -765 -1423 -731
rect -1457 -833 -1423 -799
rect -1457 -901 -1423 -867
rect -1457 -969 -1423 -935
rect -1361 935 -1327 969
rect -1361 867 -1327 901
rect -1361 799 -1327 833
rect -1361 731 -1327 765
rect -1361 663 -1327 697
rect -1361 595 -1327 629
rect -1361 527 -1327 561
rect -1361 459 -1327 493
rect -1361 391 -1327 425
rect -1361 323 -1327 357
rect -1361 255 -1327 289
rect -1361 187 -1327 221
rect -1361 119 -1327 153
rect -1361 51 -1327 85
rect -1361 -17 -1327 17
rect -1361 -85 -1327 -51
rect -1361 -153 -1327 -119
rect -1361 -221 -1327 -187
rect -1361 -289 -1327 -255
rect -1361 -357 -1327 -323
rect -1361 -425 -1327 -391
rect -1361 -493 -1327 -459
rect -1361 -561 -1327 -527
rect -1361 -629 -1327 -595
rect -1361 -697 -1327 -663
rect -1361 -765 -1327 -731
rect -1361 -833 -1327 -799
rect -1361 -901 -1327 -867
rect -1361 -969 -1327 -935
rect -1265 935 -1231 969
rect -1265 867 -1231 901
rect -1265 799 -1231 833
rect -1265 731 -1231 765
rect -1265 663 -1231 697
rect -1265 595 -1231 629
rect -1265 527 -1231 561
rect -1265 459 -1231 493
rect -1265 391 -1231 425
rect -1265 323 -1231 357
rect -1265 255 -1231 289
rect -1265 187 -1231 221
rect -1265 119 -1231 153
rect -1265 51 -1231 85
rect -1265 -17 -1231 17
rect -1265 -85 -1231 -51
rect -1265 -153 -1231 -119
rect -1265 -221 -1231 -187
rect -1265 -289 -1231 -255
rect -1265 -357 -1231 -323
rect -1265 -425 -1231 -391
rect -1265 -493 -1231 -459
rect -1265 -561 -1231 -527
rect -1265 -629 -1231 -595
rect -1265 -697 -1231 -663
rect -1265 -765 -1231 -731
rect -1265 -833 -1231 -799
rect -1265 -901 -1231 -867
rect -1265 -969 -1231 -935
rect -1169 935 -1135 969
rect -1169 867 -1135 901
rect -1169 799 -1135 833
rect -1169 731 -1135 765
rect -1169 663 -1135 697
rect -1169 595 -1135 629
rect -1169 527 -1135 561
rect -1169 459 -1135 493
rect -1169 391 -1135 425
rect -1169 323 -1135 357
rect -1169 255 -1135 289
rect -1169 187 -1135 221
rect -1169 119 -1135 153
rect -1169 51 -1135 85
rect -1169 -17 -1135 17
rect -1169 -85 -1135 -51
rect -1169 -153 -1135 -119
rect -1169 -221 -1135 -187
rect -1169 -289 -1135 -255
rect -1169 -357 -1135 -323
rect -1169 -425 -1135 -391
rect -1169 -493 -1135 -459
rect -1169 -561 -1135 -527
rect -1169 -629 -1135 -595
rect -1169 -697 -1135 -663
rect -1169 -765 -1135 -731
rect -1169 -833 -1135 -799
rect -1169 -901 -1135 -867
rect -1169 -969 -1135 -935
rect -1073 935 -1039 969
rect -1073 867 -1039 901
rect -1073 799 -1039 833
rect -1073 731 -1039 765
rect -1073 663 -1039 697
rect -1073 595 -1039 629
rect -1073 527 -1039 561
rect -1073 459 -1039 493
rect -1073 391 -1039 425
rect -1073 323 -1039 357
rect -1073 255 -1039 289
rect -1073 187 -1039 221
rect -1073 119 -1039 153
rect -1073 51 -1039 85
rect -1073 -17 -1039 17
rect -1073 -85 -1039 -51
rect -1073 -153 -1039 -119
rect -1073 -221 -1039 -187
rect -1073 -289 -1039 -255
rect -1073 -357 -1039 -323
rect -1073 -425 -1039 -391
rect -1073 -493 -1039 -459
rect -1073 -561 -1039 -527
rect -1073 -629 -1039 -595
rect -1073 -697 -1039 -663
rect -1073 -765 -1039 -731
rect -1073 -833 -1039 -799
rect -1073 -901 -1039 -867
rect -1073 -969 -1039 -935
rect -977 935 -943 969
rect -977 867 -943 901
rect -977 799 -943 833
rect -977 731 -943 765
rect -977 663 -943 697
rect -977 595 -943 629
rect -977 527 -943 561
rect -977 459 -943 493
rect -977 391 -943 425
rect -977 323 -943 357
rect -977 255 -943 289
rect -977 187 -943 221
rect -977 119 -943 153
rect -977 51 -943 85
rect -977 -17 -943 17
rect -977 -85 -943 -51
rect -977 -153 -943 -119
rect -977 -221 -943 -187
rect -977 -289 -943 -255
rect -977 -357 -943 -323
rect -977 -425 -943 -391
rect -977 -493 -943 -459
rect -977 -561 -943 -527
rect -977 -629 -943 -595
rect -977 -697 -943 -663
rect -977 -765 -943 -731
rect -977 -833 -943 -799
rect -977 -901 -943 -867
rect -977 -969 -943 -935
rect -881 935 -847 969
rect -881 867 -847 901
rect -881 799 -847 833
rect -881 731 -847 765
rect -881 663 -847 697
rect -881 595 -847 629
rect -881 527 -847 561
rect -881 459 -847 493
rect -881 391 -847 425
rect -881 323 -847 357
rect -881 255 -847 289
rect -881 187 -847 221
rect -881 119 -847 153
rect -881 51 -847 85
rect -881 -17 -847 17
rect -881 -85 -847 -51
rect -881 -153 -847 -119
rect -881 -221 -847 -187
rect -881 -289 -847 -255
rect -881 -357 -847 -323
rect -881 -425 -847 -391
rect -881 -493 -847 -459
rect -881 -561 -847 -527
rect -881 -629 -847 -595
rect -881 -697 -847 -663
rect -881 -765 -847 -731
rect -881 -833 -847 -799
rect -881 -901 -847 -867
rect -881 -969 -847 -935
rect -785 935 -751 969
rect -785 867 -751 901
rect -785 799 -751 833
rect -785 731 -751 765
rect -785 663 -751 697
rect -785 595 -751 629
rect -785 527 -751 561
rect -785 459 -751 493
rect -785 391 -751 425
rect -785 323 -751 357
rect -785 255 -751 289
rect -785 187 -751 221
rect -785 119 -751 153
rect -785 51 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -51
rect -785 -153 -751 -119
rect -785 -221 -751 -187
rect -785 -289 -751 -255
rect -785 -357 -751 -323
rect -785 -425 -751 -391
rect -785 -493 -751 -459
rect -785 -561 -751 -527
rect -785 -629 -751 -595
rect -785 -697 -751 -663
rect -785 -765 -751 -731
rect -785 -833 -751 -799
rect -785 -901 -751 -867
rect -785 -969 -751 -935
rect -689 935 -655 969
rect -689 867 -655 901
rect -689 799 -655 833
rect -689 731 -655 765
rect -689 663 -655 697
rect -689 595 -655 629
rect -689 527 -655 561
rect -689 459 -655 493
rect -689 391 -655 425
rect -689 323 -655 357
rect -689 255 -655 289
rect -689 187 -655 221
rect -689 119 -655 153
rect -689 51 -655 85
rect -689 -17 -655 17
rect -689 -85 -655 -51
rect -689 -153 -655 -119
rect -689 -221 -655 -187
rect -689 -289 -655 -255
rect -689 -357 -655 -323
rect -689 -425 -655 -391
rect -689 -493 -655 -459
rect -689 -561 -655 -527
rect -689 -629 -655 -595
rect -689 -697 -655 -663
rect -689 -765 -655 -731
rect -689 -833 -655 -799
rect -689 -901 -655 -867
rect -689 -969 -655 -935
rect -593 935 -559 969
rect -593 867 -559 901
rect -593 799 -559 833
rect -593 731 -559 765
rect -593 663 -559 697
rect -593 595 -559 629
rect -593 527 -559 561
rect -593 459 -559 493
rect -593 391 -559 425
rect -593 323 -559 357
rect -593 255 -559 289
rect -593 187 -559 221
rect -593 119 -559 153
rect -593 51 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -51
rect -593 -153 -559 -119
rect -593 -221 -559 -187
rect -593 -289 -559 -255
rect -593 -357 -559 -323
rect -593 -425 -559 -391
rect -593 -493 -559 -459
rect -593 -561 -559 -527
rect -593 -629 -559 -595
rect -593 -697 -559 -663
rect -593 -765 -559 -731
rect -593 -833 -559 -799
rect -593 -901 -559 -867
rect -593 -969 -559 -935
rect -497 935 -463 969
rect -497 867 -463 901
rect -497 799 -463 833
rect -497 731 -463 765
rect -497 663 -463 697
rect -497 595 -463 629
rect -497 527 -463 561
rect -497 459 -463 493
rect -497 391 -463 425
rect -497 323 -463 357
rect -497 255 -463 289
rect -497 187 -463 221
rect -497 119 -463 153
rect -497 51 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -51
rect -497 -153 -463 -119
rect -497 -221 -463 -187
rect -497 -289 -463 -255
rect -497 -357 -463 -323
rect -497 -425 -463 -391
rect -497 -493 -463 -459
rect -497 -561 -463 -527
rect -497 -629 -463 -595
rect -497 -697 -463 -663
rect -497 -765 -463 -731
rect -497 -833 -463 -799
rect -497 -901 -463 -867
rect -497 -969 -463 -935
rect -401 935 -367 969
rect -401 867 -367 901
rect -401 799 -367 833
rect -401 731 -367 765
rect -401 663 -367 697
rect -401 595 -367 629
rect -401 527 -367 561
rect -401 459 -367 493
rect -401 391 -367 425
rect -401 323 -367 357
rect -401 255 -367 289
rect -401 187 -367 221
rect -401 119 -367 153
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -401 -153 -367 -119
rect -401 -221 -367 -187
rect -401 -289 -367 -255
rect -401 -357 -367 -323
rect -401 -425 -367 -391
rect -401 -493 -367 -459
rect -401 -561 -367 -527
rect -401 -629 -367 -595
rect -401 -697 -367 -663
rect -401 -765 -367 -731
rect -401 -833 -367 -799
rect -401 -901 -367 -867
rect -401 -969 -367 -935
rect -305 935 -271 969
rect -305 867 -271 901
rect -305 799 -271 833
rect -305 731 -271 765
rect -305 663 -271 697
rect -305 595 -271 629
rect -305 527 -271 561
rect -305 459 -271 493
rect -305 391 -271 425
rect -305 323 -271 357
rect -305 255 -271 289
rect -305 187 -271 221
rect -305 119 -271 153
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -305 -153 -271 -119
rect -305 -221 -271 -187
rect -305 -289 -271 -255
rect -305 -357 -271 -323
rect -305 -425 -271 -391
rect -305 -493 -271 -459
rect -305 -561 -271 -527
rect -305 -629 -271 -595
rect -305 -697 -271 -663
rect -305 -765 -271 -731
rect -305 -833 -271 -799
rect -305 -901 -271 -867
rect -305 -969 -271 -935
rect -209 935 -175 969
rect -209 867 -175 901
rect -209 799 -175 833
rect -209 731 -175 765
rect -209 663 -175 697
rect -209 595 -175 629
rect -209 527 -175 561
rect -209 459 -175 493
rect -209 391 -175 425
rect -209 323 -175 357
rect -209 255 -175 289
rect -209 187 -175 221
rect -209 119 -175 153
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -209 -153 -175 -119
rect -209 -221 -175 -187
rect -209 -289 -175 -255
rect -209 -357 -175 -323
rect -209 -425 -175 -391
rect -209 -493 -175 -459
rect -209 -561 -175 -527
rect -209 -629 -175 -595
rect -209 -697 -175 -663
rect -209 -765 -175 -731
rect -209 -833 -175 -799
rect -209 -901 -175 -867
rect -209 -969 -175 -935
rect -113 935 -79 969
rect -113 867 -79 901
rect -113 799 -79 833
rect -113 731 -79 765
rect -113 663 -79 697
rect -113 595 -79 629
rect -113 527 -79 561
rect -113 459 -79 493
rect -113 391 -79 425
rect -113 323 -79 357
rect -113 255 -79 289
rect -113 187 -79 221
rect -113 119 -79 153
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -113 -153 -79 -119
rect -113 -221 -79 -187
rect -113 -289 -79 -255
rect -113 -357 -79 -323
rect -113 -425 -79 -391
rect -113 -493 -79 -459
rect -113 -561 -79 -527
rect -113 -629 -79 -595
rect -113 -697 -79 -663
rect -113 -765 -79 -731
rect -113 -833 -79 -799
rect -113 -901 -79 -867
rect -113 -969 -79 -935
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect 79 935 113 969
rect 79 867 113 901
rect 79 799 113 833
rect 79 731 113 765
rect 79 663 113 697
rect 79 595 113 629
rect 79 527 113 561
rect 79 459 113 493
rect 79 391 113 425
rect 79 323 113 357
rect 79 255 113 289
rect 79 187 113 221
rect 79 119 113 153
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 79 -153 113 -119
rect 79 -221 113 -187
rect 79 -289 113 -255
rect 79 -357 113 -323
rect 79 -425 113 -391
rect 79 -493 113 -459
rect 79 -561 113 -527
rect 79 -629 113 -595
rect 79 -697 113 -663
rect 79 -765 113 -731
rect 79 -833 113 -799
rect 79 -901 113 -867
rect 79 -969 113 -935
rect 175 935 209 969
rect 175 867 209 901
rect 175 799 209 833
rect 175 731 209 765
rect 175 663 209 697
rect 175 595 209 629
rect 175 527 209 561
rect 175 459 209 493
rect 175 391 209 425
rect 175 323 209 357
rect 175 255 209 289
rect 175 187 209 221
rect 175 119 209 153
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 175 -153 209 -119
rect 175 -221 209 -187
rect 175 -289 209 -255
rect 175 -357 209 -323
rect 175 -425 209 -391
rect 175 -493 209 -459
rect 175 -561 209 -527
rect 175 -629 209 -595
rect 175 -697 209 -663
rect 175 -765 209 -731
rect 175 -833 209 -799
rect 175 -901 209 -867
rect 175 -969 209 -935
rect 271 935 305 969
rect 271 867 305 901
rect 271 799 305 833
rect 271 731 305 765
rect 271 663 305 697
rect 271 595 305 629
rect 271 527 305 561
rect 271 459 305 493
rect 271 391 305 425
rect 271 323 305 357
rect 271 255 305 289
rect 271 187 305 221
rect 271 119 305 153
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
rect 271 -153 305 -119
rect 271 -221 305 -187
rect 271 -289 305 -255
rect 271 -357 305 -323
rect 271 -425 305 -391
rect 271 -493 305 -459
rect 271 -561 305 -527
rect 271 -629 305 -595
rect 271 -697 305 -663
rect 271 -765 305 -731
rect 271 -833 305 -799
rect 271 -901 305 -867
rect 271 -969 305 -935
rect 367 935 401 969
rect 367 867 401 901
rect 367 799 401 833
rect 367 731 401 765
rect 367 663 401 697
rect 367 595 401 629
rect 367 527 401 561
rect 367 459 401 493
rect 367 391 401 425
rect 367 323 401 357
rect 367 255 401 289
rect 367 187 401 221
rect 367 119 401 153
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 367 -153 401 -119
rect 367 -221 401 -187
rect 367 -289 401 -255
rect 367 -357 401 -323
rect 367 -425 401 -391
rect 367 -493 401 -459
rect 367 -561 401 -527
rect 367 -629 401 -595
rect 367 -697 401 -663
rect 367 -765 401 -731
rect 367 -833 401 -799
rect 367 -901 401 -867
rect 367 -969 401 -935
rect 463 935 497 969
rect 463 867 497 901
rect 463 799 497 833
rect 463 731 497 765
rect 463 663 497 697
rect 463 595 497 629
rect 463 527 497 561
rect 463 459 497 493
rect 463 391 497 425
rect 463 323 497 357
rect 463 255 497 289
rect 463 187 497 221
rect 463 119 497 153
rect 463 51 497 85
rect 463 -17 497 17
rect 463 -85 497 -51
rect 463 -153 497 -119
rect 463 -221 497 -187
rect 463 -289 497 -255
rect 463 -357 497 -323
rect 463 -425 497 -391
rect 463 -493 497 -459
rect 463 -561 497 -527
rect 463 -629 497 -595
rect 463 -697 497 -663
rect 463 -765 497 -731
rect 463 -833 497 -799
rect 463 -901 497 -867
rect 463 -969 497 -935
rect 559 935 593 969
rect 559 867 593 901
rect 559 799 593 833
rect 559 731 593 765
rect 559 663 593 697
rect 559 595 593 629
rect 559 527 593 561
rect 559 459 593 493
rect 559 391 593 425
rect 559 323 593 357
rect 559 255 593 289
rect 559 187 593 221
rect 559 119 593 153
rect 559 51 593 85
rect 559 -17 593 17
rect 559 -85 593 -51
rect 559 -153 593 -119
rect 559 -221 593 -187
rect 559 -289 593 -255
rect 559 -357 593 -323
rect 559 -425 593 -391
rect 559 -493 593 -459
rect 559 -561 593 -527
rect 559 -629 593 -595
rect 559 -697 593 -663
rect 559 -765 593 -731
rect 559 -833 593 -799
rect 559 -901 593 -867
rect 559 -969 593 -935
rect 655 935 689 969
rect 655 867 689 901
rect 655 799 689 833
rect 655 731 689 765
rect 655 663 689 697
rect 655 595 689 629
rect 655 527 689 561
rect 655 459 689 493
rect 655 391 689 425
rect 655 323 689 357
rect 655 255 689 289
rect 655 187 689 221
rect 655 119 689 153
rect 655 51 689 85
rect 655 -17 689 17
rect 655 -85 689 -51
rect 655 -153 689 -119
rect 655 -221 689 -187
rect 655 -289 689 -255
rect 655 -357 689 -323
rect 655 -425 689 -391
rect 655 -493 689 -459
rect 655 -561 689 -527
rect 655 -629 689 -595
rect 655 -697 689 -663
rect 655 -765 689 -731
rect 655 -833 689 -799
rect 655 -901 689 -867
rect 655 -969 689 -935
rect 751 935 785 969
rect 751 867 785 901
rect 751 799 785 833
rect 751 731 785 765
rect 751 663 785 697
rect 751 595 785 629
rect 751 527 785 561
rect 751 459 785 493
rect 751 391 785 425
rect 751 323 785 357
rect 751 255 785 289
rect 751 187 785 221
rect 751 119 785 153
rect 751 51 785 85
rect 751 -17 785 17
rect 751 -85 785 -51
rect 751 -153 785 -119
rect 751 -221 785 -187
rect 751 -289 785 -255
rect 751 -357 785 -323
rect 751 -425 785 -391
rect 751 -493 785 -459
rect 751 -561 785 -527
rect 751 -629 785 -595
rect 751 -697 785 -663
rect 751 -765 785 -731
rect 751 -833 785 -799
rect 751 -901 785 -867
rect 751 -969 785 -935
rect 847 935 881 969
rect 847 867 881 901
rect 847 799 881 833
rect 847 731 881 765
rect 847 663 881 697
rect 847 595 881 629
rect 847 527 881 561
rect 847 459 881 493
rect 847 391 881 425
rect 847 323 881 357
rect 847 255 881 289
rect 847 187 881 221
rect 847 119 881 153
rect 847 51 881 85
rect 847 -17 881 17
rect 847 -85 881 -51
rect 847 -153 881 -119
rect 847 -221 881 -187
rect 847 -289 881 -255
rect 847 -357 881 -323
rect 847 -425 881 -391
rect 847 -493 881 -459
rect 847 -561 881 -527
rect 847 -629 881 -595
rect 847 -697 881 -663
rect 847 -765 881 -731
rect 847 -833 881 -799
rect 847 -901 881 -867
rect 847 -969 881 -935
rect 943 935 977 969
rect 943 867 977 901
rect 943 799 977 833
rect 943 731 977 765
rect 943 663 977 697
rect 943 595 977 629
rect 943 527 977 561
rect 943 459 977 493
rect 943 391 977 425
rect 943 323 977 357
rect 943 255 977 289
rect 943 187 977 221
rect 943 119 977 153
rect 943 51 977 85
rect 943 -17 977 17
rect 943 -85 977 -51
rect 943 -153 977 -119
rect 943 -221 977 -187
rect 943 -289 977 -255
rect 943 -357 977 -323
rect 943 -425 977 -391
rect 943 -493 977 -459
rect 943 -561 977 -527
rect 943 -629 977 -595
rect 943 -697 977 -663
rect 943 -765 977 -731
rect 943 -833 977 -799
rect 943 -901 977 -867
rect 943 -969 977 -935
rect 1039 935 1073 969
rect 1039 867 1073 901
rect 1039 799 1073 833
rect 1039 731 1073 765
rect 1039 663 1073 697
rect 1039 595 1073 629
rect 1039 527 1073 561
rect 1039 459 1073 493
rect 1039 391 1073 425
rect 1039 323 1073 357
rect 1039 255 1073 289
rect 1039 187 1073 221
rect 1039 119 1073 153
rect 1039 51 1073 85
rect 1039 -17 1073 17
rect 1039 -85 1073 -51
rect 1039 -153 1073 -119
rect 1039 -221 1073 -187
rect 1039 -289 1073 -255
rect 1039 -357 1073 -323
rect 1039 -425 1073 -391
rect 1039 -493 1073 -459
rect 1039 -561 1073 -527
rect 1039 -629 1073 -595
rect 1039 -697 1073 -663
rect 1039 -765 1073 -731
rect 1039 -833 1073 -799
rect 1039 -901 1073 -867
rect 1039 -969 1073 -935
rect 1135 935 1169 969
rect 1135 867 1169 901
rect 1135 799 1169 833
rect 1135 731 1169 765
rect 1135 663 1169 697
rect 1135 595 1169 629
rect 1135 527 1169 561
rect 1135 459 1169 493
rect 1135 391 1169 425
rect 1135 323 1169 357
rect 1135 255 1169 289
rect 1135 187 1169 221
rect 1135 119 1169 153
rect 1135 51 1169 85
rect 1135 -17 1169 17
rect 1135 -85 1169 -51
rect 1135 -153 1169 -119
rect 1135 -221 1169 -187
rect 1135 -289 1169 -255
rect 1135 -357 1169 -323
rect 1135 -425 1169 -391
rect 1135 -493 1169 -459
rect 1135 -561 1169 -527
rect 1135 -629 1169 -595
rect 1135 -697 1169 -663
rect 1135 -765 1169 -731
rect 1135 -833 1169 -799
rect 1135 -901 1169 -867
rect 1135 -969 1169 -935
rect 1231 935 1265 969
rect 1231 867 1265 901
rect 1231 799 1265 833
rect 1231 731 1265 765
rect 1231 663 1265 697
rect 1231 595 1265 629
rect 1231 527 1265 561
rect 1231 459 1265 493
rect 1231 391 1265 425
rect 1231 323 1265 357
rect 1231 255 1265 289
rect 1231 187 1265 221
rect 1231 119 1265 153
rect 1231 51 1265 85
rect 1231 -17 1265 17
rect 1231 -85 1265 -51
rect 1231 -153 1265 -119
rect 1231 -221 1265 -187
rect 1231 -289 1265 -255
rect 1231 -357 1265 -323
rect 1231 -425 1265 -391
rect 1231 -493 1265 -459
rect 1231 -561 1265 -527
rect 1231 -629 1265 -595
rect 1231 -697 1265 -663
rect 1231 -765 1265 -731
rect 1231 -833 1265 -799
rect 1231 -901 1265 -867
rect 1231 -969 1265 -935
rect 1327 935 1361 969
rect 1327 867 1361 901
rect 1327 799 1361 833
rect 1327 731 1361 765
rect 1327 663 1361 697
rect 1327 595 1361 629
rect 1327 527 1361 561
rect 1327 459 1361 493
rect 1327 391 1361 425
rect 1327 323 1361 357
rect 1327 255 1361 289
rect 1327 187 1361 221
rect 1327 119 1361 153
rect 1327 51 1361 85
rect 1327 -17 1361 17
rect 1327 -85 1361 -51
rect 1327 -153 1361 -119
rect 1327 -221 1361 -187
rect 1327 -289 1361 -255
rect 1327 -357 1361 -323
rect 1327 -425 1361 -391
rect 1327 -493 1361 -459
rect 1327 -561 1361 -527
rect 1327 -629 1361 -595
rect 1327 -697 1361 -663
rect 1327 -765 1361 -731
rect 1327 -833 1361 -799
rect 1327 -901 1361 -867
rect 1327 -969 1361 -935
rect 1423 935 1457 969
rect 1423 867 1457 901
rect 1423 799 1457 833
rect 1423 731 1457 765
rect 1423 663 1457 697
rect 1423 595 1457 629
rect 1423 527 1457 561
rect 1423 459 1457 493
rect 1423 391 1457 425
rect 1423 323 1457 357
rect 1423 255 1457 289
rect 1423 187 1457 221
rect 1423 119 1457 153
rect 1423 51 1457 85
rect 1423 -17 1457 17
rect 1423 -85 1457 -51
rect 1423 -153 1457 -119
rect 1423 -221 1457 -187
rect 1423 -289 1457 -255
rect 1423 -357 1457 -323
rect 1423 -425 1457 -391
rect 1423 -493 1457 -459
rect 1423 -561 1457 -527
rect 1423 -629 1457 -595
rect 1423 -697 1457 -663
rect 1423 -765 1457 -731
rect 1423 -833 1457 -799
rect 1423 -901 1457 -867
rect 1423 -969 1457 -935
rect 1519 935 1553 969
rect 1519 867 1553 901
rect 1519 799 1553 833
rect 1519 731 1553 765
rect 1519 663 1553 697
rect 1519 595 1553 629
rect 1519 527 1553 561
rect 1519 459 1553 493
rect 1519 391 1553 425
rect 1519 323 1553 357
rect 1519 255 1553 289
rect 1519 187 1553 221
rect 1519 119 1553 153
rect 1519 51 1553 85
rect 1519 -17 1553 17
rect 1519 -85 1553 -51
rect 1519 -153 1553 -119
rect 1519 -221 1553 -187
rect 1519 -289 1553 -255
rect 1519 -357 1553 -323
rect 1519 -425 1553 -391
rect 1519 -493 1553 -459
rect 1519 -561 1553 -527
rect 1519 -629 1553 -595
rect 1519 -697 1553 -663
rect 1519 -765 1553 -731
rect 1519 -833 1553 -799
rect 1519 -901 1553 -867
rect 1519 -969 1553 -935
rect 1615 935 1649 969
rect 1615 867 1649 901
rect 1615 799 1649 833
rect 1615 731 1649 765
rect 1615 663 1649 697
rect 1615 595 1649 629
rect 1615 527 1649 561
rect 1615 459 1649 493
rect 1615 391 1649 425
rect 1615 323 1649 357
rect 1615 255 1649 289
rect 1615 187 1649 221
rect 1615 119 1649 153
rect 1615 51 1649 85
rect 1615 -17 1649 17
rect 1615 -85 1649 -51
rect 1615 -153 1649 -119
rect 1615 -221 1649 -187
rect 1615 -289 1649 -255
rect 1615 -357 1649 -323
rect 1615 -425 1649 -391
rect 1615 -493 1649 -459
rect 1615 -561 1649 -527
rect 1615 -629 1649 -595
rect 1615 -697 1649 -663
rect 1615 -765 1649 -731
rect 1615 -833 1649 -799
rect 1615 -901 1649 -867
rect 1615 -969 1649 -935
rect 1711 935 1745 969
rect 1711 867 1745 901
rect 1711 799 1745 833
rect 1711 731 1745 765
rect 1711 663 1745 697
rect 1711 595 1745 629
rect 1711 527 1745 561
rect 1711 459 1745 493
rect 1711 391 1745 425
rect 1711 323 1745 357
rect 1711 255 1745 289
rect 1711 187 1745 221
rect 1711 119 1745 153
rect 1711 51 1745 85
rect 1711 -17 1745 17
rect 1711 -85 1745 -51
rect 1711 -153 1745 -119
rect 1711 -221 1745 -187
rect 1711 -289 1745 -255
rect 1711 -357 1745 -323
rect 1711 -425 1745 -391
rect 1711 -493 1745 -459
rect 1711 -561 1745 -527
rect 1711 -629 1745 -595
rect 1711 -697 1745 -663
rect 1711 -765 1745 -731
rect 1711 -833 1745 -799
rect 1711 -901 1745 -867
rect 1711 -969 1745 -935
rect 1807 935 1841 969
rect 1807 867 1841 901
rect 1807 799 1841 833
rect 1807 731 1841 765
rect 1807 663 1841 697
rect 1807 595 1841 629
rect 1807 527 1841 561
rect 1807 459 1841 493
rect 1807 391 1841 425
rect 1807 323 1841 357
rect 1807 255 1841 289
rect 1807 187 1841 221
rect 1807 119 1841 153
rect 1807 51 1841 85
rect 1807 -17 1841 17
rect 1807 -85 1841 -51
rect 1807 -153 1841 -119
rect 1807 -221 1841 -187
rect 1807 -289 1841 -255
rect 1807 -357 1841 -323
rect 1807 -425 1841 -391
rect 1807 -493 1841 -459
rect 1807 -561 1841 -527
rect 1807 -629 1841 -595
rect 1807 -697 1841 -663
rect 1807 -765 1841 -731
rect 1807 -833 1841 -799
rect 1807 -901 1841 -867
rect 1807 -969 1841 -935
rect 1903 935 1937 969
rect 1903 867 1937 901
rect 1903 799 1937 833
rect 1903 731 1937 765
rect 1903 663 1937 697
rect 1903 595 1937 629
rect 1903 527 1937 561
rect 1903 459 1937 493
rect 1903 391 1937 425
rect 1903 323 1937 357
rect 1903 255 1937 289
rect 1903 187 1937 221
rect 1903 119 1937 153
rect 1903 51 1937 85
rect 1903 -17 1937 17
rect 1903 -85 1937 -51
rect 1903 -153 1937 -119
rect 1903 -221 1937 -187
rect 1903 -289 1937 -255
rect 1903 -357 1937 -323
rect 1903 -425 1937 -391
rect 1903 -493 1937 -459
rect 1903 -561 1937 -527
rect 1903 -629 1937 -595
rect 1903 -697 1937 -663
rect 1903 -765 1937 -731
rect 1903 -833 1937 -799
rect 1903 -901 1937 -867
rect 1903 -969 1937 -935
rect 1999 935 2033 969
rect 1999 867 2033 901
rect 1999 799 2033 833
rect 1999 731 2033 765
rect 1999 663 2033 697
rect 1999 595 2033 629
rect 1999 527 2033 561
rect 1999 459 2033 493
rect 1999 391 2033 425
rect 1999 323 2033 357
rect 1999 255 2033 289
rect 1999 187 2033 221
rect 1999 119 2033 153
rect 1999 51 2033 85
rect 1999 -17 2033 17
rect 1999 -85 2033 -51
rect 1999 -153 2033 -119
rect 1999 -221 2033 -187
rect 1999 -289 2033 -255
rect 1999 -357 2033 -323
rect 1999 -425 2033 -391
rect 1999 -493 2033 -459
rect 1999 -561 2033 -527
rect 1999 -629 2033 -595
rect 1999 -697 2033 -663
rect 1999 -765 2033 -731
rect 1999 -833 2033 -799
rect 1999 -901 2033 -867
rect 1999 -969 2033 -935
rect 2095 935 2129 969
rect 2095 867 2129 901
rect 2095 799 2129 833
rect 2095 731 2129 765
rect 2095 663 2129 697
rect 2095 595 2129 629
rect 2095 527 2129 561
rect 2095 459 2129 493
rect 2095 391 2129 425
rect 2095 323 2129 357
rect 2095 255 2129 289
rect 2095 187 2129 221
rect 2095 119 2129 153
rect 2095 51 2129 85
rect 2095 -17 2129 17
rect 2095 -85 2129 -51
rect 2095 -153 2129 -119
rect 2095 -221 2129 -187
rect 2095 -289 2129 -255
rect 2095 -357 2129 -323
rect 2095 -425 2129 -391
rect 2095 -493 2129 -459
rect 2095 -561 2129 -527
rect 2095 -629 2129 -595
rect 2095 -697 2129 -663
rect 2095 -765 2129 -731
rect 2095 -833 2129 -799
rect 2095 -901 2129 -867
rect 2095 -969 2129 -935
rect 2191 935 2225 969
rect 2191 867 2225 901
rect 2191 799 2225 833
rect 2191 731 2225 765
rect 2191 663 2225 697
rect 2191 595 2225 629
rect 2191 527 2225 561
rect 2191 459 2225 493
rect 2191 391 2225 425
rect 2191 323 2225 357
rect 2191 255 2225 289
rect 2191 187 2225 221
rect 2191 119 2225 153
rect 2191 51 2225 85
rect 2191 -17 2225 17
rect 2191 -85 2225 -51
rect 2191 -153 2225 -119
rect 2191 -221 2225 -187
rect 2191 -289 2225 -255
rect 2191 -357 2225 -323
rect 2191 -425 2225 -391
rect 2191 -493 2225 -459
rect 2191 -561 2225 -527
rect 2191 -629 2225 -595
rect 2191 -697 2225 -663
rect 2191 -765 2225 -731
rect 2191 -833 2225 -799
rect 2191 -901 2225 -867
rect 2191 -969 2225 -935
rect 2287 935 2321 969
rect 2287 867 2321 901
rect 2287 799 2321 833
rect 2287 731 2321 765
rect 2287 663 2321 697
rect 2287 595 2321 629
rect 2287 527 2321 561
rect 2287 459 2321 493
rect 2287 391 2321 425
rect 2287 323 2321 357
rect 2287 255 2321 289
rect 2287 187 2321 221
rect 2287 119 2321 153
rect 2287 51 2321 85
rect 2287 -17 2321 17
rect 2287 -85 2321 -51
rect 2287 -153 2321 -119
rect 2287 -221 2321 -187
rect 2287 -289 2321 -255
rect 2287 -357 2321 -323
rect 2287 -425 2321 -391
rect 2287 -493 2321 -459
rect 2287 -561 2321 -527
rect 2287 -629 2321 -595
rect 2287 -697 2321 -663
rect 2287 -765 2321 -731
rect 2287 -833 2321 -799
rect 2287 -901 2321 -867
rect 2287 -969 2321 -935
rect 2383 935 2417 969
rect 2383 867 2417 901
rect 2383 799 2417 833
rect 2383 731 2417 765
rect 2383 663 2417 697
rect 2383 595 2417 629
rect 2383 527 2417 561
rect 2383 459 2417 493
rect 2383 391 2417 425
rect 2383 323 2417 357
rect 2383 255 2417 289
rect 2383 187 2417 221
rect 2383 119 2417 153
rect 2383 51 2417 85
rect 2383 -17 2417 17
rect 2383 -85 2417 -51
rect 2383 -153 2417 -119
rect 2383 -221 2417 -187
rect 2383 -289 2417 -255
rect 2383 -357 2417 -323
rect 2383 -425 2417 -391
rect 2383 -493 2417 -459
rect 2383 -561 2417 -527
rect 2383 -629 2417 -595
rect 2383 -697 2417 -663
rect 2383 -765 2417 -731
rect 2383 -833 2417 -799
rect 2383 -901 2417 -867
rect 2383 -969 2417 -935
rect 2479 935 2513 969
rect 2479 867 2513 901
rect 2479 799 2513 833
rect 2479 731 2513 765
rect 2479 663 2513 697
rect 2479 595 2513 629
rect 2479 527 2513 561
rect 2479 459 2513 493
rect 2479 391 2513 425
rect 2479 323 2513 357
rect 2479 255 2513 289
rect 2479 187 2513 221
rect 2479 119 2513 153
rect 2479 51 2513 85
rect 2479 -17 2513 17
rect 2479 -85 2513 -51
rect 2479 -153 2513 -119
rect 2479 -221 2513 -187
rect 2479 -289 2513 -255
rect 2479 -357 2513 -323
rect 2479 -425 2513 -391
rect 2479 -493 2513 -459
rect 2479 -561 2513 -527
rect 2479 -629 2513 -595
rect 2479 -697 2513 -663
rect 2479 -765 2513 -731
rect 2479 -833 2513 -799
rect 2479 -901 2513 -867
rect 2479 -969 2513 -935
rect 2575 935 2609 969
rect 2575 867 2609 901
rect 2575 799 2609 833
rect 2575 731 2609 765
rect 2575 663 2609 697
rect 2575 595 2609 629
rect 2575 527 2609 561
rect 2575 459 2609 493
rect 2575 391 2609 425
rect 2575 323 2609 357
rect 2575 255 2609 289
rect 2575 187 2609 221
rect 2575 119 2609 153
rect 2575 51 2609 85
rect 2575 -17 2609 17
rect 2575 -85 2609 -51
rect 2575 -153 2609 -119
rect 2575 -221 2609 -187
rect 2575 -289 2609 -255
rect 2575 -357 2609 -323
rect 2575 -425 2609 -391
rect 2575 -493 2609 -459
rect 2575 -561 2609 -527
rect 2575 -629 2609 -595
rect 2575 -697 2609 -663
rect 2575 -765 2609 -731
rect 2575 -833 2609 -799
rect 2575 -901 2609 -867
rect 2575 -969 2609 -935
rect 2671 935 2705 969
rect 2671 867 2705 901
rect 2671 799 2705 833
rect 2671 731 2705 765
rect 2671 663 2705 697
rect 2671 595 2705 629
rect 2671 527 2705 561
rect 2671 459 2705 493
rect 2671 391 2705 425
rect 2671 323 2705 357
rect 2671 255 2705 289
rect 2671 187 2705 221
rect 2671 119 2705 153
rect 2671 51 2705 85
rect 2671 -17 2705 17
rect 2671 -85 2705 -51
rect 2671 -153 2705 -119
rect 2671 -221 2705 -187
rect 2671 -289 2705 -255
rect 2671 -357 2705 -323
rect 2671 -425 2705 -391
rect 2671 -493 2705 -459
rect 2671 -561 2705 -527
rect 2671 -629 2705 -595
rect 2671 -697 2705 -663
rect 2671 -765 2705 -731
rect 2671 -833 2705 -799
rect 2671 -901 2705 -867
rect 2671 -969 2705 -935
rect 2767 935 2801 969
rect 2767 867 2801 901
rect 2767 799 2801 833
rect 2767 731 2801 765
rect 2767 663 2801 697
rect 2767 595 2801 629
rect 2767 527 2801 561
rect 2767 459 2801 493
rect 2767 391 2801 425
rect 2767 323 2801 357
rect 2767 255 2801 289
rect 2767 187 2801 221
rect 2767 119 2801 153
rect 2767 51 2801 85
rect 2767 -17 2801 17
rect 2767 -85 2801 -51
rect 2767 -153 2801 -119
rect 2767 -221 2801 -187
rect 2767 -289 2801 -255
rect 2767 -357 2801 -323
rect 2767 -425 2801 -391
rect 2767 -493 2801 -459
rect 2767 -561 2801 -527
rect 2767 -629 2801 -595
rect 2767 -697 2801 -663
rect 2767 -765 2801 -731
rect 2767 -833 2801 -799
rect 2767 -901 2801 -867
rect 2767 -969 2801 -935
rect 2863 935 2897 969
rect 2863 867 2897 901
rect 2863 799 2897 833
rect 2863 731 2897 765
rect 2863 663 2897 697
rect 2863 595 2897 629
rect 2863 527 2897 561
rect 2863 459 2897 493
rect 2863 391 2897 425
rect 2863 323 2897 357
rect 2863 255 2897 289
rect 2863 187 2897 221
rect 2863 119 2897 153
rect 2863 51 2897 85
rect 2863 -17 2897 17
rect 2863 -85 2897 -51
rect 2863 -153 2897 -119
rect 2863 -221 2897 -187
rect 2863 -289 2897 -255
rect 2863 -357 2897 -323
rect 2863 -425 2897 -391
rect 2863 -493 2897 -459
rect 2863 -561 2897 -527
rect 2863 -629 2897 -595
rect 2863 -697 2897 -663
rect 2863 -765 2897 -731
rect 2863 -833 2897 -799
rect 2863 -901 2897 -867
rect 2863 -969 2897 -935
rect 2959 935 2993 969
rect 2959 867 2993 901
rect 2959 799 2993 833
rect 2959 731 2993 765
rect 2959 663 2993 697
rect 2959 595 2993 629
rect 2959 527 2993 561
rect 2959 459 2993 493
rect 2959 391 2993 425
rect 2959 323 2993 357
rect 2959 255 2993 289
rect 2959 187 2993 221
rect 2959 119 2993 153
rect 2959 51 2993 85
rect 2959 -17 2993 17
rect 2959 -85 2993 -51
rect 2959 -153 2993 -119
rect 2959 -221 2993 -187
rect 2959 -289 2993 -255
rect 2959 -357 2993 -323
rect 2959 -425 2993 -391
rect 2959 -493 2993 -459
rect 2959 -561 2993 -527
rect 2959 -629 2993 -595
rect 2959 -697 2993 -663
rect 2959 -765 2993 -731
rect 2959 -833 2993 -799
rect 2959 -901 2993 -867
rect 2959 -969 2993 -935
rect 3055 935 3089 969
rect 3055 867 3089 901
rect 3055 799 3089 833
rect 3055 731 3089 765
rect 3055 663 3089 697
rect 3055 595 3089 629
rect 3055 527 3089 561
rect 3055 459 3089 493
rect 3055 391 3089 425
rect 3055 323 3089 357
rect 3055 255 3089 289
rect 3055 187 3089 221
rect 3055 119 3089 153
rect 3055 51 3089 85
rect 3055 -17 3089 17
rect 3055 -85 3089 -51
rect 3055 -153 3089 -119
rect 3055 -221 3089 -187
rect 3055 -289 3089 -255
rect 3055 -357 3089 -323
rect 3055 -425 3089 -391
rect 3055 -493 3089 -459
rect 3055 -561 3089 -527
rect 3055 -629 3089 -595
rect 3055 -697 3089 -663
rect 3055 -765 3089 -731
rect 3055 -833 3089 -799
rect 3055 -901 3089 -867
rect 3055 -969 3089 -935
rect 3151 935 3185 969
rect 3151 867 3185 901
rect 3151 799 3185 833
rect 3151 731 3185 765
rect 3151 663 3185 697
rect 3151 595 3185 629
rect 3151 527 3185 561
rect 3151 459 3185 493
rect 3151 391 3185 425
rect 3151 323 3185 357
rect 3151 255 3185 289
rect 3151 187 3185 221
rect 3151 119 3185 153
rect 3151 51 3185 85
rect 3151 -17 3185 17
rect 3151 -85 3185 -51
rect 3151 -153 3185 -119
rect 3151 -221 3185 -187
rect 3151 -289 3185 -255
rect 3151 -357 3185 -323
rect 3151 -425 3185 -391
rect 3151 -493 3185 -459
rect 3151 -561 3185 -527
rect 3151 -629 3185 -595
rect 3151 -697 3185 -663
rect 3151 -765 3185 -731
rect 3151 -833 3185 -799
rect 3151 -901 3185 -867
rect 3151 -969 3185 -935
rect 3247 935 3281 969
rect 3247 867 3281 901
rect 3247 799 3281 833
rect 3247 731 3281 765
rect 3247 663 3281 697
rect 3247 595 3281 629
rect 3247 527 3281 561
rect 3247 459 3281 493
rect 3247 391 3281 425
rect 3247 323 3281 357
rect 3247 255 3281 289
rect 3247 187 3281 221
rect 3247 119 3281 153
rect 3247 51 3281 85
rect 3247 -17 3281 17
rect 3247 -85 3281 -51
rect 3247 -153 3281 -119
rect 3247 -221 3281 -187
rect 3247 -289 3281 -255
rect 3247 -357 3281 -323
rect 3247 -425 3281 -391
rect 3247 -493 3281 -459
rect 3247 -561 3281 -527
rect 3247 -629 3281 -595
rect 3247 -697 3281 -663
rect 3247 -765 3281 -731
rect 3247 -833 3281 -799
rect 3247 -901 3281 -867
rect 3247 -969 3281 -935
rect 3343 935 3377 969
rect 3343 867 3377 901
rect 3343 799 3377 833
rect 3343 731 3377 765
rect 3343 663 3377 697
rect 3343 595 3377 629
rect 3343 527 3377 561
rect 3343 459 3377 493
rect 3343 391 3377 425
rect 3343 323 3377 357
rect 3343 255 3377 289
rect 3343 187 3377 221
rect 3343 119 3377 153
rect 3343 51 3377 85
rect 3343 -17 3377 17
rect 3343 -85 3377 -51
rect 3343 -153 3377 -119
rect 3343 -221 3377 -187
rect 3343 -289 3377 -255
rect 3343 -357 3377 -323
rect 3343 -425 3377 -391
rect 3343 -493 3377 -459
rect 3343 -561 3377 -527
rect 3343 -629 3377 -595
rect 3343 -697 3377 -663
rect 3343 -765 3377 -731
rect 3343 -833 3377 -799
rect 3343 -901 3377 -867
rect 3343 -969 3377 -935
rect 3439 935 3473 969
rect 3439 867 3473 901
rect 3439 799 3473 833
rect 3439 731 3473 765
rect 3439 663 3473 697
rect 3439 595 3473 629
rect 3439 527 3473 561
rect 3439 459 3473 493
rect 3439 391 3473 425
rect 3439 323 3473 357
rect 3439 255 3473 289
rect 3439 187 3473 221
rect 3439 119 3473 153
rect 3439 51 3473 85
rect 3439 -17 3473 17
rect 3439 -85 3473 -51
rect 3439 -153 3473 -119
rect 3439 -221 3473 -187
rect 3439 -289 3473 -255
rect 3439 -357 3473 -323
rect 3439 -425 3473 -391
rect 3439 -493 3473 -459
rect 3439 -561 3473 -527
rect 3439 -629 3473 -595
rect 3439 -697 3473 -663
rect 3439 -765 3473 -731
rect 3439 -833 3473 -799
rect 3439 -901 3473 -867
rect 3439 -969 3473 -935
rect 3535 935 3569 969
rect 3535 867 3569 901
rect 3535 799 3569 833
rect 3535 731 3569 765
rect 3535 663 3569 697
rect 3535 595 3569 629
rect 3535 527 3569 561
rect 3535 459 3569 493
rect 3535 391 3569 425
rect 3535 323 3569 357
rect 3535 255 3569 289
rect 3535 187 3569 221
rect 3535 119 3569 153
rect 3535 51 3569 85
rect 3535 -17 3569 17
rect 3535 -85 3569 -51
rect 3535 -153 3569 -119
rect 3535 -221 3569 -187
rect 3535 -289 3569 -255
rect 3535 -357 3569 -323
rect 3535 -425 3569 -391
rect 3535 -493 3569 -459
rect 3535 -561 3569 -527
rect 3535 -629 3569 -595
rect 3535 -697 3569 -663
rect 3535 -765 3569 -731
rect 3535 -833 3569 -799
rect 3535 -901 3569 -867
rect 3535 -969 3569 -935
rect 3631 935 3665 969
rect 3631 867 3665 901
rect 3631 799 3665 833
rect 3631 731 3665 765
rect 3631 663 3665 697
rect 3631 595 3665 629
rect 3631 527 3665 561
rect 3631 459 3665 493
rect 3631 391 3665 425
rect 3631 323 3665 357
rect 3631 255 3665 289
rect 3631 187 3665 221
rect 3631 119 3665 153
rect 3631 51 3665 85
rect 3631 -17 3665 17
rect 3631 -85 3665 -51
rect 3631 -153 3665 -119
rect 3631 -221 3665 -187
rect 3631 -289 3665 -255
rect 3631 -357 3665 -323
rect 3631 -425 3665 -391
rect 3631 -493 3665 -459
rect 3631 -561 3665 -527
rect 3631 -629 3665 -595
rect 3631 -697 3665 -663
rect 3631 -765 3665 -731
rect 3631 -833 3665 -799
rect 3631 -901 3665 -867
rect 3631 -969 3665 -935
rect 3727 935 3761 969
rect 3727 867 3761 901
rect 3727 799 3761 833
rect 3727 731 3761 765
rect 3727 663 3761 697
rect 3727 595 3761 629
rect 3727 527 3761 561
rect 3727 459 3761 493
rect 3727 391 3761 425
rect 3727 323 3761 357
rect 3727 255 3761 289
rect 3727 187 3761 221
rect 3727 119 3761 153
rect 3727 51 3761 85
rect 3727 -17 3761 17
rect 3727 -85 3761 -51
rect 3727 -153 3761 -119
rect 3727 -221 3761 -187
rect 3727 -289 3761 -255
rect 3727 -357 3761 -323
rect 3727 -425 3761 -391
rect 3727 -493 3761 -459
rect 3727 -561 3761 -527
rect 3727 -629 3761 -595
rect 3727 -697 3761 -663
rect 3727 -765 3761 -731
rect 3727 -833 3761 -799
rect 3727 -901 3761 -867
rect 3727 -969 3761 -935
rect 3823 935 3857 969
rect 3823 867 3857 901
rect 3823 799 3857 833
rect 3823 731 3857 765
rect 3823 663 3857 697
rect 3823 595 3857 629
rect 3823 527 3857 561
rect 3823 459 3857 493
rect 3823 391 3857 425
rect 3823 323 3857 357
rect 3823 255 3857 289
rect 3823 187 3857 221
rect 3823 119 3857 153
rect 3823 51 3857 85
rect 3823 -17 3857 17
rect 3823 -85 3857 -51
rect 3823 -153 3857 -119
rect 3823 -221 3857 -187
rect 3823 -289 3857 -255
rect 3823 -357 3857 -323
rect 3823 -425 3857 -391
rect 3823 -493 3857 -459
rect 3823 -561 3857 -527
rect 3823 -629 3857 -595
rect 3823 -697 3857 -663
rect 3823 -765 3857 -731
rect 3823 -833 3857 -799
rect 3823 -901 3857 -867
rect 3823 -969 3857 -935
rect 3919 935 3953 969
rect 3919 867 3953 901
rect 3919 799 3953 833
rect 3919 731 3953 765
rect 3919 663 3953 697
rect 3919 595 3953 629
rect 3919 527 3953 561
rect 3919 459 3953 493
rect 3919 391 3953 425
rect 3919 323 3953 357
rect 3919 255 3953 289
rect 3919 187 3953 221
rect 3919 119 3953 153
rect 3919 51 3953 85
rect 3919 -17 3953 17
rect 3919 -85 3953 -51
rect 3919 -153 3953 -119
rect 3919 -221 3953 -187
rect 3919 -289 3953 -255
rect 3919 -357 3953 -323
rect 3919 -425 3953 -391
rect 3919 -493 3953 -459
rect 3919 -561 3953 -527
rect 3919 -629 3953 -595
rect 3919 -697 3953 -663
rect 3919 -765 3953 -731
rect 3919 -833 3953 -799
rect 3919 -901 3953 -867
rect 3919 -969 3953 -935
rect 4015 935 4049 969
rect 4015 867 4049 901
rect 4015 799 4049 833
rect 4015 731 4049 765
rect 4015 663 4049 697
rect 4015 595 4049 629
rect 4015 527 4049 561
rect 4015 459 4049 493
rect 4015 391 4049 425
rect 4015 323 4049 357
rect 4015 255 4049 289
rect 4015 187 4049 221
rect 4015 119 4049 153
rect 4015 51 4049 85
rect 4015 -17 4049 17
rect 4015 -85 4049 -51
rect 4015 -153 4049 -119
rect 4015 -221 4049 -187
rect 4015 -289 4049 -255
rect 4015 -357 4049 -323
rect 4015 -425 4049 -391
rect 4015 -493 4049 -459
rect 4015 -561 4049 -527
rect 4015 -629 4049 -595
rect 4015 -697 4049 -663
rect 4015 -765 4049 -731
rect 4015 -833 4049 -799
rect 4015 -901 4049 -867
rect 4015 -969 4049 -935
rect 4111 935 4145 969
rect 4111 867 4145 901
rect 4111 799 4145 833
rect 4111 731 4145 765
rect 4111 663 4145 697
rect 4111 595 4145 629
rect 4111 527 4145 561
rect 4111 459 4145 493
rect 4111 391 4145 425
rect 4111 323 4145 357
rect 4111 255 4145 289
rect 4111 187 4145 221
rect 4111 119 4145 153
rect 4111 51 4145 85
rect 4111 -17 4145 17
rect 4111 -85 4145 -51
rect 4111 -153 4145 -119
rect 4111 -221 4145 -187
rect 4111 -289 4145 -255
rect 4111 -357 4145 -323
rect 4111 -425 4145 -391
rect 4111 -493 4145 -459
rect 4111 -561 4145 -527
rect 4111 -629 4145 -595
rect 4111 -697 4145 -663
rect 4111 -765 4145 -731
rect 4111 -833 4145 -799
rect 4111 -901 4145 -867
rect 4111 -969 4145 -935
rect 4207 935 4241 969
rect 4207 867 4241 901
rect 4207 799 4241 833
rect 4207 731 4241 765
rect 4207 663 4241 697
rect 4207 595 4241 629
rect 4207 527 4241 561
rect 4207 459 4241 493
rect 4207 391 4241 425
rect 4207 323 4241 357
rect 4207 255 4241 289
rect 4207 187 4241 221
rect 4207 119 4241 153
rect 4207 51 4241 85
rect 4207 -17 4241 17
rect 4207 -85 4241 -51
rect 4207 -153 4241 -119
rect 4207 -221 4241 -187
rect 4207 -289 4241 -255
rect 4207 -357 4241 -323
rect 4207 -425 4241 -391
rect 4207 -493 4241 -459
rect 4207 -561 4241 -527
rect 4207 -629 4241 -595
rect 4207 -697 4241 -663
rect 4207 -765 4241 -731
rect 4207 -833 4241 -799
rect 4207 -901 4241 -867
rect 4207 -969 4241 -935
rect 4303 935 4337 969
rect 4303 867 4337 901
rect 4303 799 4337 833
rect 4303 731 4337 765
rect 4303 663 4337 697
rect 4303 595 4337 629
rect 4303 527 4337 561
rect 4303 459 4337 493
rect 4303 391 4337 425
rect 4303 323 4337 357
rect 4303 255 4337 289
rect 4303 187 4337 221
rect 4303 119 4337 153
rect 4303 51 4337 85
rect 4303 -17 4337 17
rect 4303 -85 4337 -51
rect 4303 -153 4337 -119
rect 4303 -221 4337 -187
rect 4303 -289 4337 -255
rect 4303 -357 4337 -323
rect 4303 -425 4337 -391
rect 4303 -493 4337 -459
rect 4303 -561 4337 -527
rect 4303 -629 4337 -595
rect 4303 -697 4337 -663
rect 4303 -765 4337 -731
rect 4303 -833 4337 -799
rect 4303 -901 4337 -867
rect 4303 -969 4337 -935
rect 4399 935 4433 969
rect 4399 867 4433 901
rect 4399 799 4433 833
rect 4399 731 4433 765
rect 4399 663 4433 697
rect 4399 595 4433 629
rect 4399 527 4433 561
rect 4399 459 4433 493
rect 4399 391 4433 425
rect 4399 323 4433 357
rect 4399 255 4433 289
rect 4399 187 4433 221
rect 4399 119 4433 153
rect 4399 51 4433 85
rect 4399 -17 4433 17
rect 4399 -85 4433 -51
rect 4399 -153 4433 -119
rect 4399 -221 4433 -187
rect 4399 -289 4433 -255
rect 4399 -357 4433 -323
rect 4399 -425 4433 -391
rect 4399 -493 4433 -459
rect 4399 -561 4433 -527
rect 4399 -629 4433 -595
rect 4399 -697 4433 -663
rect 4399 -765 4433 -731
rect 4399 -833 4433 -799
rect 4399 -901 4433 -867
rect 4399 -969 4433 -935
rect 4495 935 4529 969
rect 4495 867 4529 901
rect 4495 799 4529 833
rect 4495 731 4529 765
rect 4495 663 4529 697
rect 4495 595 4529 629
rect 4495 527 4529 561
rect 4495 459 4529 493
rect 4495 391 4529 425
rect 4495 323 4529 357
rect 4495 255 4529 289
rect 4495 187 4529 221
rect 4495 119 4529 153
rect 4495 51 4529 85
rect 4495 -17 4529 17
rect 4495 -85 4529 -51
rect 4495 -153 4529 -119
rect 4495 -221 4529 -187
rect 4495 -289 4529 -255
rect 4495 -357 4529 -323
rect 4495 -425 4529 -391
rect 4495 -493 4529 -459
rect 4495 -561 4529 -527
rect 4495 -629 4529 -595
rect 4495 -697 4529 -663
rect 4495 -765 4529 -731
rect 4495 -833 4529 -799
rect 4495 -901 4529 -867
rect 4495 -969 4529 -935
rect 4591 935 4625 969
rect 4591 867 4625 901
rect 4591 799 4625 833
rect 4591 731 4625 765
rect 4591 663 4625 697
rect 4591 595 4625 629
rect 4591 527 4625 561
rect 4591 459 4625 493
rect 4591 391 4625 425
rect 4591 323 4625 357
rect 4591 255 4625 289
rect 4591 187 4625 221
rect 4591 119 4625 153
rect 4591 51 4625 85
rect 4591 -17 4625 17
rect 4591 -85 4625 -51
rect 4591 -153 4625 -119
rect 4591 -221 4625 -187
rect 4591 -289 4625 -255
rect 4591 -357 4625 -323
rect 4591 -425 4625 -391
rect 4591 -493 4625 -459
rect 4591 -561 4625 -527
rect 4591 -629 4625 -595
rect 4591 -697 4625 -663
rect 4591 -765 4625 -731
rect 4591 -833 4625 -799
rect 4591 -901 4625 -867
rect 4591 -969 4625 -935
rect 4687 935 4721 969
rect 4687 867 4721 901
rect 4687 799 4721 833
rect 4687 731 4721 765
rect 4687 663 4721 697
rect 4687 595 4721 629
rect 4687 527 4721 561
rect 4687 459 4721 493
rect 4687 391 4721 425
rect 4687 323 4721 357
rect 4687 255 4721 289
rect 4687 187 4721 221
rect 4687 119 4721 153
rect 4687 51 4721 85
rect 4687 -17 4721 17
rect 4687 -85 4721 -51
rect 4687 -153 4721 -119
rect 4687 -221 4721 -187
rect 4687 -289 4721 -255
rect 4687 -357 4721 -323
rect 4687 -425 4721 -391
rect 4687 -493 4721 -459
rect 4687 -561 4721 -527
rect 4687 -629 4721 -595
rect 4687 -697 4721 -663
rect 4687 -765 4721 -731
rect 4687 -833 4721 -799
rect 4687 -901 4721 -867
rect 4687 -969 4721 -935
rect 4783 935 4817 969
rect 4783 867 4817 901
rect 4783 799 4817 833
rect 4783 731 4817 765
rect 4783 663 4817 697
rect 4783 595 4817 629
rect 4783 527 4817 561
rect 4783 459 4817 493
rect 4783 391 4817 425
rect 4783 323 4817 357
rect 4783 255 4817 289
rect 4783 187 4817 221
rect 4783 119 4817 153
rect 4783 51 4817 85
rect 4783 -17 4817 17
rect 4783 -85 4817 -51
rect 4783 -153 4817 -119
rect 4783 -221 4817 -187
rect 4783 -289 4817 -255
rect 4783 -357 4817 -323
rect 4783 -425 4817 -391
rect 4783 -493 4817 -459
rect 4783 -561 4817 -527
rect 4783 -629 4817 -595
rect 4783 -697 4817 -663
rect 4783 -765 4817 -731
rect 4783 -833 4817 -799
rect 4783 -901 4817 -867
rect 4783 -969 4817 -935
<< psubdiff >>
rect -4931 1140 -4811 1174
rect -4777 1140 -4743 1174
rect -4709 1140 -4675 1174
rect -4641 1140 -4607 1174
rect -4573 1140 -4539 1174
rect -4505 1140 -4471 1174
rect -4437 1140 -4403 1174
rect -4369 1140 -4335 1174
rect -4301 1140 -4267 1174
rect -4233 1140 -4199 1174
rect -4165 1140 -4131 1174
rect -4097 1140 -4063 1174
rect -4029 1140 -3995 1174
rect -3961 1140 -3927 1174
rect -3893 1140 -3859 1174
rect -3825 1140 -3791 1174
rect -3757 1140 -3723 1174
rect -3689 1140 -3655 1174
rect -3621 1140 -3587 1174
rect -3553 1140 -3519 1174
rect -3485 1140 -3451 1174
rect -3417 1140 -3383 1174
rect -3349 1140 -3315 1174
rect -3281 1140 -3247 1174
rect -3213 1140 -3179 1174
rect -3145 1140 -3111 1174
rect -3077 1140 -3043 1174
rect -3009 1140 -2975 1174
rect -2941 1140 -2907 1174
rect -2873 1140 -2839 1174
rect -2805 1140 -2771 1174
rect -2737 1140 -2703 1174
rect -2669 1140 -2635 1174
rect -2601 1140 -2567 1174
rect -2533 1140 -2499 1174
rect -2465 1140 -2431 1174
rect -2397 1140 -2363 1174
rect -2329 1140 -2295 1174
rect -2261 1140 -2227 1174
rect -2193 1140 -2159 1174
rect -2125 1140 -2091 1174
rect -2057 1140 -2023 1174
rect -1989 1140 -1955 1174
rect -1921 1140 -1887 1174
rect -1853 1140 -1819 1174
rect -1785 1140 -1751 1174
rect -1717 1140 -1683 1174
rect -1649 1140 -1615 1174
rect -1581 1140 -1547 1174
rect -1513 1140 -1479 1174
rect -1445 1140 -1411 1174
rect -1377 1140 -1343 1174
rect -1309 1140 -1275 1174
rect -1241 1140 -1207 1174
rect -1173 1140 -1139 1174
rect -1105 1140 -1071 1174
rect -1037 1140 -1003 1174
rect -969 1140 -935 1174
rect -901 1140 -867 1174
rect -833 1140 -799 1174
rect -765 1140 -731 1174
rect -697 1140 -663 1174
rect -629 1140 -595 1174
rect -561 1140 -527 1174
rect -493 1140 -459 1174
rect -425 1140 -391 1174
rect -357 1140 -323 1174
rect -289 1140 -255 1174
rect -221 1140 -187 1174
rect -153 1140 -119 1174
rect -85 1140 -51 1174
rect -17 1140 17 1174
rect 51 1140 85 1174
rect 119 1140 153 1174
rect 187 1140 221 1174
rect 255 1140 289 1174
rect 323 1140 357 1174
rect 391 1140 425 1174
rect 459 1140 493 1174
rect 527 1140 561 1174
rect 595 1140 629 1174
rect 663 1140 697 1174
rect 731 1140 765 1174
rect 799 1140 833 1174
rect 867 1140 901 1174
rect 935 1140 969 1174
rect 1003 1140 1037 1174
rect 1071 1140 1105 1174
rect 1139 1140 1173 1174
rect 1207 1140 1241 1174
rect 1275 1140 1309 1174
rect 1343 1140 1377 1174
rect 1411 1140 1445 1174
rect 1479 1140 1513 1174
rect 1547 1140 1581 1174
rect 1615 1140 1649 1174
rect 1683 1140 1717 1174
rect 1751 1140 1785 1174
rect 1819 1140 1853 1174
rect 1887 1140 1921 1174
rect 1955 1140 1989 1174
rect 2023 1140 2057 1174
rect 2091 1140 2125 1174
rect 2159 1140 2193 1174
rect 2227 1140 2261 1174
rect 2295 1140 2329 1174
rect 2363 1140 2397 1174
rect 2431 1140 2465 1174
rect 2499 1140 2533 1174
rect 2567 1140 2601 1174
rect 2635 1140 2669 1174
rect 2703 1140 2737 1174
rect 2771 1140 2805 1174
rect 2839 1140 2873 1174
rect 2907 1140 2941 1174
rect 2975 1140 3009 1174
rect 3043 1140 3077 1174
rect 3111 1140 3145 1174
rect 3179 1140 3213 1174
rect 3247 1140 3281 1174
rect 3315 1140 3349 1174
rect 3383 1140 3417 1174
rect 3451 1140 3485 1174
rect 3519 1140 3553 1174
rect 3587 1140 3621 1174
rect 3655 1140 3689 1174
rect 3723 1140 3757 1174
rect 3791 1140 3825 1174
rect 3859 1140 3893 1174
rect 3927 1140 3961 1174
rect 3995 1140 4029 1174
rect 4063 1140 4097 1174
rect 4131 1140 4165 1174
rect 4199 1140 4233 1174
rect 4267 1140 4301 1174
rect 4335 1140 4369 1174
rect 4403 1140 4437 1174
rect 4471 1140 4505 1174
rect 4539 1140 4573 1174
rect 4607 1140 4641 1174
rect 4675 1140 4709 1174
rect 4743 1140 4777 1174
rect 4811 1140 4931 1174
rect -4931 1071 -4897 1140
rect -4931 1003 -4897 1037
rect 4897 1071 4931 1140
rect 4897 1003 4931 1037
rect -4931 935 -4897 969
rect -4931 867 -4897 901
rect -4931 799 -4897 833
rect -4931 731 -4897 765
rect -4931 663 -4897 697
rect -4931 595 -4897 629
rect -4931 527 -4897 561
rect -4931 459 -4897 493
rect -4931 391 -4897 425
rect -4931 323 -4897 357
rect -4931 255 -4897 289
rect -4931 187 -4897 221
rect -4931 119 -4897 153
rect -4931 51 -4897 85
rect -4931 -17 -4897 17
rect -4931 -85 -4897 -51
rect -4931 -153 -4897 -119
rect -4931 -221 -4897 -187
rect -4931 -289 -4897 -255
rect -4931 -357 -4897 -323
rect -4931 -425 -4897 -391
rect -4931 -493 -4897 -459
rect -4931 -561 -4897 -527
rect -4931 -629 -4897 -595
rect -4931 -697 -4897 -663
rect -4931 -765 -4897 -731
rect -4931 -833 -4897 -799
rect -4931 -901 -4897 -867
rect -4931 -969 -4897 -935
rect 4897 935 4931 969
rect 4897 867 4931 901
rect 4897 799 4931 833
rect 4897 731 4931 765
rect 4897 663 4931 697
rect 4897 595 4931 629
rect 4897 527 4931 561
rect 4897 459 4931 493
rect 4897 391 4931 425
rect 4897 323 4931 357
rect 4897 255 4931 289
rect 4897 187 4931 221
rect 4897 119 4931 153
rect 4897 51 4931 85
rect 4897 -17 4931 17
rect 4897 -85 4931 -51
rect 4897 -153 4931 -119
rect 4897 -221 4931 -187
rect 4897 -289 4931 -255
rect 4897 -357 4931 -323
rect 4897 -425 4931 -391
rect 4897 -493 4931 -459
rect 4897 -561 4931 -527
rect 4897 -629 4931 -595
rect 4897 -697 4931 -663
rect 4897 -765 4931 -731
rect 4897 -833 4931 -799
rect 4897 -901 4931 -867
rect 4897 -969 4931 -935
rect -4931 -1037 -4897 -1003
rect -4931 -1140 -4897 -1071
rect 4897 -1037 4931 -1003
rect 4897 -1140 4931 -1071
rect -4931 -1174 -4811 -1140
rect -4777 -1174 -4743 -1140
rect -4709 -1174 -4675 -1140
rect -4641 -1174 -4607 -1140
rect -4573 -1174 -4539 -1140
rect -4505 -1174 -4471 -1140
rect -4437 -1174 -4403 -1140
rect -4369 -1174 -4335 -1140
rect -4301 -1174 -4267 -1140
rect -4233 -1174 -4199 -1140
rect -4165 -1174 -4131 -1140
rect -4097 -1174 -4063 -1140
rect -4029 -1174 -3995 -1140
rect -3961 -1174 -3927 -1140
rect -3893 -1174 -3859 -1140
rect -3825 -1174 -3791 -1140
rect -3757 -1174 -3723 -1140
rect -3689 -1174 -3655 -1140
rect -3621 -1174 -3587 -1140
rect -3553 -1174 -3519 -1140
rect -3485 -1174 -3451 -1140
rect -3417 -1174 -3383 -1140
rect -3349 -1174 -3315 -1140
rect -3281 -1174 -3247 -1140
rect -3213 -1174 -3179 -1140
rect -3145 -1174 -3111 -1140
rect -3077 -1174 -3043 -1140
rect -3009 -1174 -2975 -1140
rect -2941 -1174 -2907 -1140
rect -2873 -1174 -2839 -1140
rect -2805 -1174 -2771 -1140
rect -2737 -1174 -2703 -1140
rect -2669 -1174 -2635 -1140
rect -2601 -1174 -2567 -1140
rect -2533 -1174 -2499 -1140
rect -2465 -1174 -2431 -1140
rect -2397 -1174 -2363 -1140
rect -2329 -1174 -2295 -1140
rect -2261 -1174 -2227 -1140
rect -2193 -1174 -2159 -1140
rect -2125 -1174 -2091 -1140
rect -2057 -1174 -2023 -1140
rect -1989 -1174 -1955 -1140
rect -1921 -1174 -1887 -1140
rect -1853 -1174 -1819 -1140
rect -1785 -1174 -1751 -1140
rect -1717 -1174 -1683 -1140
rect -1649 -1174 -1615 -1140
rect -1581 -1174 -1547 -1140
rect -1513 -1174 -1479 -1140
rect -1445 -1174 -1411 -1140
rect -1377 -1174 -1343 -1140
rect -1309 -1174 -1275 -1140
rect -1241 -1174 -1207 -1140
rect -1173 -1174 -1139 -1140
rect -1105 -1174 -1071 -1140
rect -1037 -1174 -1003 -1140
rect -969 -1174 -935 -1140
rect -901 -1174 -867 -1140
rect -833 -1174 -799 -1140
rect -765 -1174 -731 -1140
rect -697 -1174 -663 -1140
rect -629 -1174 -595 -1140
rect -561 -1174 -527 -1140
rect -493 -1174 -459 -1140
rect -425 -1174 -391 -1140
rect -357 -1174 -323 -1140
rect -289 -1174 -255 -1140
rect -221 -1174 -187 -1140
rect -153 -1174 -119 -1140
rect -85 -1174 -51 -1140
rect -17 -1174 17 -1140
rect 51 -1174 85 -1140
rect 119 -1174 153 -1140
rect 187 -1174 221 -1140
rect 255 -1174 289 -1140
rect 323 -1174 357 -1140
rect 391 -1174 425 -1140
rect 459 -1174 493 -1140
rect 527 -1174 561 -1140
rect 595 -1174 629 -1140
rect 663 -1174 697 -1140
rect 731 -1174 765 -1140
rect 799 -1174 833 -1140
rect 867 -1174 901 -1140
rect 935 -1174 969 -1140
rect 1003 -1174 1037 -1140
rect 1071 -1174 1105 -1140
rect 1139 -1174 1173 -1140
rect 1207 -1174 1241 -1140
rect 1275 -1174 1309 -1140
rect 1343 -1174 1377 -1140
rect 1411 -1174 1445 -1140
rect 1479 -1174 1513 -1140
rect 1547 -1174 1581 -1140
rect 1615 -1174 1649 -1140
rect 1683 -1174 1717 -1140
rect 1751 -1174 1785 -1140
rect 1819 -1174 1853 -1140
rect 1887 -1174 1921 -1140
rect 1955 -1174 1989 -1140
rect 2023 -1174 2057 -1140
rect 2091 -1174 2125 -1140
rect 2159 -1174 2193 -1140
rect 2227 -1174 2261 -1140
rect 2295 -1174 2329 -1140
rect 2363 -1174 2397 -1140
rect 2431 -1174 2465 -1140
rect 2499 -1174 2533 -1140
rect 2567 -1174 2601 -1140
rect 2635 -1174 2669 -1140
rect 2703 -1174 2737 -1140
rect 2771 -1174 2805 -1140
rect 2839 -1174 2873 -1140
rect 2907 -1174 2941 -1140
rect 2975 -1174 3009 -1140
rect 3043 -1174 3077 -1140
rect 3111 -1174 3145 -1140
rect 3179 -1174 3213 -1140
rect 3247 -1174 3281 -1140
rect 3315 -1174 3349 -1140
rect 3383 -1174 3417 -1140
rect 3451 -1174 3485 -1140
rect 3519 -1174 3553 -1140
rect 3587 -1174 3621 -1140
rect 3655 -1174 3689 -1140
rect 3723 -1174 3757 -1140
rect 3791 -1174 3825 -1140
rect 3859 -1174 3893 -1140
rect 3927 -1174 3961 -1140
rect 3995 -1174 4029 -1140
rect 4063 -1174 4097 -1140
rect 4131 -1174 4165 -1140
rect 4199 -1174 4233 -1140
rect 4267 -1174 4301 -1140
rect 4335 -1174 4369 -1140
rect 4403 -1174 4437 -1140
rect 4471 -1174 4505 -1140
rect 4539 -1174 4573 -1140
rect 4607 -1174 4641 -1140
rect 4675 -1174 4709 -1140
rect 4743 -1174 4777 -1140
rect 4811 -1174 4931 -1140
<< psubdiffcont >>
rect -4811 1140 -4777 1174
rect -4743 1140 -4709 1174
rect -4675 1140 -4641 1174
rect -4607 1140 -4573 1174
rect -4539 1140 -4505 1174
rect -4471 1140 -4437 1174
rect -4403 1140 -4369 1174
rect -4335 1140 -4301 1174
rect -4267 1140 -4233 1174
rect -4199 1140 -4165 1174
rect -4131 1140 -4097 1174
rect -4063 1140 -4029 1174
rect -3995 1140 -3961 1174
rect -3927 1140 -3893 1174
rect -3859 1140 -3825 1174
rect -3791 1140 -3757 1174
rect -3723 1140 -3689 1174
rect -3655 1140 -3621 1174
rect -3587 1140 -3553 1174
rect -3519 1140 -3485 1174
rect -3451 1140 -3417 1174
rect -3383 1140 -3349 1174
rect -3315 1140 -3281 1174
rect -3247 1140 -3213 1174
rect -3179 1140 -3145 1174
rect -3111 1140 -3077 1174
rect -3043 1140 -3009 1174
rect -2975 1140 -2941 1174
rect -2907 1140 -2873 1174
rect -2839 1140 -2805 1174
rect -2771 1140 -2737 1174
rect -2703 1140 -2669 1174
rect -2635 1140 -2601 1174
rect -2567 1140 -2533 1174
rect -2499 1140 -2465 1174
rect -2431 1140 -2397 1174
rect -2363 1140 -2329 1174
rect -2295 1140 -2261 1174
rect -2227 1140 -2193 1174
rect -2159 1140 -2125 1174
rect -2091 1140 -2057 1174
rect -2023 1140 -1989 1174
rect -1955 1140 -1921 1174
rect -1887 1140 -1853 1174
rect -1819 1140 -1785 1174
rect -1751 1140 -1717 1174
rect -1683 1140 -1649 1174
rect -1615 1140 -1581 1174
rect -1547 1140 -1513 1174
rect -1479 1140 -1445 1174
rect -1411 1140 -1377 1174
rect -1343 1140 -1309 1174
rect -1275 1140 -1241 1174
rect -1207 1140 -1173 1174
rect -1139 1140 -1105 1174
rect -1071 1140 -1037 1174
rect -1003 1140 -969 1174
rect -935 1140 -901 1174
rect -867 1140 -833 1174
rect -799 1140 -765 1174
rect -731 1140 -697 1174
rect -663 1140 -629 1174
rect -595 1140 -561 1174
rect -527 1140 -493 1174
rect -459 1140 -425 1174
rect -391 1140 -357 1174
rect -323 1140 -289 1174
rect -255 1140 -221 1174
rect -187 1140 -153 1174
rect -119 1140 -85 1174
rect -51 1140 -17 1174
rect 17 1140 51 1174
rect 85 1140 119 1174
rect 153 1140 187 1174
rect 221 1140 255 1174
rect 289 1140 323 1174
rect 357 1140 391 1174
rect 425 1140 459 1174
rect 493 1140 527 1174
rect 561 1140 595 1174
rect 629 1140 663 1174
rect 697 1140 731 1174
rect 765 1140 799 1174
rect 833 1140 867 1174
rect 901 1140 935 1174
rect 969 1140 1003 1174
rect 1037 1140 1071 1174
rect 1105 1140 1139 1174
rect 1173 1140 1207 1174
rect 1241 1140 1275 1174
rect 1309 1140 1343 1174
rect 1377 1140 1411 1174
rect 1445 1140 1479 1174
rect 1513 1140 1547 1174
rect 1581 1140 1615 1174
rect 1649 1140 1683 1174
rect 1717 1140 1751 1174
rect 1785 1140 1819 1174
rect 1853 1140 1887 1174
rect 1921 1140 1955 1174
rect 1989 1140 2023 1174
rect 2057 1140 2091 1174
rect 2125 1140 2159 1174
rect 2193 1140 2227 1174
rect 2261 1140 2295 1174
rect 2329 1140 2363 1174
rect 2397 1140 2431 1174
rect 2465 1140 2499 1174
rect 2533 1140 2567 1174
rect 2601 1140 2635 1174
rect 2669 1140 2703 1174
rect 2737 1140 2771 1174
rect 2805 1140 2839 1174
rect 2873 1140 2907 1174
rect 2941 1140 2975 1174
rect 3009 1140 3043 1174
rect 3077 1140 3111 1174
rect 3145 1140 3179 1174
rect 3213 1140 3247 1174
rect 3281 1140 3315 1174
rect 3349 1140 3383 1174
rect 3417 1140 3451 1174
rect 3485 1140 3519 1174
rect 3553 1140 3587 1174
rect 3621 1140 3655 1174
rect 3689 1140 3723 1174
rect 3757 1140 3791 1174
rect 3825 1140 3859 1174
rect 3893 1140 3927 1174
rect 3961 1140 3995 1174
rect 4029 1140 4063 1174
rect 4097 1140 4131 1174
rect 4165 1140 4199 1174
rect 4233 1140 4267 1174
rect 4301 1140 4335 1174
rect 4369 1140 4403 1174
rect 4437 1140 4471 1174
rect 4505 1140 4539 1174
rect 4573 1140 4607 1174
rect 4641 1140 4675 1174
rect 4709 1140 4743 1174
rect 4777 1140 4811 1174
rect -4931 1037 -4897 1071
rect -4931 969 -4897 1003
rect 4897 1037 4931 1071
rect -4931 901 -4897 935
rect -4931 833 -4897 867
rect -4931 765 -4897 799
rect -4931 697 -4897 731
rect -4931 629 -4897 663
rect -4931 561 -4897 595
rect -4931 493 -4897 527
rect -4931 425 -4897 459
rect -4931 357 -4897 391
rect -4931 289 -4897 323
rect -4931 221 -4897 255
rect -4931 153 -4897 187
rect -4931 85 -4897 119
rect -4931 17 -4897 51
rect -4931 -51 -4897 -17
rect -4931 -119 -4897 -85
rect -4931 -187 -4897 -153
rect -4931 -255 -4897 -221
rect -4931 -323 -4897 -289
rect -4931 -391 -4897 -357
rect -4931 -459 -4897 -425
rect -4931 -527 -4897 -493
rect -4931 -595 -4897 -561
rect -4931 -663 -4897 -629
rect -4931 -731 -4897 -697
rect -4931 -799 -4897 -765
rect -4931 -867 -4897 -833
rect -4931 -935 -4897 -901
rect -4931 -1003 -4897 -969
rect 4897 969 4931 1003
rect 4897 901 4931 935
rect 4897 833 4931 867
rect 4897 765 4931 799
rect 4897 697 4931 731
rect 4897 629 4931 663
rect 4897 561 4931 595
rect 4897 493 4931 527
rect 4897 425 4931 459
rect 4897 357 4931 391
rect 4897 289 4931 323
rect 4897 221 4931 255
rect 4897 153 4931 187
rect 4897 85 4931 119
rect 4897 17 4931 51
rect 4897 -51 4931 -17
rect 4897 -119 4931 -85
rect 4897 -187 4931 -153
rect 4897 -255 4931 -221
rect 4897 -323 4931 -289
rect 4897 -391 4931 -357
rect 4897 -459 4931 -425
rect 4897 -527 4931 -493
rect 4897 -595 4931 -561
rect 4897 -663 4931 -629
rect 4897 -731 4931 -697
rect 4897 -799 4931 -765
rect 4897 -867 4931 -833
rect 4897 -935 4931 -901
rect -4931 -1071 -4897 -1037
rect 4897 -1003 4931 -969
rect 4897 -1071 4931 -1037
rect -4811 -1174 -4777 -1140
rect -4743 -1174 -4709 -1140
rect -4675 -1174 -4641 -1140
rect -4607 -1174 -4573 -1140
rect -4539 -1174 -4505 -1140
rect -4471 -1174 -4437 -1140
rect -4403 -1174 -4369 -1140
rect -4335 -1174 -4301 -1140
rect -4267 -1174 -4233 -1140
rect -4199 -1174 -4165 -1140
rect -4131 -1174 -4097 -1140
rect -4063 -1174 -4029 -1140
rect -3995 -1174 -3961 -1140
rect -3927 -1174 -3893 -1140
rect -3859 -1174 -3825 -1140
rect -3791 -1174 -3757 -1140
rect -3723 -1174 -3689 -1140
rect -3655 -1174 -3621 -1140
rect -3587 -1174 -3553 -1140
rect -3519 -1174 -3485 -1140
rect -3451 -1174 -3417 -1140
rect -3383 -1174 -3349 -1140
rect -3315 -1174 -3281 -1140
rect -3247 -1174 -3213 -1140
rect -3179 -1174 -3145 -1140
rect -3111 -1174 -3077 -1140
rect -3043 -1174 -3009 -1140
rect -2975 -1174 -2941 -1140
rect -2907 -1174 -2873 -1140
rect -2839 -1174 -2805 -1140
rect -2771 -1174 -2737 -1140
rect -2703 -1174 -2669 -1140
rect -2635 -1174 -2601 -1140
rect -2567 -1174 -2533 -1140
rect -2499 -1174 -2465 -1140
rect -2431 -1174 -2397 -1140
rect -2363 -1174 -2329 -1140
rect -2295 -1174 -2261 -1140
rect -2227 -1174 -2193 -1140
rect -2159 -1174 -2125 -1140
rect -2091 -1174 -2057 -1140
rect -2023 -1174 -1989 -1140
rect -1955 -1174 -1921 -1140
rect -1887 -1174 -1853 -1140
rect -1819 -1174 -1785 -1140
rect -1751 -1174 -1717 -1140
rect -1683 -1174 -1649 -1140
rect -1615 -1174 -1581 -1140
rect -1547 -1174 -1513 -1140
rect -1479 -1174 -1445 -1140
rect -1411 -1174 -1377 -1140
rect -1343 -1174 -1309 -1140
rect -1275 -1174 -1241 -1140
rect -1207 -1174 -1173 -1140
rect -1139 -1174 -1105 -1140
rect -1071 -1174 -1037 -1140
rect -1003 -1174 -969 -1140
rect -935 -1174 -901 -1140
rect -867 -1174 -833 -1140
rect -799 -1174 -765 -1140
rect -731 -1174 -697 -1140
rect -663 -1174 -629 -1140
rect -595 -1174 -561 -1140
rect -527 -1174 -493 -1140
rect -459 -1174 -425 -1140
rect -391 -1174 -357 -1140
rect -323 -1174 -289 -1140
rect -255 -1174 -221 -1140
rect -187 -1174 -153 -1140
rect -119 -1174 -85 -1140
rect -51 -1174 -17 -1140
rect 17 -1174 51 -1140
rect 85 -1174 119 -1140
rect 153 -1174 187 -1140
rect 221 -1174 255 -1140
rect 289 -1174 323 -1140
rect 357 -1174 391 -1140
rect 425 -1174 459 -1140
rect 493 -1174 527 -1140
rect 561 -1174 595 -1140
rect 629 -1174 663 -1140
rect 697 -1174 731 -1140
rect 765 -1174 799 -1140
rect 833 -1174 867 -1140
rect 901 -1174 935 -1140
rect 969 -1174 1003 -1140
rect 1037 -1174 1071 -1140
rect 1105 -1174 1139 -1140
rect 1173 -1174 1207 -1140
rect 1241 -1174 1275 -1140
rect 1309 -1174 1343 -1140
rect 1377 -1174 1411 -1140
rect 1445 -1174 1479 -1140
rect 1513 -1174 1547 -1140
rect 1581 -1174 1615 -1140
rect 1649 -1174 1683 -1140
rect 1717 -1174 1751 -1140
rect 1785 -1174 1819 -1140
rect 1853 -1174 1887 -1140
rect 1921 -1174 1955 -1140
rect 1989 -1174 2023 -1140
rect 2057 -1174 2091 -1140
rect 2125 -1174 2159 -1140
rect 2193 -1174 2227 -1140
rect 2261 -1174 2295 -1140
rect 2329 -1174 2363 -1140
rect 2397 -1174 2431 -1140
rect 2465 -1174 2499 -1140
rect 2533 -1174 2567 -1140
rect 2601 -1174 2635 -1140
rect 2669 -1174 2703 -1140
rect 2737 -1174 2771 -1140
rect 2805 -1174 2839 -1140
rect 2873 -1174 2907 -1140
rect 2941 -1174 2975 -1140
rect 3009 -1174 3043 -1140
rect 3077 -1174 3111 -1140
rect 3145 -1174 3179 -1140
rect 3213 -1174 3247 -1140
rect 3281 -1174 3315 -1140
rect 3349 -1174 3383 -1140
rect 3417 -1174 3451 -1140
rect 3485 -1174 3519 -1140
rect 3553 -1174 3587 -1140
rect 3621 -1174 3655 -1140
rect 3689 -1174 3723 -1140
rect 3757 -1174 3791 -1140
rect 3825 -1174 3859 -1140
rect 3893 -1174 3927 -1140
rect 3961 -1174 3995 -1140
rect 4029 -1174 4063 -1140
rect 4097 -1174 4131 -1140
rect 4165 -1174 4199 -1140
rect 4233 -1174 4267 -1140
rect 4301 -1174 4335 -1140
rect 4369 -1174 4403 -1140
rect 4437 -1174 4471 -1140
rect 4505 -1174 4539 -1140
rect 4573 -1174 4607 -1140
rect 4641 -1174 4675 -1140
rect 4709 -1174 4743 -1140
rect 4777 -1174 4811 -1140
<< poly >>
rect -4689 1072 -4623 1088
rect -4689 1038 -4673 1072
rect -4639 1038 -4623 1072
rect -4767 1000 -4737 1026
rect -4689 1022 -4623 1038
rect -4497 1072 -4431 1088
rect -4497 1038 -4481 1072
rect -4447 1038 -4431 1072
rect -4671 1000 -4641 1022
rect -4575 1000 -4545 1026
rect -4497 1022 -4431 1038
rect -4305 1072 -4239 1088
rect -4305 1038 -4289 1072
rect -4255 1038 -4239 1072
rect -4479 1000 -4449 1022
rect -4383 1000 -4353 1026
rect -4305 1022 -4239 1038
rect -4113 1072 -4047 1088
rect -4113 1038 -4097 1072
rect -4063 1038 -4047 1072
rect -4287 1000 -4257 1022
rect -4191 1000 -4161 1026
rect -4113 1022 -4047 1038
rect -3921 1072 -3855 1088
rect -3921 1038 -3905 1072
rect -3871 1038 -3855 1072
rect -4095 1000 -4065 1022
rect -3999 1000 -3969 1026
rect -3921 1022 -3855 1038
rect -3729 1072 -3663 1088
rect -3729 1038 -3713 1072
rect -3679 1038 -3663 1072
rect -3903 1000 -3873 1022
rect -3807 1000 -3777 1026
rect -3729 1022 -3663 1038
rect -3537 1072 -3471 1088
rect -3537 1038 -3521 1072
rect -3487 1038 -3471 1072
rect -3711 1000 -3681 1022
rect -3615 1000 -3585 1026
rect -3537 1022 -3471 1038
rect -3345 1072 -3279 1088
rect -3345 1038 -3329 1072
rect -3295 1038 -3279 1072
rect -3519 1000 -3489 1022
rect -3423 1000 -3393 1026
rect -3345 1022 -3279 1038
rect -3153 1072 -3087 1088
rect -3153 1038 -3137 1072
rect -3103 1038 -3087 1072
rect -3327 1000 -3297 1022
rect -3231 1000 -3201 1026
rect -3153 1022 -3087 1038
rect -2961 1072 -2895 1088
rect -2961 1038 -2945 1072
rect -2911 1038 -2895 1072
rect -3135 1000 -3105 1022
rect -3039 1000 -3009 1026
rect -2961 1022 -2895 1038
rect -2769 1072 -2703 1088
rect -2769 1038 -2753 1072
rect -2719 1038 -2703 1072
rect -2943 1000 -2913 1022
rect -2847 1000 -2817 1026
rect -2769 1022 -2703 1038
rect -2577 1072 -2511 1088
rect -2577 1038 -2561 1072
rect -2527 1038 -2511 1072
rect -2751 1000 -2721 1022
rect -2655 1000 -2625 1026
rect -2577 1022 -2511 1038
rect -2385 1072 -2319 1088
rect -2385 1038 -2369 1072
rect -2335 1038 -2319 1072
rect -2559 1000 -2529 1022
rect -2463 1000 -2433 1026
rect -2385 1022 -2319 1038
rect -2193 1072 -2127 1088
rect -2193 1038 -2177 1072
rect -2143 1038 -2127 1072
rect -2367 1000 -2337 1022
rect -2271 1000 -2241 1026
rect -2193 1022 -2127 1038
rect -2001 1072 -1935 1088
rect -2001 1038 -1985 1072
rect -1951 1038 -1935 1072
rect -2175 1000 -2145 1022
rect -2079 1000 -2049 1026
rect -2001 1022 -1935 1038
rect -1809 1072 -1743 1088
rect -1809 1038 -1793 1072
rect -1759 1038 -1743 1072
rect -1983 1000 -1953 1022
rect -1887 1000 -1857 1026
rect -1809 1022 -1743 1038
rect -1617 1072 -1551 1088
rect -1617 1038 -1601 1072
rect -1567 1038 -1551 1072
rect -1791 1000 -1761 1022
rect -1695 1000 -1665 1026
rect -1617 1022 -1551 1038
rect -1425 1072 -1359 1088
rect -1425 1038 -1409 1072
rect -1375 1038 -1359 1072
rect -1599 1000 -1569 1022
rect -1503 1000 -1473 1026
rect -1425 1022 -1359 1038
rect -1233 1072 -1167 1088
rect -1233 1038 -1217 1072
rect -1183 1038 -1167 1072
rect -1407 1000 -1377 1022
rect -1311 1000 -1281 1026
rect -1233 1022 -1167 1038
rect -1041 1072 -975 1088
rect -1041 1038 -1025 1072
rect -991 1038 -975 1072
rect -1215 1000 -1185 1022
rect -1119 1000 -1089 1026
rect -1041 1022 -975 1038
rect -849 1072 -783 1088
rect -849 1038 -833 1072
rect -799 1038 -783 1072
rect -1023 1000 -993 1022
rect -927 1000 -897 1026
rect -849 1022 -783 1038
rect -657 1072 -591 1088
rect -657 1038 -641 1072
rect -607 1038 -591 1072
rect -831 1000 -801 1022
rect -735 1000 -705 1026
rect -657 1022 -591 1038
rect -465 1072 -399 1088
rect -465 1038 -449 1072
rect -415 1038 -399 1072
rect -639 1000 -609 1022
rect -543 1000 -513 1026
rect -465 1022 -399 1038
rect -273 1072 -207 1088
rect -273 1038 -257 1072
rect -223 1038 -207 1072
rect -447 1000 -417 1022
rect -351 1000 -321 1026
rect -273 1022 -207 1038
rect -81 1072 -15 1088
rect -81 1038 -65 1072
rect -31 1038 -15 1072
rect -255 1000 -225 1022
rect -159 1000 -129 1026
rect -81 1022 -15 1038
rect 111 1072 177 1088
rect 111 1038 127 1072
rect 161 1038 177 1072
rect -63 1000 -33 1022
rect 33 1000 63 1026
rect 111 1022 177 1038
rect 303 1072 369 1088
rect 303 1038 319 1072
rect 353 1038 369 1072
rect 129 1000 159 1022
rect 225 1000 255 1026
rect 303 1022 369 1038
rect 495 1072 561 1088
rect 495 1038 511 1072
rect 545 1038 561 1072
rect 321 1000 351 1022
rect 417 1000 447 1026
rect 495 1022 561 1038
rect 687 1072 753 1088
rect 687 1038 703 1072
rect 737 1038 753 1072
rect 513 1000 543 1022
rect 609 1000 639 1026
rect 687 1022 753 1038
rect 879 1072 945 1088
rect 879 1038 895 1072
rect 929 1038 945 1072
rect 705 1000 735 1022
rect 801 1000 831 1026
rect 879 1022 945 1038
rect 1071 1072 1137 1088
rect 1071 1038 1087 1072
rect 1121 1038 1137 1072
rect 897 1000 927 1022
rect 993 1000 1023 1026
rect 1071 1022 1137 1038
rect 1263 1072 1329 1088
rect 1263 1038 1279 1072
rect 1313 1038 1329 1072
rect 1089 1000 1119 1022
rect 1185 1000 1215 1026
rect 1263 1022 1329 1038
rect 1455 1072 1521 1088
rect 1455 1038 1471 1072
rect 1505 1038 1521 1072
rect 1281 1000 1311 1022
rect 1377 1000 1407 1026
rect 1455 1022 1521 1038
rect 1647 1072 1713 1088
rect 1647 1038 1663 1072
rect 1697 1038 1713 1072
rect 1473 1000 1503 1022
rect 1569 1000 1599 1026
rect 1647 1022 1713 1038
rect 1839 1072 1905 1088
rect 1839 1038 1855 1072
rect 1889 1038 1905 1072
rect 1665 1000 1695 1022
rect 1761 1000 1791 1026
rect 1839 1022 1905 1038
rect 2031 1072 2097 1088
rect 2031 1038 2047 1072
rect 2081 1038 2097 1072
rect 1857 1000 1887 1022
rect 1953 1000 1983 1026
rect 2031 1022 2097 1038
rect 2223 1072 2289 1088
rect 2223 1038 2239 1072
rect 2273 1038 2289 1072
rect 2049 1000 2079 1022
rect 2145 1000 2175 1026
rect 2223 1022 2289 1038
rect 2415 1072 2481 1088
rect 2415 1038 2431 1072
rect 2465 1038 2481 1072
rect 2241 1000 2271 1022
rect 2337 1000 2367 1026
rect 2415 1022 2481 1038
rect 2607 1072 2673 1088
rect 2607 1038 2623 1072
rect 2657 1038 2673 1072
rect 2433 1000 2463 1022
rect 2529 1000 2559 1026
rect 2607 1022 2673 1038
rect 2799 1072 2865 1088
rect 2799 1038 2815 1072
rect 2849 1038 2865 1072
rect 2625 1000 2655 1022
rect 2721 1000 2751 1026
rect 2799 1022 2865 1038
rect 2991 1072 3057 1088
rect 2991 1038 3007 1072
rect 3041 1038 3057 1072
rect 2817 1000 2847 1022
rect 2913 1000 2943 1026
rect 2991 1022 3057 1038
rect 3183 1072 3249 1088
rect 3183 1038 3199 1072
rect 3233 1038 3249 1072
rect 3009 1000 3039 1022
rect 3105 1000 3135 1026
rect 3183 1022 3249 1038
rect 3375 1072 3441 1088
rect 3375 1038 3391 1072
rect 3425 1038 3441 1072
rect 3201 1000 3231 1022
rect 3297 1000 3327 1026
rect 3375 1022 3441 1038
rect 3567 1072 3633 1088
rect 3567 1038 3583 1072
rect 3617 1038 3633 1072
rect 3393 1000 3423 1022
rect 3489 1000 3519 1026
rect 3567 1022 3633 1038
rect 3759 1072 3825 1088
rect 3759 1038 3775 1072
rect 3809 1038 3825 1072
rect 3585 1000 3615 1022
rect 3681 1000 3711 1026
rect 3759 1022 3825 1038
rect 3951 1072 4017 1088
rect 3951 1038 3967 1072
rect 4001 1038 4017 1072
rect 3777 1000 3807 1022
rect 3873 1000 3903 1026
rect 3951 1022 4017 1038
rect 4143 1072 4209 1088
rect 4143 1038 4159 1072
rect 4193 1038 4209 1072
rect 3969 1000 3999 1022
rect 4065 1000 4095 1026
rect 4143 1022 4209 1038
rect 4335 1072 4401 1088
rect 4335 1038 4351 1072
rect 4385 1038 4401 1072
rect 4161 1000 4191 1022
rect 4257 1000 4287 1026
rect 4335 1022 4401 1038
rect 4527 1072 4593 1088
rect 4527 1038 4543 1072
rect 4577 1038 4593 1072
rect 4353 1000 4383 1022
rect 4449 1000 4479 1026
rect 4527 1022 4593 1038
rect 4719 1072 4785 1088
rect 4719 1038 4735 1072
rect 4769 1038 4785 1072
rect 4545 1000 4575 1022
rect 4641 1000 4671 1026
rect 4719 1022 4785 1038
rect 4737 1000 4767 1022
rect -4767 -1022 -4737 -1000
rect -4785 -1038 -4719 -1022
rect -4671 -1026 -4641 -1000
rect -4575 -1022 -4545 -1000
rect -4785 -1072 -4769 -1038
rect -4735 -1072 -4719 -1038
rect -4785 -1088 -4719 -1072
rect -4593 -1038 -4527 -1022
rect -4479 -1026 -4449 -1000
rect -4383 -1022 -4353 -1000
rect -4593 -1072 -4577 -1038
rect -4543 -1072 -4527 -1038
rect -4593 -1088 -4527 -1072
rect -4401 -1038 -4335 -1022
rect -4287 -1026 -4257 -1000
rect -4191 -1022 -4161 -1000
rect -4401 -1072 -4385 -1038
rect -4351 -1072 -4335 -1038
rect -4401 -1088 -4335 -1072
rect -4209 -1038 -4143 -1022
rect -4095 -1026 -4065 -1000
rect -3999 -1022 -3969 -1000
rect -4209 -1072 -4193 -1038
rect -4159 -1072 -4143 -1038
rect -4209 -1088 -4143 -1072
rect -4017 -1038 -3951 -1022
rect -3903 -1026 -3873 -1000
rect -3807 -1022 -3777 -1000
rect -4017 -1072 -4001 -1038
rect -3967 -1072 -3951 -1038
rect -4017 -1088 -3951 -1072
rect -3825 -1038 -3759 -1022
rect -3711 -1026 -3681 -1000
rect -3615 -1022 -3585 -1000
rect -3825 -1072 -3809 -1038
rect -3775 -1072 -3759 -1038
rect -3825 -1088 -3759 -1072
rect -3633 -1038 -3567 -1022
rect -3519 -1026 -3489 -1000
rect -3423 -1022 -3393 -1000
rect -3633 -1072 -3617 -1038
rect -3583 -1072 -3567 -1038
rect -3633 -1088 -3567 -1072
rect -3441 -1038 -3375 -1022
rect -3327 -1026 -3297 -1000
rect -3231 -1022 -3201 -1000
rect -3441 -1072 -3425 -1038
rect -3391 -1072 -3375 -1038
rect -3441 -1088 -3375 -1072
rect -3249 -1038 -3183 -1022
rect -3135 -1026 -3105 -1000
rect -3039 -1022 -3009 -1000
rect -3249 -1072 -3233 -1038
rect -3199 -1072 -3183 -1038
rect -3249 -1088 -3183 -1072
rect -3057 -1038 -2991 -1022
rect -2943 -1026 -2913 -1000
rect -2847 -1022 -2817 -1000
rect -3057 -1072 -3041 -1038
rect -3007 -1072 -2991 -1038
rect -3057 -1088 -2991 -1072
rect -2865 -1038 -2799 -1022
rect -2751 -1026 -2721 -1000
rect -2655 -1022 -2625 -1000
rect -2865 -1072 -2849 -1038
rect -2815 -1072 -2799 -1038
rect -2865 -1088 -2799 -1072
rect -2673 -1038 -2607 -1022
rect -2559 -1026 -2529 -1000
rect -2463 -1022 -2433 -1000
rect -2673 -1072 -2657 -1038
rect -2623 -1072 -2607 -1038
rect -2673 -1088 -2607 -1072
rect -2481 -1038 -2415 -1022
rect -2367 -1026 -2337 -1000
rect -2271 -1022 -2241 -1000
rect -2481 -1072 -2465 -1038
rect -2431 -1072 -2415 -1038
rect -2481 -1088 -2415 -1072
rect -2289 -1038 -2223 -1022
rect -2175 -1026 -2145 -1000
rect -2079 -1022 -2049 -1000
rect -2289 -1072 -2273 -1038
rect -2239 -1072 -2223 -1038
rect -2289 -1088 -2223 -1072
rect -2097 -1038 -2031 -1022
rect -1983 -1026 -1953 -1000
rect -1887 -1022 -1857 -1000
rect -2097 -1072 -2081 -1038
rect -2047 -1072 -2031 -1038
rect -2097 -1088 -2031 -1072
rect -1905 -1038 -1839 -1022
rect -1791 -1026 -1761 -1000
rect -1695 -1022 -1665 -1000
rect -1905 -1072 -1889 -1038
rect -1855 -1072 -1839 -1038
rect -1905 -1088 -1839 -1072
rect -1713 -1038 -1647 -1022
rect -1599 -1026 -1569 -1000
rect -1503 -1022 -1473 -1000
rect -1713 -1072 -1697 -1038
rect -1663 -1072 -1647 -1038
rect -1713 -1088 -1647 -1072
rect -1521 -1038 -1455 -1022
rect -1407 -1026 -1377 -1000
rect -1311 -1022 -1281 -1000
rect -1521 -1072 -1505 -1038
rect -1471 -1072 -1455 -1038
rect -1521 -1088 -1455 -1072
rect -1329 -1038 -1263 -1022
rect -1215 -1026 -1185 -1000
rect -1119 -1022 -1089 -1000
rect -1329 -1072 -1313 -1038
rect -1279 -1072 -1263 -1038
rect -1329 -1088 -1263 -1072
rect -1137 -1038 -1071 -1022
rect -1023 -1026 -993 -1000
rect -927 -1022 -897 -1000
rect -1137 -1072 -1121 -1038
rect -1087 -1072 -1071 -1038
rect -1137 -1088 -1071 -1072
rect -945 -1038 -879 -1022
rect -831 -1026 -801 -1000
rect -735 -1022 -705 -1000
rect -945 -1072 -929 -1038
rect -895 -1072 -879 -1038
rect -945 -1088 -879 -1072
rect -753 -1038 -687 -1022
rect -639 -1026 -609 -1000
rect -543 -1022 -513 -1000
rect -753 -1072 -737 -1038
rect -703 -1072 -687 -1038
rect -753 -1088 -687 -1072
rect -561 -1038 -495 -1022
rect -447 -1026 -417 -1000
rect -351 -1022 -321 -1000
rect -561 -1072 -545 -1038
rect -511 -1072 -495 -1038
rect -561 -1088 -495 -1072
rect -369 -1038 -303 -1022
rect -255 -1026 -225 -1000
rect -159 -1022 -129 -1000
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -369 -1088 -303 -1072
rect -177 -1038 -111 -1022
rect -63 -1026 -33 -1000
rect 33 -1022 63 -1000
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect -177 -1088 -111 -1072
rect 15 -1038 81 -1022
rect 129 -1026 159 -1000
rect 225 -1022 255 -1000
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 15 -1088 81 -1072
rect 207 -1038 273 -1022
rect 321 -1026 351 -1000
rect 417 -1022 447 -1000
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect 207 -1088 273 -1072
rect 399 -1038 465 -1022
rect 513 -1026 543 -1000
rect 609 -1022 639 -1000
rect 399 -1072 415 -1038
rect 449 -1072 465 -1038
rect 399 -1088 465 -1072
rect 591 -1038 657 -1022
rect 705 -1026 735 -1000
rect 801 -1022 831 -1000
rect 591 -1072 607 -1038
rect 641 -1072 657 -1038
rect 591 -1088 657 -1072
rect 783 -1038 849 -1022
rect 897 -1026 927 -1000
rect 993 -1022 1023 -1000
rect 783 -1072 799 -1038
rect 833 -1072 849 -1038
rect 783 -1088 849 -1072
rect 975 -1038 1041 -1022
rect 1089 -1026 1119 -1000
rect 1185 -1022 1215 -1000
rect 975 -1072 991 -1038
rect 1025 -1072 1041 -1038
rect 975 -1088 1041 -1072
rect 1167 -1038 1233 -1022
rect 1281 -1026 1311 -1000
rect 1377 -1022 1407 -1000
rect 1167 -1072 1183 -1038
rect 1217 -1072 1233 -1038
rect 1167 -1088 1233 -1072
rect 1359 -1038 1425 -1022
rect 1473 -1026 1503 -1000
rect 1569 -1022 1599 -1000
rect 1359 -1072 1375 -1038
rect 1409 -1072 1425 -1038
rect 1359 -1088 1425 -1072
rect 1551 -1038 1617 -1022
rect 1665 -1026 1695 -1000
rect 1761 -1022 1791 -1000
rect 1551 -1072 1567 -1038
rect 1601 -1072 1617 -1038
rect 1551 -1088 1617 -1072
rect 1743 -1038 1809 -1022
rect 1857 -1026 1887 -1000
rect 1953 -1022 1983 -1000
rect 1743 -1072 1759 -1038
rect 1793 -1072 1809 -1038
rect 1743 -1088 1809 -1072
rect 1935 -1038 2001 -1022
rect 2049 -1026 2079 -1000
rect 2145 -1022 2175 -1000
rect 1935 -1072 1951 -1038
rect 1985 -1072 2001 -1038
rect 1935 -1088 2001 -1072
rect 2127 -1038 2193 -1022
rect 2241 -1026 2271 -1000
rect 2337 -1022 2367 -1000
rect 2127 -1072 2143 -1038
rect 2177 -1072 2193 -1038
rect 2127 -1088 2193 -1072
rect 2319 -1038 2385 -1022
rect 2433 -1026 2463 -1000
rect 2529 -1022 2559 -1000
rect 2319 -1072 2335 -1038
rect 2369 -1072 2385 -1038
rect 2319 -1088 2385 -1072
rect 2511 -1038 2577 -1022
rect 2625 -1026 2655 -1000
rect 2721 -1022 2751 -1000
rect 2511 -1072 2527 -1038
rect 2561 -1072 2577 -1038
rect 2511 -1088 2577 -1072
rect 2703 -1038 2769 -1022
rect 2817 -1026 2847 -1000
rect 2913 -1022 2943 -1000
rect 2703 -1072 2719 -1038
rect 2753 -1072 2769 -1038
rect 2703 -1088 2769 -1072
rect 2895 -1038 2961 -1022
rect 3009 -1026 3039 -1000
rect 3105 -1022 3135 -1000
rect 2895 -1072 2911 -1038
rect 2945 -1072 2961 -1038
rect 2895 -1088 2961 -1072
rect 3087 -1038 3153 -1022
rect 3201 -1026 3231 -1000
rect 3297 -1022 3327 -1000
rect 3087 -1072 3103 -1038
rect 3137 -1072 3153 -1038
rect 3087 -1088 3153 -1072
rect 3279 -1038 3345 -1022
rect 3393 -1026 3423 -1000
rect 3489 -1022 3519 -1000
rect 3279 -1072 3295 -1038
rect 3329 -1072 3345 -1038
rect 3279 -1088 3345 -1072
rect 3471 -1038 3537 -1022
rect 3585 -1026 3615 -1000
rect 3681 -1022 3711 -1000
rect 3471 -1072 3487 -1038
rect 3521 -1072 3537 -1038
rect 3471 -1088 3537 -1072
rect 3663 -1038 3729 -1022
rect 3777 -1026 3807 -1000
rect 3873 -1022 3903 -1000
rect 3663 -1072 3679 -1038
rect 3713 -1072 3729 -1038
rect 3663 -1088 3729 -1072
rect 3855 -1038 3921 -1022
rect 3969 -1026 3999 -1000
rect 4065 -1022 4095 -1000
rect 3855 -1072 3871 -1038
rect 3905 -1072 3921 -1038
rect 3855 -1088 3921 -1072
rect 4047 -1038 4113 -1022
rect 4161 -1026 4191 -1000
rect 4257 -1022 4287 -1000
rect 4047 -1072 4063 -1038
rect 4097 -1072 4113 -1038
rect 4047 -1088 4113 -1072
rect 4239 -1038 4305 -1022
rect 4353 -1026 4383 -1000
rect 4449 -1022 4479 -1000
rect 4239 -1072 4255 -1038
rect 4289 -1072 4305 -1038
rect 4239 -1088 4305 -1072
rect 4431 -1038 4497 -1022
rect 4545 -1026 4575 -1000
rect 4641 -1022 4671 -1000
rect 4431 -1072 4447 -1038
rect 4481 -1072 4497 -1038
rect 4431 -1088 4497 -1072
rect 4623 -1038 4689 -1022
rect 4737 -1026 4767 -1000
rect 4623 -1072 4639 -1038
rect 4673 -1072 4689 -1038
rect 4623 -1088 4689 -1072
<< polycont >>
rect -4673 1038 -4639 1072
rect -4481 1038 -4447 1072
rect -4289 1038 -4255 1072
rect -4097 1038 -4063 1072
rect -3905 1038 -3871 1072
rect -3713 1038 -3679 1072
rect -3521 1038 -3487 1072
rect -3329 1038 -3295 1072
rect -3137 1038 -3103 1072
rect -2945 1038 -2911 1072
rect -2753 1038 -2719 1072
rect -2561 1038 -2527 1072
rect -2369 1038 -2335 1072
rect -2177 1038 -2143 1072
rect -1985 1038 -1951 1072
rect -1793 1038 -1759 1072
rect -1601 1038 -1567 1072
rect -1409 1038 -1375 1072
rect -1217 1038 -1183 1072
rect -1025 1038 -991 1072
rect -833 1038 -799 1072
rect -641 1038 -607 1072
rect -449 1038 -415 1072
rect -257 1038 -223 1072
rect -65 1038 -31 1072
rect 127 1038 161 1072
rect 319 1038 353 1072
rect 511 1038 545 1072
rect 703 1038 737 1072
rect 895 1038 929 1072
rect 1087 1038 1121 1072
rect 1279 1038 1313 1072
rect 1471 1038 1505 1072
rect 1663 1038 1697 1072
rect 1855 1038 1889 1072
rect 2047 1038 2081 1072
rect 2239 1038 2273 1072
rect 2431 1038 2465 1072
rect 2623 1038 2657 1072
rect 2815 1038 2849 1072
rect 3007 1038 3041 1072
rect 3199 1038 3233 1072
rect 3391 1038 3425 1072
rect 3583 1038 3617 1072
rect 3775 1038 3809 1072
rect 3967 1038 4001 1072
rect 4159 1038 4193 1072
rect 4351 1038 4385 1072
rect 4543 1038 4577 1072
rect 4735 1038 4769 1072
rect -4769 -1072 -4735 -1038
rect -4577 -1072 -4543 -1038
rect -4385 -1072 -4351 -1038
rect -4193 -1072 -4159 -1038
rect -4001 -1072 -3967 -1038
rect -3809 -1072 -3775 -1038
rect -3617 -1072 -3583 -1038
rect -3425 -1072 -3391 -1038
rect -3233 -1072 -3199 -1038
rect -3041 -1072 -3007 -1038
rect -2849 -1072 -2815 -1038
rect -2657 -1072 -2623 -1038
rect -2465 -1072 -2431 -1038
rect -2273 -1072 -2239 -1038
rect -2081 -1072 -2047 -1038
rect -1889 -1072 -1855 -1038
rect -1697 -1072 -1663 -1038
rect -1505 -1072 -1471 -1038
rect -1313 -1072 -1279 -1038
rect -1121 -1072 -1087 -1038
rect -929 -1072 -895 -1038
rect -737 -1072 -703 -1038
rect -545 -1072 -511 -1038
rect -353 -1072 -319 -1038
rect -161 -1072 -127 -1038
rect 31 -1072 65 -1038
rect 223 -1072 257 -1038
rect 415 -1072 449 -1038
rect 607 -1072 641 -1038
rect 799 -1072 833 -1038
rect 991 -1072 1025 -1038
rect 1183 -1072 1217 -1038
rect 1375 -1072 1409 -1038
rect 1567 -1072 1601 -1038
rect 1759 -1072 1793 -1038
rect 1951 -1072 1985 -1038
rect 2143 -1072 2177 -1038
rect 2335 -1072 2369 -1038
rect 2527 -1072 2561 -1038
rect 2719 -1072 2753 -1038
rect 2911 -1072 2945 -1038
rect 3103 -1072 3137 -1038
rect 3295 -1072 3329 -1038
rect 3487 -1072 3521 -1038
rect 3679 -1072 3713 -1038
rect 3871 -1072 3905 -1038
rect 4063 -1072 4097 -1038
rect 4255 -1072 4289 -1038
rect 4447 -1072 4481 -1038
rect 4639 -1072 4673 -1038
<< locali >>
rect -4931 1140 -4811 1174
rect -4777 1140 -4743 1174
rect -4709 1140 -4675 1174
rect -4641 1140 -4607 1174
rect -4573 1140 -4539 1174
rect -4505 1140 -4471 1174
rect -4437 1140 -4403 1174
rect -4369 1140 -4335 1174
rect -4301 1140 -4267 1174
rect -4233 1140 -4199 1174
rect -4165 1140 -4131 1174
rect -4097 1140 -4063 1174
rect -4029 1140 -3995 1174
rect -3961 1140 -3927 1174
rect -3893 1140 -3859 1174
rect -3825 1140 -3791 1174
rect -3757 1140 -3723 1174
rect -3689 1140 -3655 1174
rect -3621 1140 -3587 1174
rect -3553 1140 -3519 1174
rect -3485 1140 -3451 1174
rect -3417 1140 -3383 1174
rect -3349 1140 -3315 1174
rect -3281 1140 -3247 1174
rect -3213 1140 -3179 1174
rect -3145 1140 -3111 1174
rect -3077 1140 -3043 1174
rect -3009 1140 -2975 1174
rect -2941 1140 -2907 1174
rect -2873 1140 -2839 1174
rect -2805 1140 -2771 1174
rect -2737 1140 -2703 1174
rect -2669 1140 -2635 1174
rect -2601 1140 -2567 1174
rect -2533 1140 -2499 1174
rect -2465 1140 -2431 1174
rect -2397 1140 -2363 1174
rect -2329 1140 -2295 1174
rect -2261 1140 -2227 1174
rect -2193 1140 -2159 1174
rect -2125 1140 -2091 1174
rect -2057 1140 -2023 1174
rect -1989 1140 -1955 1174
rect -1921 1140 -1887 1174
rect -1853 1140 -1819 1174
rect -1785 1140 -1751 1174
rect -1717 1140 -1683 1174
rect -1649 1140 -1615 1174
rect -1581 1140 -1547 1174
rect -1513 1140 -1479 1174
rect -1445 1140 -1411 1174
rect -1377 1140 -1343 1174
rect -1309 1140 -1275 1174
rect -1241 1140 -1207 1174
rect -1173 1140 -1139 1174
rect -1105 1140 -1071 1174
rect -1037 1140 -1003 1174
rect -969 1140 -935 1174
rect -901 1140 -867 1174
rect -833 1140 -799 1174
rect -765 1140 -731 1174
rect -697 1140 -663 1174
rect -629 1140 -595 1174
rect -561 1140 -527 1174
rect -493 1140 -459 1174
rect -425 1140 -391 1174
rect -357 1140 -323 1174
rect -289 1140 -255 1174
rect -221 1140 -187 1174
rect -153 1140 -119 1174
rect -85 1140 -51 1174
rect -17 1140 17 1174
rect 51 1140 85 1174
rect 119 1140 153 1174
rect 187 1140 221 1174
rect 255 1140 289 1174
rect 323 1140 357 1174
rect 391 1140 425 1174
rect 459 1140 493 1174
rect 527 1140 561 1174
rect 595 1140 629 1174
rect 663 1140 697 1174
rect 731 1140 765 1174
rect 799 1140 833 1174
rect 867 1140 901 1174
rect 935 1140 969 1174
rect 1003 1140 1037 1174
rect 1071 1140 1105 1174
rect 1139 1140 1173 1174
rect 1207 1140 1241 1174
rect 1275 1140 1309 1174
rect 1343 1140 1377 1174
rect 1411 1140 1445 1174
rect 1479 1140 1513 1174
rect 1547 1140 1581 1174
rect 1615 1140 1649 1174
rect 1683 1140 1717 1174
rect 1751 1140 1785 1174
rect 1819 1140 1853 1174
rect 1887 1140 1921 1174
rect 1955 1140 1989 1174
rect 2023 1140 2057 1174
rect 2091 1140 2125 1174
rect 2159 1140 2193 1174
rect 2227 1140 2261 1174
rect 2295 1140 2329 1174
rect 2363 1140 2397 1174
rect 2431 1140 2465 1174
rect 2499 1140 2533 1174
rect 2567 1140 2601 1174
rect 2635 1140 2669 1174
rect 2703 1140 2737 1174
rect 2771 1140 2805 1174
rect 2839 1140 2873 1174
rect 2907 1140 2941 1174
rect 2975 1140 3009 1174
rect 3043 1140 3077 1174
rect 3111 1140 3145 1174
rect 3179 1140 3213 1174
rect 3247 1140 3281 1174
rect 3315 1140 3349 1174
rect 3383 1140 3417 1174
rect 3451 1140 3485 1174
rect 3519 1140 3553 1174
rect 3587 1140 3621 1174
rect 3655 1140 3689 1174
rect 3723 1140 3757 1174
rect 3791 1140 3825 1174
rect 3859 1140 3893 1174
rect 3927 1140 3961 1174
rect 3995 1140 4029 1174
rect 4063 1140 4097 1174
rect 4131 1140 4165 1174
rect 4199 1140 4233 1174
rect 4267 1140 4301 1174
rect 4335 1140 4369 1174
rect 4403 1140 4437 1174
rect 4471 1140 4505 1174
rect 4539 1140 4573 1174
rect 4607 1140 4641 1174
rect 4675 1140 4709 1174
rect 4743 1140 4777 1174
rect 4811 1140 4931 1174
rect -4931 1071 -4897 1140
rect -4689 1038 -4673 1072
rect -4639 1038 -4623 1072
rect -4497 1038 -4481 1072
rect -4447 1038 -4431 1072
rect -4305 1038 -4289 1072
rect -4255 1038 -4239 1072
rect -4113 1038 -4097 1072
rect -4063 1038 -4047 1072
rect -3921 1038 -3905 1072
rect -3871 1038 -3855 1072
rect -3729 1038 -3713 1072
rect -3679 1038 -3663 1072
rect -3537 1038 -3521 1072
rect -3487 1038 -3471 1072
rect -3345 1038 -3329 1072
rect -3295 1038 -3279 1072
rect -3153 1038 -3137 1072
rect -3103 1038 -3087 1072
rect -2961 1038 -2945 1072
rect -2911 1038 -2895 1072
rect -2769 1038 -2753 1072
rect -2719 1038 -2703 1072
rect -2577 1038 -2561 1072
rect -2527 1038 -2511 1072
rect -2385 1038 -2369 1072
rect -2335 1038 -2319 1072
rect -2193 1038 -2177 1072
rect -2143 1038 -2127 1072
rect -2001 1038 -1985 1072
rect -1951 1038 -1935 1072
rect -1809 1038 -1793 1072
rect -1759 1038 -1743 1072
rect -1617 1038 -1601 1072
rect -1567 1038 -1551 1072
rect -1425 1038 -1409 1072
rect -1375 1038 -1359 1072
rect -1233 1038 -1217 1072
rect -1183 1038 -1167 1072
rect -1041 1038 -1025 1072
rect -991 1038 -975 1072
rect -849 1038 -833 1072
rect -799 1038 -783 1072
rect -657 1038 -641 1072
rect -607 1038 -591 1072
rect -465 1038 -449 1072
rect -415 1038 -399 1072
rect -273 1038 -257 1072
rect -223 1038 -207 1072
rect -81 1038 -65 1072
rect -31 1038 -15 1072
rect 111 1038 127 1072
rect 161 1038 177 1072
rect 303 1038 319 1072
rect 353 1038 369 1072
rect 495 1038 511 1072
rect 545 1038 561 1072
rect 687 1038 703 1072
rect 737 1038 753 1072
rect 879 1038 895 1072
rect 929 1038 945 1072
rect 1071 1038 1087 1072
rect 1121 1038 1137 1072
rect 1263 1038 1279 1072
rect 1313 1038 1329 1072
rect 1455 1038 1471 1072
rect 1505 1038 1521 1072
rect 1647 1038 1663 1072
rect 1697 1038 1713 1072
rect 1839 1038 1855 1072
rect 1889 1038 1905 1072
rect 2031 1038 2047 1072
rect 2081 1038 2097 1072
rect 2223 1038 2239 1072
rect 2273 1038 2289 1072
rect 2415 1038 2431 1072
rect 2465 1038 2481 1072
rect 2607 1038 2623 1072
rect 2657 1038 2673 1072
rect 2799 1038 2815 1072
rect 2849 1038 2865 1072
rect 2991 1038 3007 1072
rect 3041 1038 3057 1072
rect 3183 1038 3199 1072
rect 3233 1038 3249 1072
rect 3375 1038 3391 1072
rect 3425 1038 3441 1072
rect 3567 1038 3583 1072
rect 3617 1038 3633 1072
rect 3759 1038 3775 1072
rect 3809 1038 3825 1072
rect 3951 1038 3967 1072
rect 4001 1038 4017 1072
rect 4143 1038 4159 1072
rect 4193 1038 4209 1072
rect 4335 1038 4351 1072
rect 4385 1038 4401 1072
rect 4527 1038 4543 1072
rect 4577 1038 4593 1072
rect 4719 1038 4735 1072
rect 4769 1038 4785 1072
rect 4897 1071 4931 1140
rect -4931 1003 -4897 1037
rect -4931 935 -4897 969
rect -4931 867 -4897 901
rect -4931 799 -4897 833
rect -4931 731 -4897 765
rect -4931 663 -4897 697
rect -4931 595 -4897 629
rect -4931 527 -4897 561
rect -4931 459 -4897 493
rect -4931 391 -4897 425
rect -4931 323 -4897 357
rect -4931 255 -4897 289
rect -4931 187 -4897 221
rect -4931 119 -4897 153
rect -4931 51 -4897 85
rect -4931 -17 -4897 17
rect -4931 -85 -4897 -51
rect -4931 -153 -4897 -119
rect -4931 -221 -4897 -187
rect -4931 -289 -4897 -255
rect -4931 -357 -4897 -323
rect -4931 -425 -4897 -391
rect -4931 -493 -4897 -459
rect -4931 -561 -4897 -527
rect -4931 -629 -4897 -595
rect -4931 -697 -4897 -663
rect -4931 -765 -4897 -731
rect -4931 -833 -4897 -799
rect -4931 -901 -4897 -867
rect -4931 -969 -4897 -935
rect -4931 -1037 -4897 -1003
rect -4817 969 -4783 1004
rect -4817 901 -4783 935
rect -4817 833 -4783 867
rect -4817 765 -4783 799
rect -4817 697 -4783 731
rect -4817 629 -4783 663
rect -4817 561 -4783 595
rect -4817 493 -4783 527
rect -4817 425 -4783 459
rect -4817 357 -4783 391
rect -4817 289 -4783 323
rect -4817 221 -4783 255
rect -4817 153 -4783 187
rect -4817 85 -4783 119
rect -4817 17 -4783 51
rect -4817 -51 -4783 -17
rect -4817 -119 -4783 -85
rect -4817 -187 -4783 -153
rect -4817 -255 -4783 -221
rect -4817 -323 -4783 -289
rect -4817 -391 -4783 -357
rect -4817 -459 -4783 -425
rect -4817 -527 -4783 -493
rect -4817 -595 -4783 -561
rect -4817 -663 -4783 -629
rect -4817 -731 -4783 -697
rect -4817 -799 -4783 -765
rect -4817 -867 -4783 -833
rect -4817 -935 -4783 -901
rect -4817 -1004 -4783 -969
rect -4721 969 -4687 1004
rect -4721 901 -4687 935
rect -4721 833 -4687 867
rect -4721 765 -4687 799
rect -4721 697 -4687 731
rect -4721 629 -4687 663
rect -4721 561 -4687 595
rect -4721 493 -4687 527
rect -4721 425 -4687 459
rect -4721 357 -4687 391
rect -4721 289 -4687 323
rect -4721 221 -4687 255
rect -4721 153 -4687 187
rect -4721 85 -4687 119
rect -4721 17 -4687 51
rect -4721 -51 -4687 -17
rect -4721 -119 -4687 -85
rect -4721 -187 -4687 -153
rect -4721 -255 -4687 -221
rect -4721 -323 -4687 -289
rect -4721 -391 -4687 -357
rect -4721 -459 -4687 -425
rect -4721 -527 -4687 -493
rect -4721 -595 -4687 -561
rect -4721 -663 -4687 -629
rect -4721 -731 -4687 -697
rect -4721 -799 -4687 -765
rect -4721 -867 -4687 -833
rect -4721 -935 -4687 -901
rect -4721 -1004 -4687 -969
rect -4625 969 -4591 1004
rect -4625 901 -4591 935
rect -4625 833 -4591 867
rect -4625 765 -4591 799
rect -4625 697 -4591 731
rect -4625 629 -4591 663
rect -4625 561 -4591 595
rect -4625 493 -4591 527
rect -4625 425 -4591 459
rect -4625 357 -4591 391
rect -4625 289 -4591 323
rect -4625 221 -4591 255
rect -4625 153 -4591 187
rect -4625 85 -4591 119
rect -4625 17 -4591 51
rect -4625 -51 -4591 -17
rect -4625 -119 -4591 -85
rect -4625 -187 -4591 -153
rect -4625 -255 -4591 -221
rect -4625 -323 -4591 -289
rect -4625 -391 -4591 -357
rect -4625 -459 -4591 -425
rect -4625 -527 -4591 -493
rect -4625 -595 -4591 -561
rect -4625 -663 -4591 -629
rect -4625 -731 -4591 -697
rect -4625 -799 -4591 -765
rect -4625 -867 -4591 -833
rect -4625 -935 -4591 -901
rect -4625 -1004 -4591 -969
rect -4529 969 -4495 1004
rect -4529 901 -4495 935
rect -4529 833 -4495 867
rect -4529 765 -4495 799
rect -4529 697 -4495 731
rect -4529 629 -4495 663
rect -4529 561 -4495 595
rect -4529 493 -4495 527
rect -4529 425 -4495 459
rect -4529 357 -4495 391
rect -4529 289 -4495 323
rect -4529 221 -4495 255
rect -4529 153 -4495 187
rect -4529 85 -4495 119
rect -4529 17 -4495 51
rect -4529 -51 -4495 -17
rect -4529 -119 -4495 -85
rect -4529 -187 -4495 -153
rect -4529 -255 -4495 -221
rect -4529 -323 -4495 -289
rect -4529 -391 -4495 -357
rect -4529 -459 -4495 -425
rect -4529 -527 -4495 -493
rect -4529 -595 -4495 -561
rect -4529 -663 -4495 -629
rect -4529 -731 -4495 -697
rect -4529 -799 -4495 -765
rect -4529 -867 -4495 -833
rect -4529 -935 -4495 -901
rect -4529 -1004 -4495 -969
rect -4433 969 -4399 1004
rect -4433 901 -4399 935
rect -4433 833 -4399 867
rect -4433 765 -4399 799
rect -4433 697 -4399 731
rect -4433 629 -4399 663
rect -4433 561 -4399 595
rect -4433 493 -4399 527
rect -4433 425 -4399 459
rect -4433 357 -4399 391
rect -4433 289 -4399 323
rect -4433 221 -4399 255
rect -4433 153 -4399 187
rect -4433 85 -4399 119
rect -4433 17 -4399 51
rect -4433 -51 -4399 -17
rect -4433 -119 -4399 -85
rect -4433 -187 -4399 -153
rect -4433 -255 -4399 -221
rect -4433 -323 -4399 -289
rect -4433 -391 -4399 -357
rect -4433 -459 -4399 -425
rect -4433 -527 -4399 -493
rect -4433 -595 -4399 -561
rect -4433 -663 -4399 -629
rect -4433 -731 -4399 -697
rect -4433 -799 -4399 -765
rect -4433 -867 -4399 -833
rect -4433 -935 -4399 -901
rect -4433 -1004 -4399 -969
rect -4337 969 -4303 1004
rect -4337 901 -4303 935
rect -4337 833 -4303 867
rect -4337 765 -4303 799
rect -4337 697 -4303 731
rect -4337 629 -4303 663
rect -4337 561 -4303 595
rect -4337 493 -4303 527
rect -4337 425 -4303 459
rect -4337 357 -4303 391
rect -4337 289 -4303 323
rect -4337 221 -4303 255
rect -4337 153 -4303 187
rect -4337 85 -4303 119
rect -4337 17 -4303 51
rect -4337 -51 -4303 -17
rect -4337 -119 -4303 -85
rect -4337 -187 -4303 -153
rect -4337 -255 -4303 -221
rect -4337 -323 -4303 -289
rect -4337 -391 -4303 -357
rect -4337 -459 -4303 -425
rect -4337 -527 -4303 -493
rect -4337 -595 -4303 -561
rect -4337 -663 -4303 -629
rect -4337 -731 -4303 -697
rect -4337 -799 -4303 -765
rect -4337 -867 -4303 -833
rect -4337 -935 -4303 -901
rect -4337 -1004 -4303 -969
rect -4241 969 -4207 1004
rect -4241 901 -4207 935
rect -4241 833 -4207 867
rect -4241 765 -4207 799
rect -4241 697 -4207 731
rect -4241 629 -4207 663
rect -4241 561 -4207 595
rect -4241 493 -4207 527
rect -4241 425 -4207 459
rect -4241 357 -4207 391
rect -4241 289 -4207 323
rect -4241 221 -4207 255
rect -4241 153 -4207 187
rect -4241 85 -4207 119
rect -4241 17 -4207 51
rect -4241 -51 -4207 -17
rect -4241 -119 -4207 -85
rect -4241 -187 -4207 -153
rect -4241 -255 -4207 -221
rect -4241 -323 -4207 -289
rect -4241 -391 -4207 -357
rect -4241 -459 -4207 -425
rect -4241 -527 -4207 -493
rect -4241 -595 -4207 -561
rect -4241 -663 -4207 -629
rect -4241 -731 -4207 -697
rect -4241 -799 -4207 -765
rect -4241 -867 -4207 -833
rect -4241 -935 -4207 -901
rect -4241 -1004 -4207 -969
rect -4145 969 -4111 1004
rect -4145 901 -4111 935
rect -4145 833 -4111 867
rect -4145 765 -4111 799
rect -4145 697 -4111 731
rect -4145 629 -4111 663
rect -4145 561 -4111 595
rect -4145 493 -4111 527
rect -4145 425 -4111 459
rect -4145 357 -4111 391
rect -4145 289 -4111 323
rect -4145 221 -4111 255
rect -4145 153 -4111 187
rect -4145 85 -4111 119
rect -4145 17 -4111 51
rect -4145 -51 -4111 -17
rect -4145 -119 -4111 -85
rect -4145 -187 -4111 -153
rect -4145 -255 -4111 -221
rect -4145 -323 -4111 -289
rect -4145 -391 -4111 -357
rect -4145 -459 -4111 -425
rect -4145 -527 -4111 -493
rect -4145 -595 -4111 -561
rect -4145 -663 -4111 -629
rect -4145 -731 -4111 -697
rect -4145 -799 -4111 -765
rect -4145 -867 -4111 -833
rect -4145 -935 -4111 -901
rect -4145 -1004 -4111 -969
rect -4049 969 -4015 1004
rect -4049 901 -4015 935
rect -4049 833 -4015 867
rect -4049 765 -4015 799
rect -4049 697 -4015 731
rect -4049 629 -4015 663
rect -4049 561 -4015 595
rect -4049 493 -4015 527
rect -4049 425 -4015 459
rect -4049 357 -4015 391
rect -4049 289 -4015 323
rect -4049 221 -4015 255
rect -4049 153 -4015 187
rect -4049 85 -4015 119
rect -4049 17 -4015 51
rect -4049 -51 -4015 -17
rect -4049 -119 -4015 -85
rect -4049 -187 -4015 -153
rect -4049 -255 -4015 -221
rect -4049 -323 -4015 -289
rect -4049 -391 -4015 -357
rect -4049 -459 -4015 -425
rect -4049 -527 -4015 -493
rect -4049 -595 -4015 -561
rect -4049 -663 -4015 -629
rect -4049 -731 -4015 -697
rect -4049 -799 -4015 -765
rect -4049 -867 -4015 -833
rect -4049 -935 -4015 -901
rect -4049 -1004 -4015 -969
rect -3953 969 -3919 1004
rect -3953 901 -3919 935
rect -3953 833 -3919 867
rect -3953 765 -3919 799
rect -3953 697 -3919 731
rect -3953 629 -3919 663
rect -3953 561 -3919 595
rect -3953 493 -3919 527
rect -3953 425 -3919 459
rect -3953 357 -3919 391
rect -3953 289 -3919 323
rect -3953 221 -3919 255
rect -3953 153 -3919 187
rect -3953 85 -3919 119
rect -3953 17 -3919 51
rect -3953 -51 -3919 -17
rect -3953 -119 -3919 -85
rect -3953 -187 -3919 -153
rect -3953 -255 -3919 -221
rect -3953 -323 -3919 -289
rect -3953 -391 -3919 -357
rect -3953 -459 -3919 -425
rect -3953 -527 -3919 -493
rect -3953 -595 -3919 -561
rect -3953 -663 -3919 -629
rect -3953 -731 -3919 -697
rect -3953 -799 -3919 -765
rect -3953 -867 -3919 -833
rect -3953 -935 -3919 -901
rect -3953 -1004 -3919 -969
rect -3857 969 -3823 1004
rect -3857 901 -3823 935
rect -3857 833 -3823 867
rect -3857 765 -3823 799
rect -3857 697 -3823 731
rect -3857 629 -3823 663
rect -3857 561 -3823 595
rect -3857 493 -3823 527
rect -3857 425 -3823 459
rect -3857 357 -3823 391
rect -3857 289 -3823 323
rect -3857 221 -3823 255
rect -3857 153 -3823 187
rect -3857 85 -3823 119
rect -3857 17 -3823 51
rect -3857 -51 -3823 -17
rect -3857 -119 -3823 -85
rect -3857 -187 -3823 -153
rect -3857 -255 -3823 -221
rect -3857 -323 -3823 -289
rect -3857 -391 -3823 -357
rect -3857 -459 -3823 -425
rect -3857 -527 -3823 -493
rect -3857 -595 -3823 -561
rect -3857 -663 -3823 -629
rect -3857 -731 -3823 -697
rect -3857 -799 -3823 -765
rect -3857 -867 -3823 -833
rect -3857 -935 -3823 -901
rect -3857 -1004 -3823 -969
rect -3761 969 -3727 1004
rect -3761 901 -3727 935
rect -3761 833 -3727 867
rect -3761 765 -3727 799
rect -3761 697 -3727 731
rect -3761 629 -3727 663
rect -3761 561 -3727 595
rect -3761 493 -3727 527
rect -3761 425 -3727 459
rect -3761 357 -3727 391
rect -3761 289 -3727 323
rect -3761 221 -3727 255
rect -3761 153 -3727 187
rect -3761 85 -3727 119
rect -3761 17 -3727 51
rect -3761 -51 -3727 -17
rect -3761 -119 -3727 -85
rect -3761 -187 -3727 -153
rect -3761 -255 -3727 -221
rect -3761 -323 -3727 -289
rect -3761 -391 -3727 -357
rect -3761 -459 -3727 -425
rect -3761 -527 -3727 -493
rect -3761 -595 -3727 -561
rect -3761 -663 -3727 -629
rect -3761 -731 -3727 -697
rect -3761 -799 -3727 -765
rect -3761 -867 -3727 -833
rect -3761 -935 -3727 -901
rect -3761 -1004 -3727 -969
rect -3665 969 -3631 1004
rect -3665 901 -3631 935
rect -3665 833 -3631 867
rect -3665 765 -3631 799
rect -3665 697 -3631 731
rect -3665 629 -3631 663
rect -3665 561 -3631 595
rect -3665 493 -3631 527
rect -3665 425 -3631 459
rect -3665 357 -3631 391
rect -3665 289 -3631 323
rect -3665 221 -3631 255
rect -3665 153 -3631 187
rect -3665 85 -3631 119
rect -3665 17 -3631 51
rect -3665 -51 -3631 -17
rect -3665 -119 -3631 -85
rect -3665 -187 -3631 -153
rect -3665 -255 -3631 -221
rect -3665 -323 -3631 -289
rect -3665 -391 -3631 -357
rect -3665 -459 -3631 -425
rect -3665 -527 -3631 -493
rect -3665 -595 -3631 -561
rect -3665 -663 -3631 -629
rect -3665 -731 -3631 -697
rect -3665 -799 -3631 -765
rect -3665 -867 -3631 -833
rect -3665 -935 -3631 -901
rect -3665 -1004 -3631 -969
rect -3569 969 -3535 1004
rect -3569 901 -3535 935
rect -3569 833 -3535 867
rect -3569 765 -3535 799
rect -3569 697 -3535 731
rect -3569 629 -3535 663
rect -3569 561 -3535 595
rect -3569 493 -3535 527
rect -3569 425 -3535 459
rect -3569 357 -3535 391
rect -3569 289 -3535 323
rect -3569 221 -3535 255
rect -3569 153 -3535 187
rect -3569 85 -3535 119
rect -3569 17 -3535 51
rect -3569 -51 -3535 -17
rect -3569 -119 -3535 -85
rect -3569 -187 -3535 -153
rect -3569 -255 -3535 -221
rect -3569 -323 -3535 -289
rect -3569 -391 -3535 -357
rect -3569 -459 -3535 -425
rect -3569 -527 -3535 -493
rect -3569 -595 -3535 -561
rect -3569 -663 -3535 -629
rect -3569 -731 -3535 -697
rect -3569 -799 -3535 -765
rect -3569 -867 -3535 -833
rect -3569 -935 -3535 -901
rect -3569 -1004 -3535 -969
rect -3473 969 -3439 1004
rect -3473 901 -3439 935
rect -3473 833 -3439 867
rect -3473 765 -3439 799
rect -3473 697 -3439 731
rect -3473 629 -3439 663
rect -3473 561 -3439 595
rect -3473 493 -3439 527
rect -3473 425 -3439 459
rect -3473 357 -3439 391
rect -3473 289 -3439 323
rect -3473 221 -3439 255
rect -3473 153 -3439 187
rect -3473 85 -3439 119
rect -3473 17 -3439 51
rect -3473 -51 -3439 -17
rect -3473 -119 -3439 -85
rect -3473 -187 -3439 -153
rect -3473 -255 -3439 -221
rect -3473 -323 -3439 -289
rect -3473 -391 -3439 -357
rect -3473 -459 -3439 -425
rect -3473 -527 -3439 -493
rect -3473 -595 -3439 -561
rect -3473 -663 -3439 -629
rect -3473 -731 -3439 -697
rect -3473 -799 -3439 -765
rect -3473 -867 -3439 -833
rect -3473 -935 -3439 -901
rect -3473 -1004 -3439 -969
rect -3377 969 -3343 1004
rect -3377 901 -3343 935
rect -3377 833 -3343 867
rect -3377 765 -3343 799
rect -3377 697 -3343 731
rect -3377 629 -3343 663
rect -3377 561 -3343 595
rect -3377 493 -3343 527
rect -3377 425 -3343 459
rect -3377 357 -3343 391
rect -3377 289 -3343 323
rect -3377 221 -3343 255
rect -3377 153 -3343 187
rect -3377 85 -3343 119
rect -3377 17 -3343 51
rect -3377 -51 -3343 -17
rect -3377 -119 -3343 -85
rect -3377 -187 -3343 -153
rect -3377 -255 -3343 -221
rect -3377 -323 -3343 -289
rect -3377 -391 -3343 -357
rect -3377 -459 -3343 -425
rect -3377 -527 -3343 -493
rect -3377 -595 -3343 -561
rect -3377 -663 -3343 -629
rect -3377 -731 -3343 -697
rect -3377 -799 -3343 -765
rect -3377 -867 -3343 -833
rect -3377 -935 -3343 -901
rect -3377 -1004 -3343 -969
rect -3281 969 -3247 1004
rect -3281 901 -3247 935
rect -3281 833 -3247 867
rect -3281 765 -3247 799
rect -3281 697 -3247 731
rect -3281 629 -3247 663
rect -3281 561 -3247 595
rect -3281 493 -3247 527
rect -3281 425 -3247 459
rect -3281 357 -3247 391
rect -3281 289 -3247 323
rect -3281 221 -3247 255
rect -3281 153 -3247 187
rect -3281 85 -3247 119
rect -3281 17 -3247 51
rect -3281 -51 -3247 -17
rect -3281 -119 -3247 -85
rect -3281 -187 -3247 -153
rect -3281 -255 -3247 -221
rect -3281 -323 -3247 -289
rect -3281 -391 -3247 -357
rect -3281 -459 -3247 -425
rect -3281 -527 -3247 -493
rect -3281 -595 -3247 -561
rect -3281 -663 -3247 -629
rect -3281 -731 -3247 -697
rect -3281 -799 -3247 -765
rect -3281 -867 -3247 -833
rect -3281 -935 -3247 -901
rect -3281 -1004 -3247 -969
rect -3185 969 -3151 1004
rect -3185 901 -3151 935
rect -3185 833 -3151 867
rect -3185 765 -3151 799
rect -3185 697 -3151 731
rect -3185 629 -3151 663
rect -3185 561 -3151 595
rect -3185 493 -3151 527
rect -3185 425 -3151 459
rect -3185 357 -3151 391
rect -3185 289 -3151 323
rect -3185 221 -3151 255
rect -3185 153 -3151 187
rect -3185 85 -3151 119
rect -3185 17 -3151 51
rect -3185 -51 -3151 -17
rect -3185 -119 -3151 -85
rect -3185 -187 -3151 -153
rect -3185 -255 -3151 -221
rect -3185 -323 -3151 -289
rect -3185 -391 -3151 -357
rect -3185 -459 -3151 -425
rect -3185 -527 -3151 -493
rect -3185 -595 -3151 -561
rect -3185 -663 -3151 -629
rect -3185 -731 -3151 -697
rect -3185 -799 -3151 -765
rect -3185 -867 -3151 -833
rect -3185 -935 -3151 -901
rect -3185 -1004 -3151 -969
rect -3089 969 -3055 1004
rect -3089 901 -3055 935
rect -3089 833 -3055 867
rect -3089 765 -3055 799
rect -3089 697 -3055 731
rect -3089 629 -3055 663
rect -3089 561 -3055 595
rect -3089 493 -3055 527
rect -3089 425 -3055 459
rect -3089 357 -3055 391
rect -3089 289 -3055 323
rect -3089 221 -3055 255
rect -3089 153 -3055 187
rect -3089 85 -3055 119
rect -3089 17 -3055 51
rect -3089 -51 -3055 -17
rect -3089 -119 -3055 -85
rect -3089 -187 -3055 -153
rect -3089 -255 -3055 -221
rect -3089 -323 -3055 -289
rect -3089 -391 -3055 -357
rect -3089 -459 -3055 -425
rect -3089 -527 -3055 -493
rect -3089 -595 -3055 -561
rect -3089 -663 -3055 -629
rect -3089 -731 -3055 -697
rect -3089 -799 -3055 -765
rect -3089 -867 -3055 -833
rect -3089 -935 -3055 -901
rect -3089 -1004 -3055 -969
rect -2993 969 -2959 1004
rect -2993 901 -2959 935
rect -2993 833 -2959 867
rect -2993 765 -2959 799
rect -2993 697 -2959 731
rect -2993 629 -2959 663
rect -2993 561 -2959 595
rect -2993 493 -2959 527
rect -2993 425 -2959 459
rect -2993 357 -2959 391
rect -2993 289 -2959 323
rect -2993 221 -2959 255
rect -2993 153 -2959 187
rect -2993 85 -2959 119
rect -2993 17 -2959 51
rect -2993 -51 -2959 -17
rect -2993 -119 -2959 -85
rect -2993 -187 -2959 -153
rect -2993 -255 -2959 -221
rect -2993 -323 -2959 -289
rect -2993 -391 -2959 -357
rect -2993 -459 -2959 -425
rect -2993 -527 -2959 -493
rect -2993 -595 -2959 -561
rect -2993 -663 -2959 -629
rect -2993 -731 -2959 -697
rect -2993 -799 -2959 -765
rect -2993 -867 -2959 -833
rect -2993 -935 -2959 -901
rect -2993 -1004 -2959 -969
rect -2897 969 -2863 1004
rect -2897 901 -2863 935
rect -2897 833 -2863 867
rect -2897 765 -2863 799
rect -2897 697 -2863 731
rect -2897 629 -2863 663
rect -2897 561 -2863 595
rect -2897 493 -2863 527
rect -2897 425 -2863 459
rect -2897 357 -2863 391
rect -2897 289 -2863 323
rect -2897 221 -2863 255
rect -2897 153 -2863 187
rect -2897 85 -2863 119
rect -2897 17 -2863 51
rect -2897 -51 -2863 -17
rect -2897 -119 -2863 -85
rect -2897 -187 -2863 -153
rect -2897 -255 -2863 -221
rect -2897 -323 -2863 -289
rect -2897 -391 -2863 -357
rect -2897 -459 -2863 -425
rect -2897 -527 -2863 -493
rect -2897 -595 -2863 -561
rect -2897 -663 -2863 -629
rect -2897 -731 -2863 -697
rect -2897 -799 -2863 -765
rect -2897 -867 -2863 -833
rect -2897 -935 -2863 -901
rect -2897 -1004 -2863 -969
rect -2801 969 -2767 1004
rect -2801 901 -2767 935
rect -2801 833 -2767 867
rect -2801 765 -2767 799
rect -2801 697 -2767 731
rect -2801 629 -2767 663
rect -2801 561 -2767 595
rect -2801 493 -2767 527
rect -2801 425 -2767 459
rect -2801 357 -2767 391
rect -2801 289 -2767 323
rect -2801 221 -2767 255
rect -2801 153 -2767 187
rect -2801 85 -2767 119
rect -2801 17 -2767 51
rect -2801 -51 -2767 -17
rect -2801 -119 -2767 -85
rect -2801 -187 -2767 -153
rect -2801 -255 -2767 -221
rect -2801 -323 -2767 -289
rect -2801 -391 -2767 -357
rect -2801 -459 -2767 -425
rect -2801 -527 -2767 -493
rect -2801 -595 -2767 -561
rect -2801 -663 -2767 -629
rect -2801 -731 -2767 -697
rect -2801 -799 -2767 -765
rect -2801 -867 -2767 -833
rect -2801 -935 -2767 -901
rect -2801 -1004 -2767 -969
rect -2705 969 -2671 1004
rect -2705 901 -2671 935
rect -2705 833 -2671 867
rect -2705 765 -2671 799
rect -2705 697 -2671 731
rect -2705 629 -2671 663
rect -2705 561 -2671 595
rect -2705 493 -2671 527
rect -2705 425 -2671 459
rect -2705 357 -2671 391
rect -2705 289 -2671 323
rect -2705 221 -2671 255
rect -2705 153 -2671 187
rect -2705 85 -2671 119
rect -2705 17 -2671 51
rect -2705 -51 -2671 -17
rect -2705 -119 -2671 -85
rect -2705 -187 -2671 -153
rect -2705 -255 -2671 -221
rect -2705 -323 -2671 -289
rect -2705 -391 -2671 -357
rect -2705 -459 -2671 -425
rect -2705 -527 -2671 -493
rect -2705 -595 -2671 -561
rect -2705 -663 -2671 -629
rect -2705 -731 -2671 -697
rect -2705 -799 -2671 -765
rect -2705 -867 -2671 -833
rect -2705 -935 -2671 -901
rect -2705 -1004 -2671 -969
rect -2609 969 -2575 1004
rect -2609 901 -2575 935
rect -2609 833 -2575 867
rect -2609 765 -2575 799
rect -2609 697 -2575 731
rect -2609 629 -2575 663
rect -2609 561 -2575 595
rect -2609 493 -2575 527
rect -2609 425 -2575 459
rect -2609 357 -2575 391
rect -2609 289 -2575 323
rect -2609 221 -2575 255
rect -2609 153 -2575 187
rect -2609 85 -2575 119
rect -2609 17 -2575 51
rect -2609 -51 -2575 -17
rect -2609 -119 -2575 -85
rect -2609 -187 -2575 -153
rect -2609 -255 -2575 -221
rect -2609 -323 -2575 -289
rect -2609 -391 -2575 -357
rect -2609 -459 -2575 -425
rect -2609 -527 -2575 -493
rect -2609 -595 -2575 -561
rect -2609 -663 -2575 -629
rect -2609 -731 -2575 -697
rect -2609 -799 -2575 -765
rect -2609 -867 -2575 -833
rect -2609 -935 -2575 -901
rect -2609 -1004 -2575 -969
rect -2513 969 -2479 1004
rect -2513 901 -2479 935
rect -2513 833 -2479 867
rect -2513 765 -2479 799
rect -2513 697 -2479 731
rect -2513 629 -2479 663
rect -2513 561 -2479 595
rect -2513 493 -2479 527
rect -2513 425 -2479 459
rect -2513 357 -2479 391
rect -2513 289 -2479 323
rect -2513 221 -2479 255
rect -2513 153 -2479 187
rect -2513 85 -2479 119
rect -2513 17 -2479 51
rect -2513 -51 -2479 -17
rect -2513 -119 -2479 -85
rect -2513 -187 -2479 -153
rect -2513 -255 -2479 -221
rect -2513 -323 -2479 -289
rect -2513 -391 -2479 -357
rect -2513 -459 -2479 -425
rect -2513 -527 -2479 -493
rect -2513 -595 -2479 -561
rect -2513 -663 -2479 -629
rect -2513 -731 -2479 -697
rect -2513 -799 -2479 -765
rect -2513 -867 -2479 -833
rect -2513 -935 -2479 -901
rect -2513 -1004 -2479 -969
rect -2417 969 -2383 1004
rect -2417 901 -2383 935
rect -2417 833 -2383 867
rect -2417 765 -2383 799
rect -2417 697 -2383 731
rect -2417 629 -2383 663
rect -2417 561 -2383 595
rect -2417 493 -2383 527
rect -2417 425 -2383 459
rect -2417 357 -2383 391
rect -2417 289 -2383 323
rect -2417 221 -2383 255
rect -2417 153 -2383 187
rect -2417 85 -2383 119
rect -2417 17 -2383 51
rect -2417 -51 -2383 -17
rect -2417 -119 -2383 -85
rect -2417 -187 -2383 -153
rect -2417 -255 -2383 -221
rect -2417 -323 -2383 -289
rect -2417 -391 -2383 -357
rect -2417 -459 -2383 -425
rect -2417 -527 -2383 -493
rect -2417 -595 -2383 -561
rect -2417 -663 -2383 -629
rect -2417 -731 -2383 -697
rect -2417 -799 -2383 -765
rect -2417 -867 -2383 -833
rect -2417 -935 -2383 -901
rect -2417 -1004 -2383 -969
rect -2321 969 -2287 1004
rect -2321 901 -2287 935
rect -2321 833 -2287 867
rect -2321 765 -2287 799
rect -2321 697 -2287 731
rect -2321 629 -2287 663
rect -2321 561 -2287 595
rect -2321 493 -2287 527
rect -2321 425 -2287 459
rect -2321 357 -2287 391
rect -2321 289 -2287 323
rect -2321 221 -2287 255
rect -2321 153 -2287 187
rect -2321 85 -2287 119
rect -2321 17 -2287 51
rect -2321 -51 -2287 -17
rect -2321 -119 -2287 -85
rect -2321 -187 -2287 -153
rect -2321 -255 -2287 -221
rect -2321 -323 -2287 -289
rect -2321 -391 -2287 -357
rect -2321 -459 -2287 -425
rect -2321 -527 -2287 -493
rect -2321 -595 -2287 -561
rect -2321 -663 -2287 -629
rect -2321 -731 -2287 -697
rect -2321 -799 -2287 -765
rect -2321 -867 -2287 -833
rect -2321 -935 -2287 -901
rect -2321 -1004 -2287 -969
rect -2225 969 -2191 1004
rect -2225 901 -2191 935
rect -2225 833 -2191 867
rect -2225 765 -2191 799
rect -2225 697 -2191 731
rect -2225 629 -2191 663
rect -2225 561 -2191 595
rect -2225 493 -2191 527
rect -2225 425 -2191 459
rect -2225 357 -2191 391
rect -2225 289 -2191 323
rect -2225 221 -2191 255
rect -2225 153 -2191 187
rect -2225 85 -2191 119
rect -2225 17 -2191 51
rect -2225 -51 -2191 -17
rect -2225 -119 -2191 -85
rect -2225 -187 -2191 -153
rect -2225 -255 -2191 -221
rect -2225 -323 -2191 -289
rect -2225 -391 -2191 -357
rect -2225 -459 -2191 -425
rect -2225 -527 -2191 -493
rect -2225 -595 -2191 -561
rect -2225 -663 -2191 -629
rect -2225 -731 -2191 -697
rect -2225 -799 -2191 -765
rect -2225 -867 -2191 -833
rect -2225 -935 -2191 -901
rect -2225 -1004 -2191 -969
rect -2129 969 -2095 1004
rect -2129 901 -2095 935
rect -2129 833 -2095 867
rect -2129 765 -2095 799
rect -2129 697 -2095 731
rect -2129 629 -2095 663
rect -2129 561 -2095 595
rect -2129 493 -2095 527
rect -2129 425 -2095 459
rect -2129 357 -2095 391
rect -2129 289 -2095 323
rect -2129 221 -2095 255
rect -2129 153 -2095 187
rect -2129 85 -2095 119
rect -2129 17 -2095 51
rect -2129 -51 -2095 -17
rect -2129 -119 -2095 -85
rect -2129 -187 -2095 -153
rect -2129 -255 -2095 -221
rect -2129 -323 -2095 -289
rect -2129 -391 -2095 -357
rect -2129 -459 -2095 -425
rect -2129 -527 -2095 -493
rect -2129 -595 -2095 -561
rect -2129 -663 -2095 -629
rect -2129 -731 -2095 -697
rect -2129 -799 -2095 -765
rect -2129 -867 -2095 -833
rect -2129 -935 -2095 -901
rect -2129 -1004 -2095 -969
rect -2033 969 -1999 1004
rect -2033 901 -1999 935
rect -2033 833 -1999 867
rect -2033 765 -1999 799
rect -2033 697 -1999 731
rect -2033 629 -1999 663
rect -2033 561 -1999 595
rect -2033 493 -1999 527
rect -2033 425 -1999 459
rect -2033 357 -1999 391
rect -2033 289 -1999 323
rect -2033 221 -1999 255
rect -2033 153 -1999 187
rect -2033 85 -1999 119
rect -2033 17 -1999 51
rect -2033 -51 -1999 -17
rect -2033 -119 -1999 -85
rect -2033 -187 -1999 -153
rect -2033 -255 -1999 -221
rect -2033 -323 -1999 -289
rect -2033 -391 -1999 -357
rect -2033 -459 -1999 -425
rect -2033 -527 -1999 -493
rect -2033 -595 -1999 -561
rect -2033 -663 -1999 -629
rect -2033 -731 -1999 -697
rect -2033 -799 -1999 -765
rect -2033 -867 -1999 -833
rect -2033 -935 -1999 -901
rect -2033 -1004 -1999 -969
rect -1937 969 -1903 1004
rect -1937 901 -1903 935
rect -1937 833 -1903 867
rect -1937 765 -1903 799
rect -1937 697 -1903 731
rect -1937 629 -1903 663
rect -1937 561 -1903 595
rect -1937 493 -1903 527
rect -1937 425 -1903 459
rect -1937 357 -1903 391
rect -1937 289 -1903 323
rect -1937 221 -1903 255
rect -1937 153 -1903 187
rect -1937 85 -1903 119
rect -1937 17 -1903 51
rect -1937 -51 -1903 -17
rect -1937 -119 -1903 -85
rect -1937 -187 -1903 -153
rect -1937 -255 -1903 -221
rect -1937 -323 -1903 -289
rect -1937 -391 -1903 -357
rect -1937 -459 -1903 -425
rect -1937 -527 -1903 -493
rect -1937 -595 -1903 -561
rect -1937 -663 -1903 -629
rect -1937 -731 -1903 -697
rect -1937 -799 -1903 -765
rect -1937 -867 -1903 -833
rect -1937 -935 -1903 -901
rect -1937 -1004 -1903 -969
rect -1841 969 -1807 1004
rect -1841 901 -1807 935
rect -1841 833 -1807 867
rect -1841 765 -1807 799
rect -1841 697 -1807 731
rect -1841 629 -1807 663
rect -1841 561 -1807 595
rect -1841 493 -1807 527
rect -1841 425 -1807 459
rect -1841 357 -1807 391
rect -1841 289 -1807 323
rect -1841 221 -1807 255
rect -1841 153 -1807 187
rect -1841 85 -1807 119
rect -1841 17 -1807 51
rect -1841 -51 -1807 -17
rect -1841 -119 -1807 -85
rect -1841 -187 -1807 -153
rect -1841 -255 -1807 -221
rect -1841 -323 -1807 -289
rect -1841 -391 -1807 -357
rect -1841 -459 -1807 -425
rect -1841 -527 -1807 -493
rect -1841 -595 -1807 -561
rect -1841 -663 -1807 -629
rect -1841 -731 -1807 -697
rect -1841 -799 -1807 -765
rect -1841 -867 -1807 -833
rect -1841 -935 -1807 -901
rect -1841 -1004 -1807 -969
rect -1745 969 -1711 1004
rect -1745 901 -1711 935
rect -1745 833 -1711 867
rect -1745 765 -1711 799
rect -1745 697 -1711 731
rect -1745 629 -1711 663
rect -1745 561 -1711 595
rect -1745 493 -1711 527
rect -1745 425 -1711 459
rect -1745 357 -1711 391
rect -1745 289 -1711 323
rect -1745 221 -1711 255
rect -1745 153 -1711 187
rect -1745 85 -1711 119
rect -1745 17 -1711 51
rect -1745 -51 -1711 -17
rect -1745 -119 -1711 -85
rect -1745 -187 -1711 -153
rect -1745 -255 -1711 -221
rect -1745 -323 -1711 -289
rect -1745 -391 -1711 -357
rect -1745 -459 -1711 -425
rect -1745 -527 -1711 -493
rect -1745 -595 -1711 -561
rect -1745 -663 -1711 -629
rect -1745 -731 -1711 -697
rect -1745 -799 -1711 -765
rect -1745 -867 -1711 -833
rect -1745 -935 -1711 -901
rect -1745 -1004 -1711 -969
rect -1649 969 -1615 1004
rect -1649 901 -1615 935
rect -1649 833 -1615 867
rect -1649 765 -1615 799
rect -1649 697 -1615 731
rect -1649 629 -1615 663
rect -1649 561 -1615 595
rect -1649 493 -1615 527
rect -1649 425 -1615 459
rect -1649 357 -1615 391
rect -1649 289 -1615 323
rect -1649 221 -1615 255
rect -1649 153 -1615 187
rect -1649 85 -1615 119
rect -1649 17 -1615 51
rect -1649 -51 -1615 -17
rect -1649 -119 -1615 -85
rect -1649 -187 -1615 -153
rect -1649 -255 -1615 -221
rect -1649 -323 -1615 -289
rect -1649 -391 -1615 -357
rect -1649 -459 -1615 -425
rect -1649 -527 -1615 -493
rect -1649 -595 -1615 -561
rect -1649 -663 -1615 -629
rect -1649 -731 -1615 -697
rect -1649 -799 -1615 -765
rect -1649 -867 -1615 -833
rect -1649 -935 -1615 -901
rect -1649 -1004 -1615 -969
rect -1553 969 -1519 1004
rect -1553 901 -1519 935
rect -1553 833 -1519 867
rect -1553 765 -1519 799
rect -1553 697 -1519 731
rect -1553 629 -1519 663
rect -1553 561 -1519 595
rect -1553 493 -1519 527
rect -1553 425 -1519 459
rect -1553 357 -1519 391
rect -1553 289 -1519 323
rect -1553 221 -1519 255
rect -1553 153 -1519 187
rect -1553 85 -1519 119
rect -1553 17 -1519 51
rect -1553 -51 -1519 -17
rect -1553 -119 -1519 -85
rect -1553 -187 -1519 -153
rect -1553 -255 -1519 -221
rect -1553 -323 -1519 -289
rect -1553 -391 -1519 -357
rect -1553 -459 -1519 -425
rect -1553 -527 -1519 -493
rect -1553 -595 -1519 -561
rect -1553 -663 -1519 -629
rect -1553 -731 -1519 -697
rect -1553 -799 -1519 -765
rect -1553 -867 -1519 -833
rect -1553 -935 -1519 -901
rect -1553 -1004 -1519 -969
rect -1457 969 -1423 1004
rect -1457 901 -1423 935
rect -1457 833 -1423 867
rect -1457 765 -1423 799
rect -1457 697 -1423 731
rect -1457 629 -1423 663
rect -1457 561 -1423 595
rect -1457 493 -1423 527
rect -1457 425 -1423 459
rect -1457 357 -1423 391
rect -1457 289 -1423 323
rect -1457 221 -1423 255
rect -1457 153 -1423 187
rect -1457 85 -1423 119
rect -1457 17 -1423 51
rect -1457 -51 -1423 -17
rect -1457 -119 -1423 -85
rect -1457 -187 -1423 -153
rect -1457 -255 -1423 -221
rect -1457 -323 -1423 -289
rect -1457 -391 -1423 -357
rect -1457 -459 -1423 -425
rect -1457 -527 -1423 -493
rect -1457 -595 -1423 -561
rect -1457 -663 -1423 -629
rect -1457 -731 -1423 -697
rect -1457 -799 -1423 -765
rect -1457 -867 -1423 -833
rect -1457 -935 -1423 -901
rect -1457 -1004 -1423 -969
rect -1361 969 -1327 1004
rect -1361 901 -1327 935
rect -1361 833 -1327 867
rect -1361 765 -1327 799
rect -1361 697 -1327 731
rect -1361 629 -1327 663
rect -1361 561 -1327 595
rect -1361 493 -1327 527
rect -1361 425 -1327 459
rect -1361 357 -1327 391
rect -1361 289 -1327 323
rect -1361 221 -1327 255
rect -1361 153 -1327 187
rect -1361 85 -1327 119
rect -1361 17 -1327 51
rect -1361 -51 -1327 -17
rect -1361 -119 -1327 -85
rect -1361 -187 -1327 -153
rect -1361 -255 -1327 -221
rect -1361 -323 -1327 -289
rect -1361 -391 -1327 -357
rect -1361 -459 -1327 -425
rect -1361 -527 -1327 -493
rect -1361 -595 -1327 -561
rect -1361 -663 -1327 -629
rect -1361 -731 -1327 -697
rect -1361 -799 -1327 -765
rect -1361 -867 -1327 -833
rect -1361 -935 -1327 -901
rect -1361 -1004 -1327 -969
rect -1265 969 -1231 1004
rect -1265 901 -1231 935
rect -1265 833 -1231 867
rect -1265 765 -1231 799
rect -1265 697 -1231 731
rect -1265 629 -1231 663
rect -1265 561 -1231 595
rect -1265 493 -1231 527
rect -1265 425 -1231 459
rect -1265 357 -1231 391
rect -1265 289 -1231 323
rect -1265 221 -1231 255
rect -1265 153 -1231 187
rect -1265 85 -1231 119
rect -1265 17 -1231 51
rect -1265 -51 -1231 -17
rect -1265 -119 -1231 -85
rect -1265 -187 -1231 -153
rect -1265 -255 -1231 -221
rect -1265 -323 -1231 -289
rect -1265 -391 -1231 -357
rect -1265 -459 -1231 -425
rect -1265 -527 -1231 -493
rect -1265 -595 -1231 -561
rect -1265 -663 -1231 -629
rect -1265 -731 -1231 -697
rect -1265 -799 -1231 -765
rect -1265 -867 -1231 -833
rect -1265 -935 -1231 -901
rect -1265 -1004 -1231 -969
rect -1169 969 -1135 1004
rect -1169 901 -1135 935
rect -1169 833 -1135 867
rect -1169 765 -1135 799
rect -1169 697 -1135 731
rect -1169 629 -1135 663
rect -1169 561 -1135 595
rect -1169 493 -1135 527
rect -1169 425 -1135 459
rect -1169 357 -1135 391
rect -1169 289 -1135 323
rect -1169 221 -1135 255
rect -1169 153 -1135 187
rect -1169 85 -1135 119
rect -1169 17 -1135 51
rect -1169 -51 -1135 -17
rect -1169 -119 -1135 -85
rect -1169 -187 -1135 -153
rect -1169 -255 -1135 -221
rect -1169 -323 -1135 -289
rect -1169 -391 -1135 -357
rect -1169 -459 -1135 -425
rect -1169 -527 -1135 -493
rect -1169 -595 -1135 -561
rect -1169 -663 -1135 -629
rect -1169 -731 -1135 -697
rect -1169 -799 -1135 -765
rect -1169 -867 -1135 -833
rect -1169 -935 -1135 -901
rect -1169 -1004 -1135 -969
rect -1073 969 -1039 1004
rect -1073 901 -1039 935
rect -1073 833 -1039 867
rect -1073 765 -1039 799
rect -1073 697 -1039 731
rect -1073 629 -1039 663
rect -1073 561 -1039 595
rect -1073 493 -1039 527
rect -1073 425 -1039 459
rect -1073 357 -1039 391
rect -1073 289 -1039 323
rect -1073 221 -1039 255
rect -1073 153 -1039 187
rect -1073 85 -1039 119
rect -1073 17 -1039 51
rect -1073 -51 -1039 -17
rect -1073 -119 -1039 -85
rect -1073 -187 -1039 -153
rect -1073 -255 -1039 -221
rect -1073 -323 -1039 -289
rect -1073 -391 -1039 -357
rect -1073 -459 -1039 -425
rect -1073 -527 -1039 -493
rect -1073 -595 -1039 -561
rect -1073 -663 -1039 -629
rect -1073 -731 -1039 -697
rect -1073 -799 -1039 -765
rect -1073 -867 -1039 -833
rect -1073 -935 -1039 -901
rect -1073 -1004 -1039 -969
rect -977 969 -943 1004
rect -977 901 -943 935
rect -977 833 -943 867
rect -977 765 -943 799
rect -977 697 -943 731
rect -977 629 -943 663
rect -977 561 -943 595
rect -977 493 -943 527
rect -977 425 -943 459
rect -977 357 -943 391
rect -977 289 -943 323
rect -977 221 -943 255
rect -977 153 -943 187
rect -977 85 -943 119
rect -977 17 -943 51
rect -977 -51 -943 -17
rect -977 -119 -943 -85
rect -977 -187 -943 -153
rect -977 -255 -943 -221
rect -977 -323 -943 -289
rect -977 -391 -943 -357
rect -977 -459 -943 -425
rect -977 -527 -943 -493
rect -977 -595 -943 -561
rect -977 -663 -943 -629
rect -977 -731 -943 -697
rect -977 -799 -943 -765
rect -977 -867 -943 -833
rect -977 -935 -943 -901
rect -977 -1004 -943 -969
rect -881 969 -847 1004
rect -881 901 -847 935
rect -881 833 -847 867
rect -881 765 -847 799
rect -881 697 -847 731
rect -881 629 -847 663
rect -881 561 -847 595
rect -881 493 -847 527
rect -881 425 -847 459
rect -881 357 -847 391
rect -881 289 -847 323
rect -881 221 -847 255
rect -881 153 -847 187
rect -881 85 -847 119
rect -881 17 -847 51
rect -881 -51 -847 -17
rect -881 -119 -847 -85
rect -881 -187 -847 -153
rect -881 -255 -847 -221
rect -881 -323 -847 -289
rect -881 -391 -847 -357
rect -881 -459 -847 -425
rect -881 -527 -847 -493
rect -881 -595 -847 -561
rect -881 -663 -847 -629
rect -881 -731 -847 -697
rect -881 -799 -847 -765
rect -881 -867 -847 -833
rect -881 -935 -847 -901
rect -881 -1004 -847 -969
rect -785 969 -751 1004
rect -785 901 -751 935
rect -785 833 -751 867
rect -785 765 -751 799
rect -785 697 -751 731
rect -785 629 -751 663
rect -785 561 -751 595
rect -785 493 -751 527
rect -785 425 -751 459
rect -785 357 -751 391
rect -785 289 -751 323
rect -785 221 -751 255
rect -785 153 -751 187
rect -785 85 -751 119
rect -785 17 -751 51
rect -785 -51 -751 -17
rect -785 -119 -751 -85
rect -785 -187 -751 -153
rect -785 -255 -751 -221
rect -785 -323 -751 -289
rect -785 -391 -751 -357
rect -785 -459 -751 -425
rect -785 -527 -751 -493
rect -785 -595 -751 -561
rect -785 -663 -751 -629
rect -785 -731 -751 -697
rect -785 -799 -751 -765
rect -785 -867 -751 -833
rect -785 -935 -751 -901
rect -785 -1004 -751 -969
rect -689 969 -655 1004
rect -689 901 -655 935
rect -689 833 -655 867
rect -689 765 -655 799
rect -689 697 -655 731
rect -689 629 -655 663
rect -689 561 -655 595
rect -689 493 -655 527
rect -689 425 -655 459
rect -689 357 -655 391
rect -689 289 -655 323
rect -689 221 -655 255
rect -689 153 -655 187
rect -689 85 -655 119
rect -689 17 -655 51
rect -689 -51 -655 -17
rect -689 -119 -655 -85
rect -689 -187 -655 -153
rect -689 -255 -655 -221
rect -689 -323 -655 -289
rect -689 -391 -655 -357
rect -689 -459 -655 -425
rect -689 -527 -655 -493
rect -689 -595 -655 -561
rect -689 -663 -655 -629
rect -689 -731 -655 -697
rect -689 -799 -655 -765
rect -689 -867 -655 -833
rect -689 -935 -655 -901
rect -689 -1004 -655 -969
rect -593 969 -559 1004
rect -593 901 -559 935
rect -593 833 -559 867
rect -593 765 -559 799
rect -593 697 -559 731
rect -593 629 -559 663
rect -593 561 -559 595
rect -593 493 -559 527
rect -593 425 -559 459
rect -593 357 -559 391
rect -593 289 -559 323
rect -593 221 -559 255
rect -593 153 -559 187
rect -593 85 -559 119
rect -593 17 -559 51
rect -593 -51 -559 -17
rect -593 -119 -559 -85
rect -593 -187 -559 -153
rect -593 -255 -559 -221
rect -593 -323 -559 -289
rect -593 -391 -559 -357
rect -593 -459 -559 -425
rect -593 -527 -559 -493
rect -593 -595 -559 -561
rect -593 -663 -559 -629
rect -593 -731 -559 -697
rect -593 -799 -559 -765
rect -593 -867 -559 -833
rect -593 -935 -559 -901
rect -593 -1004 -559 -969
rect -497 969 -463 1004
rect -497 901 -463 935
rect -497 833 -463 867
rect -497 765 -463 799
rect -497 697 -463 731
rect -497 629 -463 663
rect -497 561 -463 595
rect -497 493 -463 527
rect -497 425 -463 459
rect -497 357 -463 391
rect -497 289 -463 323
rect -497 221 -463 255
rect -497 153 -463 187
rect -497 85 -463 119
rect -497 17 -463 51
rect -497 -51 -463 -17
rect -497 -119 -463 -85
rect -497 -187 -463 -153
rect -497 -255 -463 -221
rect -497 -323 -463 -289
rect -497 -391 -463 -357
rect -497 -459 -463 -425
rect -497 -527 -463 -493
rect -497 -595 -463 -561
rect -497 -663 -463 -629
rect -497 -731 -463 -697
rect -497 -799 -463 -765
rect -497 -867 -463 -833
rect -497 -935 -463 -901
rect -497 -1004 -463 -969
rect -401 969 -367 1004
rect -401 901 -367 935
rect -401 833 -367 867
rect -401 765 -367 799
rect -401 697 -367 731
rect -401 629 -367 663
rect -401 561 -367 595
rect -401 493 -367 527
rect -401 425 -367 459
rect -401 357 -367 391
rect -401 289 -367 323
rect -401 221 -367 255
rect -401 153 -367 187
rect -401 85 -367 119
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -119 -367 -85
rect -401 -187 -367 -153
rect -401 -255 -367 -221
rect -401 -323 -367 -289
rect -401 -391 -367 -357
rect -401 -459 -367 -425
rect -401 -527 -367 -493
rect -401 -595 -367 -561
rect -401 -663 -367 -629
rect -401 -731 -367 -697
rect -401 -799 -367 -765
rect -401 -867 -367 -833
rect -401 -935 -367 -901
rect -401 -1004 -367 -969
rect -305 969 -271 1004
rect -305 901 -271 935
rect -305 833 -271 867
rect -305 765 -271 799
rect -305 697 -271 731
rect -305 629 -271 663
rect -305 561 -271 595
rect -305 493 -271 527
rect -305 425 -271 459
rect -305 357 -271 391
rect -305 289 -271 323
rect -305 221 -271 255
rect -305 153 -271 187
rect -305 85 -271 119
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -119 -271 -85
rect -305 -187 -271 -153
rect -305 -255 -271 -221
rect -305 -323 -271 -289
rect -305 -391 -271 -357
rect -305 -459 -271 -425
rect -305 -527 -271 -493
rect -305 -595 -271 -561
rect -305 -663 -271 -629
rect -305 -731 -271 -697
rect -305 -799 -271 -765
rect -305 -867 -271 -833
rect -305 -935 -271 -901
rect -305 -1004 -271 -969
rect -209 969 -175 1004
rect -209 901 -175 935
rect -209 833 -175 867
rect -209 765 -175 799
rect -209 697 -175 731
rect -209 629 -175 663
rect -209 561 -175 595
rect -209 493 -175 527
rect -209 425 -175 459
rect -209 357 -175 391
rect -209 289 -175 323
rect -209 221 -175 255
rect -209 153 -175 187
rect -209 85 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -85
rect -209 -187 -175 -153
rect -209 -255 -175 -221
rect -209 -323 -175 -289
rect -209 -391 -175 -357
rect -209 -459 -175 -425
rect -209 -527 -175 -493
rect -209 -595 -175 -561
rect -209 -663 -175 -629
rect -209 -731 -175 -697
rect -209 -799 -175 -765
rect -209 -867 -175 -833
rect -209 -935 -175 -901
rect -209 -1004 -175 -969
rect -113 969 -79 1004
rect -113 901 -79 935
rect -113 833 -79 867
rect -113 765 -79 799
rect -113 697 -79 731
rect -113 629 -79 663
rect -113 561 -79 595
rect -113 493 -79 527
rect -113 425 -79 459
rect -113 357 -79 391
rect -113 289 -79 323
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -113 -323 -79 -289
rect -113 -391 -79 -357
rect -113 -459 -79 -425
rect -113 -527 -79 -493
rect -113 -595 -79 -561
rect -113 -663 -79 -629
rect -113 -731 -79 -697
rect -113 -799 -79 -765
rect -113 -867 -79 -833
rect -113 -935 -79 -901
rect -113 -1004 -79 -969
rect -17 969 17 1004
rect -17 901 17 935
rect -17 833 17 867
rect -17 765 17 799
rect -17 697 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -697
rect -17 -799 17 -765
rect -17 -867 17 -833
rect -17 -935 17 -901
rect -17 -1004 17 -969
rect 79 969 113 1004
rect 79 901 113 935
rect 79 833 113 867
rect 79 765 113 799
rect 79 697 113 731
rect 79 629 113 663
rect 79 561 113 595
rect 79 493 113 527
rect 79 425 113 459
rect 79 357 113 391
rect 79 289 113 323
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 79 -323 113 -289
rect 79 -391 113 -357
rect 79 -459 113 -425
rect 79 -527 113 -493
rect 79 -595 113 -561
rect 79 -663 113 -629
rect 79 -731 113 -697
rect 79 -799 113 -765
rect 79 -867 113 -833
rect 79 -935 113 -901
rect 79 -1004 113 -969
rect 175 969 209 1004
rect 175 901 209 935
rect 175 833 209 867
rect 175 765 209 799
rect 175 697 209 731
rect 175 629 209 663
rect 175 561 209 595
rect 175 493 209 527
rect 175 425 209 459
rect 175 357 209 391
rect 175 289 209 323
rect 175 221 209 255
rect 175 153 209 187
rect 175 85 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -85
rect 175 -187 209 -153
rect 175 -255 209 -221
rect 175 -323 209 -289
rect 175 -391 209 -357
rect 175 -459 209 -425
rect 175 -527 209 -493
rect 175 -595 209 -561
rect 175 -663 209 -629
rect 175 -731 209 -697
rect 175 -799 209 -765
rect 175 -867 209 -833
rect 175 -935 209 -901
rect 175 -1004 209 -969
rect 271 969 305 1004
rect 271 901 305 935
rect 271 833 305 867
rect 271 765 305 799
rect 271 697 305 731
rect 271 629 305 663
rect 271 561 305 595
rect 271 493 305 527
rect 271 425 305 459
rect 271 357 305 391
rect 271 289 305 323
rect 271 221 305 255
rect 271 153 305 187
rect 271 85 305 119
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -119 305 -85
rect 271 -187 305 -153
rect 271 -255 305 -221
rect 271 -323 305 -289
rect 271 -391 305 -357
rect 271 -459 305 -425
rect 271 -527 305 -493
rect 271 -595 305 -561
rect 271 -663 305 -629
rect 271 -731 305 -697
rect 271 -799 305 -765
rect 271 -867 305 -833
rect 271 -935 305 -901
rect 271 -1004 305 -969
rect 367 969 401 1004
rect 367 901 401 935
rect 367 833 401 867
rect 367 765 401 799
rect 367 697 401 731
rect 367 629 401 663
rect 367 561 401 595
rect 367 493 401 527
rect 367 425 401 459
rect 367 357 401 391
rect 367 289 401 323
rect 367 221 401 255
rect 367 153 401 187
rect 367 85 401 119
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -119 401 -85
rect 367 -187 401 -153
rect 367 -255 401 -221
rect 367 -323 401 -289
rect 367 -391 401 -357
rect 367 -459 401 -425
rect 367 -527 401 -493
rect 367 -595 401 -561
rect 367 -663 401 -629
rect 367 -731 401 -697
rect 367 -799 401 -765
rect 367 -867 401 -833
rect 367 -935 401 -901
rect 367 -1004 401 -969
rect 463 969 497 1004
rect 463 901 497 935
rect 463 833 497 867
rect 463 765 497 799
rect 463 697 497 731
rect 463 629 497 663
rect 463 561 497 595
rect 463 493 497 527
rect 463 425 497 459
rect 463 357 497 391
rect 463 289 497 323
rect 463 221 497 255
rect 463 153 497 187
rect 463 85 497 119
rect 463 17 497 51
rect 463 -51 497 -17
rect 463 -119 497 -85
rect 463 -187 497 -153
rect 463 -255 497 -221
rect 463 -323 497 -289
rect 463 -391 497 -357
rect 463 -459 497 -425
rect 463 -527 497 -493
rect 463 -595 497 -561
rect 463 -663 497 -629
rect 463 -731 497 -697
rect 463 -799 497 -765
rect 463 -867 497 -833
rect 463 -935 497 -901
rect 463 -1004 497 -969
rect 559 969 593 1004
rect 559 901 593 935
rect 559 833 593 867
rect 559 765 593 799
rect 559 697 593 731
rect 559 629 593 663
rect 559 561 593 595
rect 559 493 593 527
rect 559 425 593 459
rect 559 357 593 391
rect 559 289 593 323
rect 559 221 593 255
rect 559 153 593 187
rect 559 85 593 119
rect 559 17 593 51
rect 559 -51 593 -17
rect 559 -119 593 -85
rect 559 -187 593 -153
rect 559 -255 593 -221
rect 559 -323 593 -289
rect 559 -391 593 -357
rect 559 -459 593 -425
rect 559 -527 593 -493
rect 559 -595 593 -561
rect 559 -663 593 -629
rect 559 -731 593 -697
rect 559 -799 593 -765
rect 559 -867 593 -833
rect 559 -935 593 -901
rect 559 -1004 593 -969
rect 655 969 689 1004
rect 655 901 689 935
rect 655 833 689 867
rect 655 765 689 799
rect 655 697 689 731
rect 655 629 689 663
rect 655 561 689 595
rect 655 493 689 527
rect 655 425 689 459
rect 655 357 689 391
rect 655 289 689 323
rect 655 221 689 255
rect 655 153 689 187
rect 655 85 689 119
rect 655 17 689 51
rect 655 -51 689 -17
rect 655 -119 689 -85
rect 655 -187 689 -153
rect 655 -255 689 -221
rect 655 -323 689 -289
rect 655 -391 689 -357
rect 655 -459 689 -425
rect 655 -527 689 -493
rect 655 -595 689 -561
rect 655 -663 689 -629
rect 655 -731 689 -697
rect 655 -799 689 -765
rect 655 -867 689 -833
rect 655 -935 689 -901
rect 655 -1004 689 -969
rect 751 969 785 1004
rect 751 901 785 935
rect 751 833 785 867
rect 751 765 785 799
rect 751 697 785 731
rect 751 629 785 663
rect 751 561 785 595
rect 751 493 785 527
rect 751 425 785 459
rect 751 357 785 391
rect 751 289 785 323
rect 751 221 785 255
rect 751 153 785 187
rect 751 85 785 119
rect 751 17 785 51
rect 751 -51 785 -17
rect 751 -119 785 -85
rect 751 -187 785 -153
rect 751 -255 785 -221
rect 751 -323 785 -289
rect 751 -391 785 -357
rect 751 -459 785 -425
rect 751 -527 785 -493
rect 751 -595 785 -561
rect 751 -663 785 -629
rect 751 -731 785 -697
rect 751 -799 785 -765
rect 751 -867 785 -833
rect 751 -935 785 -901
rect 751 -1004 785 -969
rect 847 969 881 1004
rect 847 901 881 935
rect 847 833 881 867
rect 847 765 881 799
rect 847 697 881 731
rect 847 629 881 663
rect 847 561 881 595
rect 847 493 881 527
rect 847 425 881 459
rect 847 357 881 391
rect 847 289 881 323
rect 847 221 881 255
rect 847 153 881 187
rect 847 85 881 119
rect 847 17 881 51
rect 847 -51 881 -17
rect 847 -119 881 -85
rect 847 -187 881 -153
rect 847 -255 881 -221
rect 847 -323 881 -289
rect 847 -391 881 -357
rect 847 -459 881 -425
rect 847 -527 881 -493
rect 847 -595 881 -561
rect 847 -663 881 -629
rect 847 -731 881 -697
rect 847 -799 881 -765
rect 847 -867 881 -833
rect 847 -935 881 -901
rect 847 -1004 881 -969
rect 943 969 977 1004
rect 943 901 977 935
rect 943 833 977 867
rect 943 765 977 799
rect 943 697 977 731
rect 943 629 977 663
rect 943 561 977 595
rect 943 493 977 527
rect 943 425 977 459
rect 943 357 977 391
rect 943 289 977 323
rect 943 221 977 255
rect 943 153 977 187
rect 943 85 977 119
rect 943 17 977 51
rect 943 -51 977 -17
rect 943 -119 977 -85
rect 943 -187 977 -153
rect 943 -255 977 -221
rect 943 -323 977 -289
rect 943 -391 977 -357
rect 943 -459 977 -425
rect 943 -527 977 -493
rect 943 -595 977 -561
rect 943 -663 977 -629
rect 943 -731 977 -697
rect 943 -799 977 -765
rect 943 -867 977 -833
rect 943 -935 977 -901
rect 943 -1004 977 -969
rect 1039 969 1073 1004
rect 1039 901 1073 935
rect 1039 833 1073 867
rect 1039 765 1073 799
rect 1039 697 1073 731
rect 1039 629 1073 663
rect 1039 561 1073 595
rect 1039 493 1073 527
rect 1039 425 1073 459
rect 1039 357 1073 391
rect 1039 289 1073 323
rect 1039 221 1073 255
rect 1039 153 1073 187
rect 1039 85 1073 119
rect 1039 17 1073 51
rect 1039 -51 1073 -17
rect 1039 -119 1073 -85
rect 1039 -187 1073 -153
rect 1039 -255 1073 -221
rect 1039 -323 1073 -289
rect 1039 -391 1073 -357
rect 1039 -459 1073 -425
rect 1039 -527 1073 -493
rect 1039 -595 1073 -561
rect 1039 -663 1073 -629
rect 1039 -731 1073 -697
rect 1039 -799 1073 -765
rect 1039 -867 1073 -833
rect 1039 -935 1073 -901
rect 1039 -1004 1073 -969
rect 1135 969 1169 1004
rect 1135 901 1169 935
rect 1135 833 1169 867
rect 1135 765 1169 799
rect 1135 697 1169 731
rect 1135 629 1169 663
rect 1135 561 1169 595
rect 1135 493 1169 527
rect 1135 425 1169 459
rect 1135 357 1169 391
rect 1135 289 1169 323
rect 1135 221 1169 255
rect 1135 153 1169 187
rect 1135 85 1169 119
rect 1135 17 1169 51
rect 1135 -51 1169 -17
rect 1135 -119 1169 -85
rect 1135 -187 1169 -153
rect 1135 -255 1169 -221
rect 1135 -323 1169 -289
rect 1135 -391 1169 -357
rect 1135 -459 1169 -425
rect 1135 -527 1169 -493
rect 1135 -595 1169 -561
rect 1135 -663 1169 -629
rect 1135 -731 1169 -697
rect 1135 -799 1169 -765
rect 1135 -867 1169 -833
rect 1135 -935 1169 -901
rect 1135 -1004 1169 -969
rect 1231 969 1265 1004
rect 1231 901 1265 935
rect 1231 833 1265 867
rect 1231 765 1265 799
rect 1231 697 1265 731
rect 1231 629 1265 663
rect 1231 561 1265 595
rect 1231 493 1265 527
rect 1231 425 1265 459
rect 1231 357 1265 391
rect 1231 289 1265 323
rect 1231 221 1265 255
rect 1231 153 1265 187
rect 1231 85 1265 119
rect 1231 17 1265 51
rect 1231 -51 1265 -17
rect 1231 -119 1265 -85
rect 1231 -187 1265 -153
rect 1231 -255 1265 -221
rect 1231 -323 1265 -289
rect 1231 -391 1265 -357
rect 1231 -459 1265 -425
rect 1231 -527 1265 -493
rect 1231 -595 1265 -561
rect 1231 -663 1265 -629
rect 1231 -731 1265 -697
rect 1231 -799 1265 -765
rect 1231 -867 1265 -833
rect 1231 -935 1265 -901
rect 1231 -1004 1265 -969
rect 1327 969 1361 1004
rect 1327 901 1361 935
rect 1327 833 1361 867
rect 1327 765 1361 799
rect 1327 697 1361 731
rect 1327 629 1361 663
rect 1327 561 1361 595
rect 1327 493 1361 527
rect 1327 425 1361 459
rect 1327 357 1361 391
rect 1327 289 1361 323
rect 1327 221 1361 255
rect 1327 153 1361 187
rect 1327 85 1361 119
rect 1327 17 1361 51
rect 1327 -51 1361 -17
rect 1327 -119 1361 -85
rect 1327 -187 1361 -153
rect 1327 -255 1361 -221
rect 1327 -323 1361 -289
rect 1327 -391 1361 -357
rect 1327 -459 1361 -425
rect 1327 -527 1361 -493
rect 1327 -595 1361 -561
rect 1327 -663 1361 -629
rect 1327 -731 1361 -697
rect 1327 -799 1361 -765
rect 1327 -867 1361 -833
rect 1327 -935 1361 -901
rect 1327 -1004 1361 -969
rect 1423 969 1457 1004
rect 1423 901 1457 935
rect 1423 833 1457 867
rect 1423 765 1457 799
rect 1423 697 1457 731
rect 1423 629 1457 663
rect 1423 561 1457 595
rect 1423 493 1457 527
rect 1423 425 1457 459
rect 1423 357 1457 391
rect 1423 289 1457 323
rect 1423 221 1457 255
rect 1423 153 1457 187
rect 1423 85 1457 119
rect 1423 17 1457 51
rect 1423 -51 1457 -17
rect 1423 -119 1457 -85
rect 1423 -187 1457 -153
rect 1423 -255 1457 -221
rect 1423 -323 1457 -289
rect 1423 -391 1457 -357
rect 1423 -459 1457 -425
rect 1423 -527 1457 -493
rect 1423 -595 1457 -561
rect 1423 -663 1457 -629
rect 1423 -731 1457 -697
rect 1423 -799 1457 -765
rect 1423 -867 1457 -833
rect 1423 -935 1457 -901
rect 1423 -1004 1457 -969
rect 1519 969 1553 1004
rect 1519 901 1553 935
rect 1519 833 1553 867
rect 1519 765 1553 799
rect 1519 697 1553 731
rect 1519 629 1553 663
rect 1519 561 1553 595
rect 1519 493 1553 527
rect 1519 425 1553 459
rect 1519 357 1553 391
rect 1519 289 1553 323
rect 1519 221 1553 255
rect 1519 153 1553 187
rect 1519 85 1553 119
rect 1519 17 1553 51
rect 1519 -51 1553 -17
rect 1519 -119 1553 -85
rect 1519 -187 1553 -153
rect 1519 -255 1553 -221
rect 1519 -323 1553 -289
rect 1519 -391 1553 -357
rect 1519 -459 1553 -425
rect 1519 -527 1553 -493
rect 1519 -595 1553 -561
rect 1519 -663 1553 -629
rect 1519 -731 1553 -697
rect 1519 -799 1553 -765
rect 1519 -867 1553 -833
rect 1519 -935 1553 -901
rect 1519 -1004 1553 -969
rect 1615 969 1649 1004
rect 1615 901 1649 935
rect 1615 833 1649 867
rect 1615 765 1649 799
rect 1615 697 1649 731
rect 1615 629 1649 663
rect 1615 561 1649 595
rect 1615 493 1649 527
rect 1615 425 1649 459
rect 1615 357 1649 391
rect 1615 289 1649 323
rect 1615 221 1649 255
rect 1615 153 1649 187
rect 1615 85 1649 119
rect 1615 17 1649 51
rect 1615 -51 1649 -17
rect 1615 -119 1649 -85
rect 1615 -187 1649 -153
rect 1615 -255 1649 -221
rect 1615 -323 1649 -289
rect 1615 -391 1649 -357
rect 1615 -459 1649 -425
rect 1615 -527 1649 -493
rect 1615 -595 1649 -561
rect 1615 -663 1649 -629
rect 1615 -731 1649 -697
rect 1615 -799 1649 -765
rect 1615 -867 1649 -833
rect 1615 -935 1649 -901
rect 1615 -1004 1649 -969
rect 1711 969 1745 1004
rect 1711 901 1745 935
rect 1711 833 1745 867
rect 1711 765 1745 799
rect 1711 697 1745 731
rect 1711 629 1745 663
rect 1711 561 1745 595
rect 1711 493 1745 527
rect 1711 425 1745 459
rect 1711 357 1745 391
rect 1711 289 1745 323
rect 1711 221 1745 255
rect 1711 153 1745 187
rect 1711 85 1745 119
rect 1711 17 1745 51
rect 1711 -51 1745 -17
rect 1711 -119 1745 -85
rect 1711 -187 1745 -153
rect 1711 -255 1745 -221
rect 1711 -323 1745 -289
rect 1711 -391 1745 -357
rect 1711 -459 1745 -425
rect 1711 -527 1745 -493
rect 1711 -595 1745 -561
rect 1711 -663 1745 -629
rect 1711 -731 1745 -697
rect 1711 -799 1745 -765
rect 1711 -867 1745 -833
rect 1711 -935 1745 -901
rect 1711 -1004 1745 -969
rect 1807 969 1841 1004
rect 1807 901 1841 935
rect 1807 833 1841 867
rect 1807 765 1841 799
rect 1807 697 1841 731
rect 1807 629 1841 663
rect 1807 561 1841 595
rect 1807 493 1841 527
rect 1807 425 1841 459
rect 1807 357 1841 391
rect 1807 289 1841 323
rect 1807 221 1841 255
rect 1807 153 1841 187
rect 1807 85 1841 119
rect 1807 17 1841 51
rect 1807 -51 1841 -17
rect 1807 -119 1841 -85
rect 1807 -187 1841 -153
rect 1807 -255 1841 -221
rect 1807 -323 1841 -289
rect 1807 -391 1841 -357
rect 1807 -459 1841 -425
rect 1807 -527 1841 -493
rect 1807 -595 1841 -561
rect 1807 -663 1841 -629
rect 1807 -731 1841 -697
rect 1807 -799 1841 -765
rect 1807 -867 1841 -833
rect 1807 -935 1841 -901
rect 1807 -1004 1841 -969
rect 1903 969 1937 1004
rect 1903 901 1937 935
rect 1903 833 1937 867
rect 1903 765 1937 799
rect 1903 697 1937 731
rect 1903 629 1937 663
rect 1903 561 1937 595
rect 1903 493 1937 527
rect 1903 425 1937 459
rect 1903 357 1937 391
rect 1903 289 1937 323
rect 1903 221 1937 255
rect 1903 153 1937 187
rect 1903 85 1937 119
rect 1903 17 1937 51
rect 1903 -51 1937 -17
rect 1903 -119 1937 -85
rect 1903 -187 1937 -153
rect 1903 -255 1937 -221
rect 1903 -323 1937 -289
rect 1903 -391 1937 -357
rect 1903 -459 1937 -425
rect 1903 -527 1937 -493
rect 1903 -595 1937 -561
rect 1903 -663 1937 -629
rect 1903 -731 1937 -697
rect 1903 -799 1937 -765
rect 1903 -867 1937 -833
rect 1903 -935 1937 -901
rect 1903 -1004 1937 -969
rect 1999 969 2033 1004
rect 1999 901 2033 935
rect 1999 833 2033 867
rect 1999 765 2033 799
rect 1999 697 2033 731
rect 1999 629 2033 663
rect 1999 561 2033 595
rect 1999 493 2033 527
rect 1999 425 2033 459
rect 1999 357 2033 391
rect 1999 289 2033 323
rect 1999 221 2033 255
rect 1999 153 2033 187
rect 1999 85 2033 119
rect 1999 17 2033 51
rect 1999 -51 2033 -17
rect 1999 -119 2033 -85
rect 1999 -187 2033 -153
rect 1999 -255 2033 -221
rect 1999 -323 2033 -289
rect 1999 -391 2033 -357
rect 1999 -459 2033 -425
rect 1999 -527 2033 -493
rect 1999 -595 2033 -561
rect 1999 -663 2033 -629
rect 1999 -731 2033 -697
rect 1999 -799 2033 -765
rect 1999 -867 2033 -833
rect 1999 -935 2033 -901
rect 1999 -1004 2033 -969
rect 2095 969 2129 1004
rect 2095 901 2129 935
rect 2095 833 2129 867
rect 2095 765 2129 799
rect 2095 697 2129 731
rect 2095 629 2129 663
rect 2095 561 2129 595
rect 2095 493 2129 527
rect 2095 425 2129 459
rect 2095 357 2129 391
rect 2095 289 2129 323
rect 2095 221 2129 255
rect 2095 153 2129 187
rect 2095 85 2129 119
rect 2095 17 2129 51
rect 2095 -51 2129 -17
rect 2095 -119 2129 -85
rect 2095 -187 2129 -153
rect 2095 -255 2129 -221
rect 2095 -323 2129 -289
rect 2095 -391 2129 -357
rect 2095 -459 2129 -425
rect 2095 -527 2129 -493
rect 2095 -595 2129 -561
rect 2095 -663 2129 -629
rect 2095 -731 2129 -697
rect 2095 -799 2129 -765
rect 2095 -867 2129 -833
rect 2095 -935 2129 -901
rect 2095 -1004 2129 -969
rect 2191 969 2225 1004
rect 2191 901 2225 935
rect 2191 833 2225 867
rect 2191 765 2225 799
rect 2191 697 2225 731
rect 2191 629 2225 663
rect 2191 561 2225 595
rect 2191 493 2225 527
rect 2191 425 2225 459
rect 2191 357 2225 391
rect 2191 289 2225 323
rect 2191 221 2225 255
rect 2191 153 2225 187
rect 2191 85 2225 119
rect 2191 17 2225 51
rect 2191 -51 2225 -17
rect 2191 -119 2225 -85
rect 2191 -187 2225 -153
rect 2191 -255 2225 -221
rect 2191 -323 2225 -289
rect 2191 -391 2225 -357
rect 2191 -459 2225 -425
rect 2191 -527 2225 -493
rect 2191 -595 2225 -561
rect 2191 -663 2225 -629
rect 2191 -731 2225 -697
rect 2191 -799 2225 -765
rect 2191 -867 2225 -833
rect 2191 -935 2225 -901
rect 2191 -1004 2225 -969
rect 2287 969 2321 1004
rect 2287 901 2321 935
rect 2287 833 2321 867
rect 2287 765 2321 799
rect 2287 697 2321 731
rect 2287 629 2321 663
rect 2287 561 2321 595
rect 2287 493 2321 527
rect 2287 425 2321 459
rect 2287 357 2321 391
rect 2287 289 2321 323
rect 2287 221 2321 255
rect 2287 153 2321 187
rect 2287 85 2321 119
rect 2287 17 2321 51
rect 2287 -51 2321 -17
rect 2287 -119 2321 -85
rect 2287 -187 2321 -153
rect 2287 -255 2321 -221
rect 2287 -323 2321 -289
rect 2287 -391 2321 -357
rect 2287 -459 2321 -425
rect 2287 -527 2321 -493
rect 2287 -595 2321 -561
rect 2287 -663 2321 -629
rect 2287 -731 2321 -697
rect 2287 -799 2321 -765
rect 2287 -867 2321 -833
rect 2287 -935 2321 -901
rect 2287 -1004 2321 -969
rect 2383 969 2417 1004
rect 2383 901 2417 935
rect 2383 833 2417 867
rect 2383 765 2417 799
rect 2383 697 2417 731
rect 2383 629 2417 663
rect 2383 561 2417 595
rect 2383 493 2417 527
rect 2383 425 2417 459
rect 2383 357 2417 391
rect 2383 289 2417 323
rect 2383 221 2417 255
rect 2383 153 2417 187
rect 2383 85 2417 119
rect 2383 17 2417 51
rect 2383 -51 2417 -17
rect 2383 -119 2417 -85
rect 2383 -187 2417 -153
rect 2383 -255 2417 -221
rect 2383 -323 2417 -289
rect 2383 -391 2417 -357
rect 2383 -459 2417 -425
rect 2383 -527 2417 -493
rect 2383 -595 2417 -561
rect 2383 -663 2417 -629
rect 2383 -731 2417 -697
rect 2383 -799 2417 -765
rect 2383 -867 2417 -833
rect 2383 -935 2417 -901
rect 2383 -1004 2417 -969
rect 2479 969 2513 1004
rect 2479 901 2513 935
rect 2479 833 2513 867
rect 2479 765 2513 799
rect 2479 697 2513 731
rect 2479 629 2513 663
rect 2479 561 2513 595
rect 2479 493 2513 527
rect 2479 425 2513 459
rect 2479 357 2513 391
rect 2479 289 2513 323
rect 2479 221 2513 255
rect 2479 153 2513 187
rect 2479 85 2513 119
rect 2479 17 2513 51
rect 2479 -51 2513 -17
rect 2479 -119 2513 -85
rect 2479 -187 2513 -153
rect 2479 -255 2513 -221
rect 2479 -323 2513 -289
rect 2479 -391 2513 -357
rect 2479 -459 2513 -425
rect 2479 -527 2513 -493
rect 2479 -595 2513 -561
rect 2479 -663 2513 -629
rect 2479 -731 2513 -697
rect 2479 -799 2513 -765
rect 2479 -867 2513 -833
rect 2479 -935 2513 -901
rect 2479 -1004 2513 -969
rect 2575 969 2609 1004
rect 2575 901 2609 935
rect 2575 833 2609 867
rect 2575 765 2609 799
rect 2575 697 2609 731
rect 2575 629 2609 663
rect 2575 561 2609 595
rect 2575 493 2609 527
rect 2575 425 2609 459
rect 2575 357 2609 391
rect 2575 289 2609 323
rect 2575 221 2609 255
rect 2575 153 2609 187
rect 2575 85 2609 119
rect 2575 17 2609 51
rect 2575 -51 2609 -17
rect 2575 -119 2609 -85
rect 2575 -187 2609 -153
rect 2575 -255 2609 -221
rect 2575 -323 2609 -289
rect 2575 -391 2609 -357
rect 2575 -459 2609 -425
rect 2575 -527 2609 -493
rect 2575 -595 2609 -561
rect 2575 -663 2609 -629
rect 2575 -731 2609 -697
rect 2575 -799 2609 -765
rect 2575 -867 2609 -833
rect 2575 -935 2609 -901
rect 2575 -1004 2609 -969
rect 2671 969 2705 1004
rect 2671 901 2705 935
rect 2671 833 2705 867
rect 2671 765 2705 799
rect 2671 697 2705 731
rect 2671 629 2705 663
rect 2671 561 2705 595
rect 2671 493 2705 527
rect 2671 425 2705 459
rect 2671 357 2705 391
rect 2671 289 2705 323
rect 2671 221 2705 255
rect 2671 153 2705 187
rect 2671 85 2705 119
rect 2671 17 2705 51
rect 2671 -51 2705 -17
rect 2671 -119 2705 -85
rect 2671 -187 2705 -153
rect 2671 -255 2705 -221
rect 2671 -323 2705 -289
rect 2671 -391 2705 -357
rect 2671 -459 2705 -425
rect 2671 -527 2705 -493
rect 2671 -595 2705 -561
rect 2671 -663 2705 -629
rect 2671 -731 2705 -697
rect 2671 -799 2705 -765
rect 2671 -867 2705 -833
rect 2671 -935 2705 -901
rect 2671 -1004 2705 -969
rect 2767 969 2801 1004
rect 2767 901 2801 935
rect 2767 833 2801 867
rect 2767 765 2801 799
rect 2767 697 2801 731
rect 2767 629 2801 663
rect 2767 561 2801 595
rect 2767 493 2801 527
rect 2767 425 2801 459
rect 2767 357 2801 391
rect 2767 289 2801 323
rect 2767 221 2801 255
rect 2767 153 2801 187
rect 2767 85 2801 119
rect 2767 17 2801 51
rect 2767 -51 2801 -17
rect 2767 -119 2801 -85
rect 2767 -187 2801 -153
rect 2767 -255 2801 -221
rect 2767 -323 2801 -289
rect 2767 -391 2801 -357
rect 2767 -459 2801 -425
rect 2767 -527 2801 -493
rect 2767 -595 2801 -561
rect 2767 -663 2801 -629
rect 2767 -731 2801 -697
rect 2767 -799 2801 -765
rect 2767 -867 2801 -833
rect 2767 -935 2801 -901
rect 2767 -1004 2801 -969
rect 2863 969 2897 1004
rect 2863 901 2897 935
rect 2863 833 2897 867
rect 2863 765 2897 799
rect 2863 697 2897 731
rect 2863 629 2897 663
rect 2863 561 2897 595
rect 2863 493 2897 527
rect 2863 425 2897 459
rect 2863 357 2897 391
rect 2863 289 2897 323
rect 2863 221 2897 255
rect 2863 153 2897 187
rect 2863 85 2897 119
rect 2863 17 2897 51
rect 2863 -51 2897 -17
rect 2863 -119 2897 -85
rect 2863 -187 2897 -153
rect 2863 -255 2897 -221
rect 2863 -323 2897 -289
rect 2863 -391 2897 -357
rect 2863 -459 2897 -425
rect 2863 -527 2897 -493
rect 2863 -595 2897 -561
rect 2863 -663 2897 -629
rect 2863 -731 2897 -697
rect 2863 -799 2897 -765
rect 2863 -867 2897 -833
rect 2863 -935 2897 -901
rect 2863 -1004 2897 -969
rect 2959 969 2993 1004
rect 2959 901 2993 935
rect 2959 833 2993 867
rect 2959 765 2993 799
rect 2959 697 2993 731
rect 2959 629 2993 663
rect 2959 561 2993 595
rect 2959 493 2993 527
rect 2959 425 2993 459
rect 2959 357 2993 391
rect 2959 289 2993 323
rect 2959 221 2993 255
rect 2959 153 2993 187
rect 2959 85 2993 119
rect 2959 17 2993 51
rect 2959 -51 2993 -17
rect 2959 -119 2993 -85
rect 2959 -187 2993 -153
rect 2959 -255 2993 -221
rect 2959 -323 2993 -289
rect 2959 -391 2993 -357
rect 2959 -459 2993 -425
rect 2959 -527 2993 -493
rect 2959 -595 2993 -561
rect 2959 -663 2993 -629
rect 2959 -731 2993 -697
rect 2959 -799 2993 -765
rect 2959 -867 2993 -833
rect 2959 -935 2993 -901
rect 2959 -1004 2993 -969
rect 3055 969 3089 1004
rect 3055 901 3089 935
rect 3055 833 3089 867
rect 3055 765 3089 799
rect 3055 697 3089 731
rect 3055 629 3089 663
rect 3055 561 3089 595
rect 3055 493 3089 527
rect 3055 425 3089 459
rect 3055 357 3089 391
rect 3055 289 3089 323
rect 3055 221 3089 255
rect 3055 153 3089 187
rect 3055 85 3089 119
rect 3055 17 3089 51
rect 3055 -51 3089 -17
rect 3055 -119 3089 -85
rect 3055 -187 3089 -153
rect 3055 -255 3089 -221
rect 3055 -323 3089 -289
rect 3055 -391 3089 -357
rect 3055 -459 3089 -425
rect 3055 -527 3089 -493
rect 3055 -595 3089 -561
rect 3055 -663 3089 -629
rect 3055 -731 3089 -697
rect 3055 -799 3089 -765
rect 3055 -867 3089 -833
rect 3055 -935 3089 -901
rect 3055 -1004 3089 -969
rect 3151 969 3185 1004
rect 3151 901 3185 935
rect 3151 833 3185 867
rect 3151 765 3185 799
rect 3151 697 3185 731
rect 3151 629 3185 663
rect 3151 561 3185 595
rect 3151 493 3185 527
rect 3151 425 3185 459
rect 3151 357 3185 391
rect 3151 289 3185 323
rect 3151 221 3185 255
rect 3151 153 3185 187
rect 3151 85 3185 119
rect 3151 17 3185 51
rect 3151 -51 3185 -17
rect 3151 -119 3185 -85
rect 3151 -187 3185 -153
rect 3151 -255 3185 -221
rect 3151 -323 3185 -289
rect 3151 -391 3185 -357
rect 3151 -459 3185 -425
rect 3151 -527 3185 -493
rect 3151 -595 3185 -561
rect 3151 -663 3185 -629
rect 3151 -731 3185 -697
rect 3151 -799 3185 -765
rect 3151 -867 3185 -833
rect 3151 -935 3185 -901
rect 3151 -1004 3185 -969
rect 3247 969 3281 1004
rect 3247 901 3281 935
rect 3247 833 3281 867
rect 3247 765 3281 799
rect 3247 697 3281 731
rect 3247 629 3281 663
rect 3247 561 3281 595
rect 3247 493 3281 527
rect 3247 425 3281 459
rect 3247 357 3281 391
rect 3247 289 3281 323
rect 3247 221 3281 255
rect 3247 153 3281 187
rect 3247 85 3281 119
rect 3247 17 3281 51
rect 3247 -51 3281 -17
rect 3247 -119 3281 -85
rect 3247 -187 3281 -153
rect 3247 -255 3281 -221
rect 3247 -323 3281 -289
rect 3247 -391 3281 -357
rect 3247 -459 3281 -425
rect 3247 -527 3281 -493
rect 3247 -595 3281 -561
rect 3247 -663 3281 -629
rect 3247 -731 3281 -697
rect 3247 -799 3281 -765
rect 3247 -867 3281 -833
rect 3247 -935 3281 -901
rect 3247 -1004 3281 -969
rect 3343 969 3377 1004
rect 3343 901 3377 935
rect 3343 833 3377 867
rect 3343 765 3377 799
rect 3343 697 3377 731
rect 3343 629 3377 663
rect 3343 561 3377 595
rect 3343 493 3377 527
rect 3343 425 3377 459
rect 3343 357 3377 391
rect 3343 289 3377 323
rect 3343 221 3377 255
rect 3343 153 3377 187
rect 3343 85 3377 119
rect 3343 17 3377 51
rect 3343 -51 3377 -17
rect 3343 -119 3377 -85
rect 3343 -187 3377 -153
rect 3343 -255 3377 -221
rect 3343 -323 3377 -289
rect 3343 -391 3377 -357
rect 3343 -459 3377 -425
rect 3343 -527 3377 -493
rect 3343 -595 3377 -561
rect 3343 -663 3377 -629
rect 3343 -731 3377 -697
rect 3343 -799 3377 -765
rect 3343 -867 3377 -833
rect 3343 -935 3377 -901
rect 3343 -1004 3377 -969
rect 3439 969 3473 1004
rect 3439 901 3473 935
rect 3439 833 3473 867
rect 3439 765 3473 799
rect 3439 697 3473 731
rect 3439 629 3473 663
rect 3439 561 3473 595
rect 3439 493 3473 527
rect 3439 425 3473 459
rect 3439 357 3473 391
rect 3439 289 3473 323
rect 3439 221 3473 255
rect 3439 153 3473 187
rect 3439 85 3473 119
rect 3439 17 3473 51
rect 3439 -51 3473 -17
rect 3439 -119 3473 -85
rect 3439 -187 3473 -153
rect 3439 -255 3473 -221
rect 3439 -323 3473 -289
rect 3439 -391 3473 -357
rect 3439 -459 3473 -425
rect 3439 -527 3473 -493
rect 3439 -595 3473 -561
rect 3439 -663 3473 -629
rect 3439 -731 3473 -697
rect 3439 -799 3473 -765
rect 3439 -867 3473 -833
rect 3439 -935 3473 -901
rect 3439 -1004 3473 -969
rect 3535 969 3569 1004
rect 3535 901 3569 935
rect 3535 833 3569 867
rect 3535 765 3569 799
rect 3535 697 3569 731
rect 3535 629 3569 663
rect 3535 561 3569 595
rect 3535 493 3569 527
rect 3535 425 3569 459
rect 3535 357 3569 391
rect 3535 289 3569 323
rect 3535 221 3569 255
rect 3535 153 3569 187
rect 3535 85 3569 119
rect 3535 17 3569 51
rect 3535 -51 3569 -17
rect 3535 -119 3569 -85
rect 3535 -187 3569 -153
rect 3535 -255 3569 -221
rect 3535 -323 3569 -289
rect 3535 -391 3569 -357
rect 3535 -459 3569 -425
rect 3535 -527 3569 -493
rect 3535 -595 3569 -561
rect 3535 -663 3569 -629
rect 3535 -731 3569 -697
rect 3535 -799 3569 -765
rect 3535 -867 3569 -833
rect 3535 -935 3569 -901
rect 3535 -1004 3569 -969
rect 3631 969 3665 1004
rect 3631 901 3665 935
rect 3631 833 3665 867
rect 3631 765 3665 799
rect 3631 697 3665 731
rect 3631 629 3665 663
rect 3631 561 3665 595
rect 3631 493 3665 527
rect 3631 425 3665 459
rect 3631 357 3665 391
rect 3631 289 3665 323
rect 3631 221 3665 255
rect 3631 153 3665 187
rect 3631 85 3665 119
rect 3631 17 3665 51
rect 3631 -51 3665 -17
rect 3631 -119 3665 -85
rect 3631 -187 3665 -153
rect 3631 -255 3665 -221
rect 3631 -323 3665 -289
rect 3631 -391 3665 -357
rect 3631 -459 3665 -425
rect 3631 -527 3665 -493
rect 3631 -595 3665 -561
rect 3631 -663 3665 -629
rect 3631 -731 3665 -697
rect 3631 -799 3665 -765
rect 3631 -867 3665 -833
rect 3631 -935 3665 -901
rect 3631 -1004 3665 -969
rect 3727 969 3761 1004
rect 3727 901 3761 935
rect 3727 833 3761 867
rect 3727 765 3761 799
rect 3727 697 3761 731
rect 3727 629 3761 663
rect 3727 561 3761 595
rect 3727 493 3761 527
rect 3727 425 3761 459
rect 3727 357 3761 391
rect 3727 289 3761 323
rect 3727 221 3761 255
rect 3727 153 3761 187
rect 3727 85 3761 119
rect 3727 17 3761 51
rect 3727 -51 3761 -17
rect 3727 -119 3761 -85
rect 3727 -187 3761 -153
rect 3727 -255 3761 -221
rect 3727 -323 3761 -289
rect 3727 -391 3761 -357
rect 3727 -459 3761 -425
rect 3727 -527 3761 -493
rect 3727 -595 3761 -561
rect 3727 -663 3761 -629
rect 3727 -731 3761 -697
rect 3727 -799 3761 -765
rect 3727 -867 3761 -833
rect 3727 -935 3761 -901
rect 3727 -1004 3761 -969
rect 3823 969 3857 1004
rect 3823 901 3857 935
rect 3823 833 3857 867
rect 3823 765 3857 799
rect 3823 697 3857 731
rect 3823 629 3857 663
rect 3823 561 3857 595
rect 3823 493 3857 527
rect 3823 425 3857 459
rect 3823 357 3857 391
rect 3823 289 3857 323
rect 3823 221 3857 255
rect 3823 153 3857 187
rect 3823 85 3857 119
rect 3823 17 3857 51
rect 3823 -51 3857 -17
rect 3823 -119 3857 -85
rect 3823 -187 3857 -153
rect 3823 -255 3857 -221
rect 3823 -323 3857 -289
rect 3823 -391 3857 -357
rect 3823 -459 3857 -425
rect 3823 -527 3857 -493
rect 3823 -595 3857 -561
rect 3823 -663 3857 -629
rect 3823 -731 3857 -697
rect 3823 -799 3857 -765
rect 3823 -867 3857 -833
rect 3823 -935 3857 -901
rect 3823 -1004 3857 -969
rect 3919 969 3953 1004
rect 3919 901 3953 935
rect 3919 833 3953 867
rect 3919 765 3953 799
rect 3919 697 3953 731
rect 3919 629 3953 663
rect 3919 561 3953 595
rect 3919 493 3953 527
rect 3919 425 3953 459
rect 3919 357 3953 391
rect 3919 289 3953 323
rect 3919 221 3953 255
rect 3919 153 3953 187
rect 3919 85 3953 119
rect 3919 17 3953 51
rect 3919 -51 3953 -17
rect 3919 -119 3953 -85
rect 3919 -187 3953 -153
rect 3919 -255 3953 -221
rect 3919 -323 3953 -289
rect 3919 -391 3953 -357
rect 3919 -459 3953 -425
rect 3919 -527 3953 -493
rect 3919 -595 3953 -561
rect 3919 -663 3953 -629
rect 3919 -731 3953 -697
rect 3919 -799 3953 -765
rect 3919 -867 3953 -833
rect 3919 -935 3953 -901
rect 3919 -1004 3953 -969
rect 4015 969 4049 1004
rect 4015 901 4049 935
rect 4015 833 4049 867
rect 4015 765 4049 799
rect 4015 697 4049 731
rect 4015 629 4049 663
rect 4015 561 4049 595
rect 4015 493 4049 527
rect 4015 425 4049 459
rect 4015 357 4049 391
rect 4015 289 4049 323
rect 4015 221 4049 255
rect 4015 153 4049 187
rect 4015 85 4049 119
rect 4015 17 4049 51
rect 4015 -51 4049 -17
rect 4015 -119 4049 -85
rect 4015 -187 4049 -153
rect 4015 -255 4049 -221
rect 4015 -323 4049 -289
rect 4015 -391 4049 -357
rect 4015 -459 4049 -425
rect 4015 -527 4049 -493
rect 4015 -595 4049 -561
rect 4015 -663 4049 -629
rect 4015 -731 4049 -697
rect 4015 -799 4049 -765
rect 4015 -867 4049 -833
rect 4015 -935 4049 -901
rect 4015 -1004 4049 -969
rect 4111 969 4145 1004
rect 4111 901 4145 935
rect 4111 833 4145 867
rect 4111 765 4145 799
rect 4111 697 4145 731
rect 4111 629 4145 663
rect 4111 561 4145 595
rect 4111 493 4145 527
rect 4111 425 4145 459
rect 4111 357 4145 391
rect 4111 289 4145 323
rect 4111 221 4145 255
rect 4111 153 4145 187
rect 4111 85 4145 119
rect 4111 17 4145 51
rect 4111 -51 4145 -17
rect 4111 -119 4145 -85
rect 4111 -187 4145 -153
rect 4111 -255 4145 -221
rect 4111 -323 4145 -289
rect 4111 -391 4145 -357
rect 4111 -459 4145 -425
rect 4111 -527 4145 -493
rect 4111 -595 4145 -561
rect 4111 -663 4145 -629
rect 4111 -731 4145 -697
rect 4111 -799 4145 -765
rect 4111 -867 4145 -833
rect 4111 -935 4145 -901
rect 4111 -1004 4145 -969
rect 4207 969 4241 1004
rect 4207 901 4241 935
rect 4207 833 4241 867
rect 4207 765 4241 799
rect 4207 697 4241 731
rect 4207 629 4241 663
rect 4207 561 4241 595
rect 4207 493 4241 527
rect 4207 425 4241 459
rect 4207 357 4241 391
rect 4207 289 4241 323
rect 4207 221 4241 255
rect 4207 153 4241 187
rect 4207 85 4241 119
rect 4207 17 4241 51
rect 4207 -51 4241 -17
rect 4207 -119 4241 -85
rect 4207 -187 4241 -153
rect 4207 -255 4241 -221
rect 4207 -323 4241 -289
rect 4207 -391 4241 -357
rect 4207 -459 4241 -425
rect 4207 -527 4241 -493
rect 4207 -595 4241 -561
rect 4207 -663 4241 -629
rect 4207 -731 4241 -697
rect 4207 -799 4241 -765
rect 4207 -867 4241 -833
rect 4207 -935 4241 -901
rect 4207 -1004 4241 -969
rect 4303 969 4337 1004
rect 4303 901 4337 935
rect 4303 833 4337 867
rect 4303 765 4337 799
rect 4303 697 4337 731
rect 4303 629 4337 663
rect 4303 561 4337 595
rect 4303 493 4337 527
rect 4303 425 4337 459
rect 4303 357 4337 391
rect 4303 289 4337 323
rect 4303 221 4337 255
rect 4303 153 4337 187
rect 4303 85 4337 119
rect 4303 17 4337 51
rect 4303 -51 4337 -17
rect 4303 -119 4337 -85
rect 4303 -187 4337 -153
rect 4303 -255 4337 -221
rect 4303 -323 4337 -289
rect 4303 -391 4337 -357
rect 4303 -459 4337 -425
rect 4303 -527 4337 -493
rect 4303 -595 4337 -561
rect 4303 -663 4337 -629
rect 4303 -731 4337 -697
rect 4303 -799 4337 -765
rect 4303 -867 4337 -833
rect 4303 -935 4337 -901
rect 4303 -1004 4337 -969
rect 4399 969 4433 1004
rect 4399 901 4433 935
rect 4399 833 4433 867
rect 4399 765 4433 799
rect 4399 697 4433 731
rect 4399 629 4433 663
rect 4399 561 4433 595
rect 4399 493 4433 527
rect 4399 425 4433 459
rect 4399 357 4433 391
rect 4399 289 4433 323
rect 4399 221 4433 255
rect 4399 153 4433 187
rect 4399 85 4433 119
rect 4399 17 4433 51
rect 4399 -51 4433 -17
rect 4399 -119 4433 -85
rect 4399 -187 4433 -153
rect 4399 -255 4433 -221
rect 4399 -323 4433 -289
rect 4399 -391 4433 -357
rect 4399 -459 4433 -425
rect 4399 -527 4433 -493
rect 4399 -595 4433 -561
rect 4399 -663 4433 -629
rect 4399 -731 4433 -697
rect 4399 -799 4433 -765
rect 4399 -867 4433 -833
rect 4399 -935 4433 -901
rect 4399 -1004 4433 -969
rect 4495 969 4529 1004
rect 4495 901 4529 935
rect 4495 833 4529 867
rect 4495 765 4529 799
rect 4495 697 4529 731
rect 4495 629 4529 663
rect 4495 561 4529 595
rect 4495 493 4529 527
rect 4495 425 4529 459
rect 4495 357 4529 391
rect 4495 289 4529 323
rect 4495 221 4529 255
rect 4495 153 4529 187
rect 4495 85 4529 119
rect 4495 17 4529 51
rect 4495 -51 4529 -17
rect 4495 -119 4529 -85
rect 4495 -187 4529 -153
rect 4495 -255 4529 -221
rect 4495 -323 4529 -289
rect 4495 -391 4529 -357
rect 4495 -459 4529 -425
rect 4495 -527 4529 -493
rect 4495 -595 4529 -561
rect 4495 -663 4529 -629
rect 4495 -731 4529 -697
rect 4495 -799 4529 -765
rect 4495 -867 4529 -833
rect 4495 -935 4529 -901
rect 4495 -1004 4529 -969
rect 4591 969 4625 1004
rect 4591 901 4625 935
rect 4591 833 4625 867
rect 4591 765 4625 799
rect 4591 697 4625 731
rect 4591 629 4625 663
rect 4591 561 4625 595
rect 4591 493 4625 527
rect 4591 425 4625 459
rect 4591 357 4625 391
rect 4591 289 4625 323
rect 4591 221 4625 255
rect 4591 153 4625 187
rect 4591 85 4625 119
rect 4591 17 4625 51
rect 4591 -51 4625 -17
rect 4591 -119 4625 -85
rect 4591 -187 4625 -153
rect 4591 -255 4625 -221
rect 4591 -323 4625 -289
rect 4591 -391 4625 -357
rect 4591 -459 4625 -425
rect 4591 -527 4625 -493
rect 4591 -595 4625 -561
rect 4591 -663 4625 -629
rect 4591 -731 4625 -697
rect 4591 -799 4625 -765
rect 4591 -867 4625 -833
rect 4591 -935 4625 -901
rect 4591 -1004 4625 -969
rect 4687 969 4721 1004
rect 4687 901 4721 935
rect 4687 833 4721 867
rect 4687 765 4721 799
rect 4687 697 4721 731
rect 4687 629 4721 663
rect 4687 561 4721 595
rect 4687 493 4721 527
rect 4687 425 4721 459
rect 4687 357 4721 391
rect 4687 289 4721 323
rect 4687 221 4721 255
rect 4687 153 4721 187
rect 4687 85 4721 119
rect 4687 17 4721 51
rect 4687 -51 4721 -17
rect 4687 -119 4721 -85
rect 4687 -187 4721 -153
rect 4687 -255 4721 -221
rect 4687 -323 4721 -289
rect 4687 -391 4721 -357
rect 4687 -459 4721 -425
rect 4687 -527 4721 -493
rect 4687 -595 4721 -561
rect 4687 -663 4721 -629
rect 4687 -731 4721 -697
rect 4687 -799 4721 -765
rect 4687 -867 4721 -833
rect 4687 -935 4721 -901
rect 4687 -1004 4721 -969
rect 4783 969 4817 1004
rect 4783 901 4817 935
rect 4783 833 4817 867
rect 4783 765 4817 799
rect 4783 697 4817 731
rect 4783 629 4817 663
rect 4783 561 4817 595
rect 4783 493 4817 527
rect 4783 425 4817 459
rect 4783 357 4817 391
rect 4783 289 4817 323
rect 4783 221 4817 255
rect 4783 153 4817 187
rect 4783 85 4817 119
rect 4783 17 4817 51
rect 4783 -51 4817 -17
rect 4783 -119 4817 -85
rect 4783 -187 4817 -153
rect 4783 -255 4817 -221
rect 4783 -323 4817 -289
rect 4783 -391 4817 -357
rect 4783 -459 4817 -425
rect 4783 -527 4817 -493
rect 4783 -595 4817 -561
rect 4783 -663 4817 -629
rect 4783 -731 4817 -697
rect 4783 -799 4817 -765
rect 4783 -867 4817 -833
rect 4783 -935 4817 -901
rect 4783 -1004 4817 -969
rect 4897 1003 4931 1037
rect 4897 935 4931 969
rect 4897 867 4931 901
rect 4897 799 4931 833
rect 4897 731 4931 765
rect 4897 663 4931 697
rect 4897 595 4931 629
rect 4897 527 4931 561
rect 4897 459 4931 493
rect 4897 391 4931 425
rect 4897 323 4931 357
rect 4897 255 4931 289
rect 4897 187 4931 221
rect 4897 119 4931 153
rect 4897 51 4931 85
rect 4897 -17 4931 17
rect 4897 -85 4931 -51
rect 4897 -153 4931 -119
rect 4897 -221 4931 -187
rect 4897 -289 4931 -255
rect 4897 -357 4931 -323
rect 4897 -425 4931 -391
rect 4897 -493 4931 -459
rect 4897 -561 4931 -527
rect 4897 -629 4931 -595
rect 4897 -697 4931 -663
rect 4897 -765 4931 -731
rect 4897 -833 4931 -799
rect 4897 -901 4931 -867
rect 4897 -969 4931 -935
rect 4897 -1037 4931 -1003
rect -4931 -1140 -4897 -1071
rect -4785 -1072 -4769 -1038
rect -4735 -1072 -4719 -1038
rect -4593 -1072 -4577 -1038
rect -4543 -1072 -4527 -1038
rect -4401 -1072 -4385 -1038
rect -4351 -1072 -4335 -1038
rect -4209 -1072 -4193 -1038
rect -4159 -1072 -4143 -1038
rect -4017 -1072 -4001 -1038
rect -3967 -1072 -3951 -1038
rect -3825 -1072 -3809 -1038
rect -3775 -1072 -3759 -1038
rect -3633 -1072 -3617 -1038
rect -3583 -1072 -3567 -1038
rect -3441 -1072 -3425 -1038
rect -3391 -1072 -3375 -1038
rect -3249 -1072 -3233 -1038
rect -3199 -1072 -3183 -1038
rect -3057 -1072 -3041 -1038
rect -3007 -1072 -2991 -1038
rect -2865 -1072 -2849 -1038
rect -2815 -1072 -2799 -1038
rect -2673 -1072 -2657 -1038
rect -2623 -1072 -2607 -1038
rect -2481 -1072 -2465 -1038
rect -2431 -1072 -2415 -1038
rect -2289 -1072 -2273 -1038
rect -2239 -1072 -2223 -1038
rect -2097 -1072 -2081 -1038
rect -2047 -1072 -2031 -1038
rect -1905 -1072 -1889 -1038
rect -1855 -1072 -1839 -1038
rect -1713 -1072 -1697 -1038
rect -1663 -1072 -1647 -1038
rect -1521 -1072 -1505 -1038
rect -1471 -1072 -1455 -1038
rect -1329 -1072 -1313 -1038
rect -1279 -1072 -1263 -1038
rect -1137 -1072 -1121 -1038
rect -1087 -1072 -1071 -1038
rect -945 -1072 -929 -1038
rect -895 -1072 -879 -1038
rect -753 -1072 -737 -1038
rect -703 -1072 -687 -1038
rect -561 -1072 -545 -1038
rect -511 -1072 -495 -1038
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect 399 -1072 415 -1038
rect 449 -1072 465 -1038
rect 591 -1072 607 -1038
rect 641 -1072 657 -1038
rect 783 -1072 799 -1038
rect 833 -1072 849 -1038
rect 975 -1072 991 -1038
rect 1025 -1072 1041 -1038
rect 1167 -1072 1183 -1038
rect 1217 -1072 1233 -1038
rect 1359 -1072 1375 -1038
rect 1409 -1072 1425 -1038
rect 1551 -1072 1567 -1038
rect 1601 -1072 1617 -1038
rect 1743 -1072 1759 -1038
rect 1793 -1072 1809 -1038
rect 1935 -1072 1951 -1038
rect 1985 -1072 2001 -1038
rect 2127 -1072 2143 -1038
rect 2177 -1072 2193 -1038
rect 2319 -1072 2335 -1038
rect 2369 -1072 2385 -1038
rect 2511 -1072 2527 -1038
rect 2561 -1072 2577 -1038
rect 2703 -1072 2719 -1038
rect 2753 -1072 2769 -1038
rect 2895 -1072 2911 -1038
rect 2945 -1072 2961 -1038
rect 3087 -1072 3103 -1038
rect 3137 -1072 3153 -1038
rect 3279 -1072 3295 -1038
rect 3329 -1072 3345 -1038
rect 3471 -1072 3487 -1038
rect 3521 -1072 3537 -1038
rect 3663 -1072 3679 -1038
rect 3713 -1072 3729 -1038
rect 3855 -1072 3871 -1038
rect 3905 -1072 3921 -1038
rect 4047 -1072 4063 -1038
rect 4097 -1072 4113 -1038
rect 4239 -1072 4255 -1038
rect 4289 -1072 4305 -1038
rect 4431 -1072 4447 -1038
rect 4481 -1072 4497 -1038
rect 4623 -1072 4639 -1038
rect 4673 -1072 4689 -1038
rect 4897 -1140 4931 -1071
rect -4931 -1174 -4811 -1140
rect -4777 -1174 -4743 -1140
rect -4709 -1174 -4675 -1140
rect -4641 -1174 -4607 -1140
rect -4573 -1174 -4539 -1140
rect -4505 -1174 -4471 -1140
rect -4437 -1174 -4403 -1140
rect -4369 -1174 -4335 -1140
rect -4301 -1174 -4267 -1140
rect -4233 -1174 -4199 -1140
rect -4165 -1174 -4131 -1140
rect -4097 -1174 -4063 -1140
rect -4029 -1174 -3995 -1140
rect -3961 -1174 -3927 -1140
rect -3893 -1174 -3859 -1140
rect -3825 -1174 -3791 -1140
rect -3757 -1174 -3723 -1140
rect -3689 -1174 -3655 -1140
rect -3621 -1174 -3587 -1140
rect -3553 -1174 -3519 -1140
rect -3485 -1174 -3451 -1140
rect -3417 -1174 -3383 -1140
rect -3349 -1174 -3315 -1140
rect -3281 -1174 -3247 -1140
rect -3213 -1174 -3179 -1140
rect -3145 -1174 -3111 -1140
rect -3077 -1174 -3043 -1140
rect -3009 -1174 -2975 -1140
rect -2941 -1174 -2907 -1140
rect -2873 -1174 -2839 -1140
rect -2805 -1174 -2771 -1140
rect -2737 -1174 -2703 -1140
rect -2669 -1174 -2635 -1140
rect -2601 -1174 -2567 -1140
rect -2533 -1174 -2499 -1140
rect -2465 -1174 -2431 -1140
rect -2397 -1174 -2363 -1140
rect -2329 -1174 -2295 -1140
rect -2261 -1174 -2227 -1140
rect -2193 -1174 -2159 -1140
rect -2125 -1174 -2091 -1140
rect -2057 -1174 -2023 -1140
rect -1989 -1174 -1955 -1140
rect -1921 -1174 -1887 -1140
rect -1853 -1174 -1819 -1140
rect -1785 -1174 -1751 -1140
rect -1717 -1174 -1683 -1140
rect -1649 -1174 -1615 -1140
rect -1581 -1174 -1547 -1140
rect -1513 -1174 -1479 -1140
rect -1445 -1174 -1411 -1140
rect -1377 -1174 -1343 -1140
rect -1309 -1174 -1275 -1140
rect -1241 -1174 -1207 -1140
rect -1173 -1174 -1139 -1140
rect -1105 -1174 -1071 -1140
rect -1037 -1174 -1003 -1140
rect -969 -1174 -935 -1140
rect -901 -1174 -867 -1140
rect -833 -1174 -799 -1140
rect -765 -1174 -731 -1140
rect -697 -1174 -663 -1140
rect -629 -1174 -595 -1140
rect -561 -1174 -527 -1140
rect -493 -1174 -459 -1140
rect -425 -1174 -391 -1140
rect -357 -1174 -323 -1140
rect -289 -1174 -255 -1140
rect -221 -1174 -187 -1140
rect -153 -1174 -119 -1140
rect -85 -1174 -51 -1140
rect -17 -1174 17 -1140
rect 51 -1174 85 -1140
rect 119 -1174 153 -1140
rect 187 -1174 221 -1140
rect 255 -1174 289 -1140
rect 323 -1174 357 -1140
rect 391 -1174 425 -1140
rect 459 -1174 493 -1140
rect 527 -1174 561 -1140
rect 595 -1174 629 -1140
rect 663 -1174 697 -1140
rect 731 -1174 765 -1140
rect 799 -1174 833 -1140
rect 867 -1174 901 -1140
rect 935 -1174 969 -1140
rect 1003 -1174 1037 -1140
rect 1071 -1174 1105 -1140
rect 1139 -1174 1173 -1140
rect 1207 -1174 1241 -1140
rect 1275 -1174 1309 -1140
rect 1343 -1174 1377 -1140
rect 1411 -1174 1445 -1140
rect 1479 -1174 1513 -1140
rect 1547 -1174 1581 -1140
rect 1615 -1174 1649 -1140
rect 1683 -1174 1717 -1140
rect 1751 -1174 1785 -1140
rect 1819 -1174 1853 -1140
rect 1887 -1174 1921 -1140
rect 1955 -1174 1989 -1140
rect 2023 -1174 2057 -1140
rect 2091 -1174 2125 -1140
rect 2159 -1174 2193 -1140
rect 2227 -1174 2261 -1140
rect 2295 -1174 2329 -1140
rect 2363 -1174 2397 -1140
rect 2431 -1174 2465 -1140
rect 2499 -1174 2533 -1140
rect 2567 -1174 2601 -1140
rect 2635 -1174 2669 -1140
rect 2703 -1174 2737 -1140
rect 2771 -1174 2805 -1140
rect 2839 -1174 2873 -1140
rect 2907 -1174 2941 -1140
rect 2975 -1174 3009 -1140
rect 3043 -1174 3077 -1140
rect 3111 -1174 3145 -1140
rect 3179 -1174 3213 -1140
rect 3247 -1174 3281 -1140
rect 3315 -1174 3349 -1140
rect 3383 -1174 3417 -1140
rect 3451 -1174 3485 -1140
rect 3519 -1174 3553 -1140
rect 3587 -1174 3621 -1140
rect 3655 -1174 3689 -1140
rect 3723 -1174 3757 -1140
rect 3791 -1174 3825 -1140
rect 3859 -1174 3893 -1140
rect 3927 -1174 3961 -1140
rect 3995 -1174 4029 -1140
rect 4063 -1174 4097 -1140
rect 4131 -1174 4165 -1140
rect 4199 -1174 4233 -1140
rect 4267 -1174 4301 -1140
rect 4335 -1174 4369 -1140
rect 4403 -1174 4437 -1140
rect 4471 -1174 4505 -1140
rect 4539 -1174 4573 -1140
rect 4607 -1174 4641 -1140
rect 4675 -1174 4709 -1140
rect 4743 -1174 4777 -1140
rect 4811 -1174 4931 -1140
<< properties >>
string FIXED_BBOX -4914 -1157 4914 1157
<< end >>
