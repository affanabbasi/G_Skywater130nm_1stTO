magic
tech sky130A
timestamp 1606471058
<< nwell >>
rect -885 -459 885 459
<< pmos >>
rect -787 -350 -587 350
rect -558 -350 -358 350
rect -329 -350 -129 350
rect -100 -350 100 350
rect 129 -350 329 350
rect 358 -350 558 350
rect 587 -350 787 350
<< pdiff >>
rect -816 344 -787 350
rect -816 -344 -810 344
rect -793 -344 -787 344
rect -816 -350 -787 -344
rect -587 344 -558 350
rect -587 -344 -581 344
rect -564 -344 -558 344
rect -587 -350 -558 -344
rect -358 344 -329 350
rect -358 -344 -352 344
rect -335 -344 -329 344
rect -358 -350 -329 -344
rect -129 344 -100 350
rect -129 -344 -123 344
rect -106 -344 -100 344
rect -129 -350 -100 -344
rect 100 344 129 350
rect 100 -344 106 344
rect 123 -344 129 344
rect 100 -350 129 -344
rect 329 344 358 350
rect 329 -344 335 344
rect 352 -344 358 344
rect 329 -350 358 -344
rect 558 344 587 350
rect 558 -344 564 344
rect 581 -344 587 344
rect 558 -350 587 -344
rect 787 344 816 350
rect 787 -344 793 344
rect 810 -344 816 344
rect 787 -350 816 -344
<< pdiffc >>
rect -810 -344 -793 344
rect -581 -344 -564 344
rect -352 -344 -335 344
rect -123 -344 -106 344
rect 106 -344 123 344
rect 335 -344 352 344
rect 564 -344 581 344
rect 793 -344 810 344
<< nsubdiff >>
rect -867 424 -819 441
rect 819 424 867 441
rect -867 393 -850 424
rect 850 393 867 424
rect -867 -424 -850 -393
rect 850 -424 867 -393
rect -867 -441 -819 -424
rect 819 -441 867 -424
<< nsubdiffcont >>
rect -819 424 819 441
rect -867 -393 -850 393
rect 850 -393 867 393
rect -819 -441 819 -424
<< poly >>
rect -787 390 -587 398
rect -787 373 -779 390
rect -595 373 -587 390
rect -787 350 -587 373
rect -558 390 -358 398
rect -558 373 -550 390
rect -366 373 -358 390
rect -558 350 -358 373
rect -329 390 -129 398
rect -329 373 -321 390
rect -137 373 -129 390
rect -329 350 -129 373
rect -100 390 100 398
rect -100 373 -92 390
rect 92 373 100 390
rect -100 350 100 373
rect 129 390 329 398
rect 129 373 137 390
rect 321 373 329 390
rect 129 350 329 373
rect 358 390 558 398
rect 358 373 366 390
rect 550 373 558 390
rect 358 350 558 373
rect 587 390 787 398
rect 587 373 595 390
rect 779 373 787 390
rect 587 350 787 373
rect -787 -373 -587 -350
rect -787 -390 -779 -373
rect -595 -390 -587 -373
rect -787 -398 -587 -390
rect -558 -373 -358 -350
rect -558 -390 -550 -373
rect -366 -390 -358 -373
rect -558 -398 -358 -390
rect -329 -373 -129 -350
rect -329 -390 -321 -373
rect -137 -390 -129 -373
rect -329 -398 -129 -390
rect -100 -373 100 -350
rect -100 -390 -92 -373
rect 92 -390 100 -373
rect -100 -398 100 -390
rect 129 -373 329 -350
rect 129 -390 137 -373
rect 321 -390 329 -373
rect 129 -398 329 -390
rect 358 -373 558 -350
rect 358 -390 366 -373
rect 550 -390 558 -373
rect 358 -398 558 -390
rect 587 -373 787 -350
rect 587 -390 595 -373
rect 779 -390 787 -373
rect 587 -398 787 -390
<< polycont >>
rect -779 373 -595 390
rect -550 373 -366 390
rect -321 373 -137 390
rect -92 373 92 390
rect 137 373 321 390
rect 366 373 550 390
rect 595 373 779 390
rect -779 -390 -595 -373
rect -550 -390 -366 -373
rect -321 -390 -137 -373
rect -92 -390 92 -373
rect 137 -390 321 -373
rect 366 -390 550 -373
rect 595 -390 779 -373
<< locali >>
rect -867 424 -819 441
rect 819 424 867 441
rect -867 393 -850 424
rect 850 393 867 424
rect -787 373 -779 390
rect -595 373 -587 390
rect -558 373 -550 390
rect -366 373 -358 390
rect -329 373 -321 390
rect -137 373 -129 390
rect -100 373 -92 390
rect 92 373 100 390
rect 129 373 137 390
rect 321 373 329 390
rect 358 373 366 390
rect 550 373 558 390
rect 587 373 595 390
rect 779 373 787 390
rect -810 344 -793 352
rect -810 -352 -793 -344
rect -581 344 -564 352
rect -581 -352 -564 -344
rect -352 344 -335 352
rect -352 -352 -335 -344
rect -123 344 -106 352
rect -123 -352 -106 -344
rect 106 344 123 352
rect 106 -352 123 -344
rect 335 344 352 352
rect 335 -352 352 -344
rect 564 344 581 352
rect 564 -352 581 -344
rect 793 344 810 352
rect 793 -352 810 -344
rect -787 -390 -779 -373
rect -595 -390 -587 -373
rect -558 -390 -550 -373
rect -366 -390 -358 -373
rect -329 -390 -321 -373
rect -137 -390 -129 -373
rect -100 -390 -92 -373
rect 92 -390 100 -373
rect 129 -390 137 -373
rect 321 -390 329 -373
rect 358 -390 366 -373
rect 550 -390 558 -373
rect 587 -390 595 -373
rect 779 -390 787 -373
rect -867 -424 -850 -393
rect 850 -424 867 -393
rect -867 -441 -819 -424
rect 819 -441 867 -424
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -858 -433 858 433
string parameters w 7 l 2 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
