magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -175 205 175 239
rect -175 -205 -141 205
rect 141 -205 175 205
rect -175 -239 175 -205
<< nmos >>
rect -15 -65 15 65
<< ndiff >>
rect -73 51 -15 65
rect -73 17 -61 51
rect -27 17 -15 51
rect -73 -17 -15 17
rect -73 -51 -61 -17
rect -27 -51 -15 -17
rect -73 -65 -15 -51
rect 15 51 73 65
rect 15 17 27 51
rect 61 17 73 51
rect 15 -17 73 17
rect 15 -51 27 -17
rect 61 -51 73 -17
rect 15 -65 73 -51
<< ndiffc >>
rect -61 17 -27 51
rect -61 -51 -27 -17
rect 27 17 61 51
rect 27 -51 61 -17
<< psubdiff >>
rect -175 205 -51 239
rect -17 205 17 239
rect 51 205 175 239
rect -175 119 -141 205
rect 141 119 175 205
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -205 -141 -119
rect 141 -205 175 -119
rect -175 -239 -51 -205
rect -17 -239 17 -205
rect 51 -239 175 -205
<< psubdiffcont >>
rect -51 205 -17 239
rect 17 205 51 239
rect -175 85 -141 119
rect 141 85 175 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -119 -141 -85
rect 141 -119 175 -85
rect -51 -239 -17 -205
rect 17 -239 51 -205
<< poly >>
rect -33 137 33 153
rect -33 103 -17 137
rect 17 103 33 137
rect -33 87 33 103
rect -15 65 15 87
rect -15 -87 15 -65
rect -33 -103 33 -87
rect -33 -137 -17 -103
rect 17 -137 33 -103
rect -33 -153 33 -137
<< polycont >>
rect -17 103 17 137
rect -17 -137 17 -103
<< locali >>
rect -175 205 -51 239
rect -17 205 17 239
rect 51 205 175 239
rect -175 119 -141 205
rect -33 103 -17 137
rect 17 103 33 137
rect 141 119 175 205
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -61 51 -27 69
rect -61 -17 -27 17
rect -61 -69 -27 -51
rect 27 51 61 69
rect 27 -17 61 17
rect 27 -69 61 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -205 -141 -119
rect -33 -137 -17 -103
rect 17 -137 33 -103
rect 141 -205 175 -119
rect -175 -239 -51 -205
rect -17 -239 17 -205
rect 51 -239 175 -205
<< properties >>
string FIXED_BBOX -158 -222 158 222
<< end >>
