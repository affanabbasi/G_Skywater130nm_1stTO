magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect -2166 -404 2166 404
<< nsubdiff >>
rect -2130 334 -2023 368
rect -1989 334 -1955 368
rect -1921 334 -1887 368
rect -1853 334 -1819 368
rect -1785 334 -1751 368
rect -1717 334 -1683 368
rect -1649 334 -1615 368
rect -1581 334 -1547 368
rect -1513 334 -1479 368
rect -1445 334 -1411 368
rect -1377 334 -1343 368
rect -1309 334 -1275 368
rect -1241 334 -1207 368
rect -1173 334 -1139 368
rect -1105 334 -1071 368
rect -1037 334 -1003 368
rect -969 334 -935 368
rect -901 334 -867 368
rect -833 334 -799 368
rect -765 334 -731 368
rect -697 334 -663 368
rect -629 334 -595 368
rect -561 334 -527 368
rect -493 334 -459 368
rect -425 334 -391 368
rect -357 334 -323 368
rect -289 334 -255 368
rect -221 334 -187 368
rect -153 334 -119 368
rect -85 334 -51 368
rect -17 334 17 368
rect 51 334 85 368
rect 119 334 153 368
rect 187 334 221 368
rect 255 334 289 368
rect 323 334 357 368
rect 391 334 425 368
rect 459 334 493 368
rect 527 334 561 368
rect 595 334 629 368
rect 663 334 697 368
rect 731 334 765 368
rect 799 334 833 368
rect 867 334 901 368
rect 935 334 969 368
rect 1003 334 1037 368
rect 1071 334 1105 368
rect 1139 334 1173 368
rect 1207 334 1241 368
rect 1275 334 1309 368
rect 1343 334 1377 368
rect 1411 334 1445 368
rect 1479 334 1513 368
rect 1547 334 1581 368
rect 1615 334 1649 368
rect 1683 334 1717 368
rect 1751 334 1785 368
rect 1819 334 1853 368
rect 1887 334 1921 368
rect 1955 334 1989 368
rect 2023 334 2130 368
rect -2130 255 -2096 334
rect 2096 255 2130 334
rect -2130 187 -2096 221
rect -2130 119 -2096 153
rect -2130 51 -2096 85
rect -2130 -17 -2096 17
rect -2130 -85 -2096 -51
rect -2130 -153 -2096 -119
rect -2130 -221 -2096 -187
rect 2096 187 2130 221
rect 2096 119 2130 153
rect 2096 51 2130 85
rect 2096 -17 2130 17
rect 2096 -85 2130 -51
rect 2096 -153 2130 -119
rect 2096 -221 2130 -187
rect -2130 -334 -2096 -255
rect 2096 -334 2130 -255
rect -2130 -368 -2023 -334
rect -1989 -368 -1955 -334
rect -1921 -368 -1887 -334
rect -1853 -368 -1819 -334
rect -1785 -368 -1751 -334
rect -1717 -368 -1683 -334
rect -1649 -368 -1615 -334
rect -1581 -368 -1547 -334
rect -1513 -368 -1479 -334
rect -1445 -368 -1411 -334
rect -1377 -368 -1343 -334
rect -1309 -368 -1275 -334
rect -1241 -368 -1207 -334
rect -1173 -368 -1139 -334
rect -1105 -368 -1071 -334
rect -1037 -368 -1003 -334
rect -969 -368 -935 -334
rect -901 -368 -867 -334
rect -833 -368 -799 -334
rect -765 -368 -731 -334
rect -697 -368 -663 -334
rect -629 -368 -595 -334
rect -561 -368 -527 -334
rect -493 -368 -459 -334
rect -425 -368 -391 -334
rect -357 -368 -323 -334
rect -289 -368 -255 -334
rect -221 -368 -187 -334
rect -153 -368 -119 -334
rect -85 -368 -51 -334
rect -17 -368 17 -334
rect 51 -368 85 -334
rect 119 -368 153 -334
rect 187 -368 221 -334
rect 255 -368 289 -334
rect 323 -368 357 -334
rect 391 -368 425 -334
rect 459 -368 493 -334
rect 527 -368 561 -334
rect 595 -368 629 -334
rect 663 -368 697 -334
rect 731 -368 765 -334
rect 799 -368 833 -334
rect 867 -368 901 -334
rect 935 -368 969 -334
rect 1003 -368 1037 -334
rect 1071 -368 1105 -334
rect 1139 -368 1173 -334
rect 1207 -368 1241 -334
rect 1275 -368 1309 -334
rect 1343 -368 1377 -334
rect 1411 -368 1445 -334
rect 1479 -368 1513 -334
rect 1547 -368 1581 -334
rect 1615 -368 1649 -334
rect 1683 -368 1717 -334
rect 1751 -368 1785 -334
rect 1819 -368 1853 -334
rect 1887 -368 1921 -334
rect 1955 -368 1989 -334
rect 2023 -368 2130 -334
<< nsubdiffcont >>
rect -2023 334 -1989 368
rect -1955 334 -1921 368
rect -1887 334 -1853 368
rect -1819 334 -1785 368
rect -1751 334 -1717 368
rect -1683 334 -1649 368
rect -1615 334 -1581 368
rect -1547 334 -1513 368
rect -1479 334 -1445 368
rect -1411 334 -1377 368
rect -1343 334 -1309 368
rect -1275 334 -1241 368
rect -1207 334 -1173 368
rect -1139 334 -1105 368
rect -1071 334 -1037 368
rect -1003 334 -969 368
rect -935 334 -901 368
rect -867 334 -833 368
rect -799 334 -765 368
rect -731 334 -697 368
rect -663 334 -629 368
rect -595 334 -561 368
rect -527 334 -493 368
rect -459 334 -425 368
rect -391 334 -357 368
rect -323 334 -289 368
rect -255 334 -221 368
rect -187 334 -153 368
rect -119 334 -85 368
rect -51 334 -17 368
rect 17 334 51 368
rect 85 334 119 368
rect 153 334 187 368
rect 221 334 255 368
rect 289 334 323 368
rect 357 334 391 368
rect 425 334 459 368
rect 493 334 527 368
rect 561 334 595 368
rect 629 334 663 368
rect 697 334 731 368
rect 765 334 799 368
rect 833 334 867 368
rect 901 334 935 368
rect 969 334 1003 368
rect 1037 334 1071 368
rect 1105 334 1139 368
rect 1173 334 1207 368
rect 1241 334 1275 368
rect 1309 334 1343 368
rect 1377 334 1411 368
rect 1445 334 1479 368
rect 1513 334 1547 368
rect 1581 334 1615 368
rect 1649 334 1683 368
rect 1717 334 1751 368
rect 1785 334 1819 368
rect 1853 334 1887 368
rect 1921 334 1955 368
rect 1989 334 2023 368
rect -2130 221 -2096 255
rect -2130 153 -2096 187
rect -2130 85 -2096 119
rect -2130 17 -2096 51
rect -2130 -51 -2096 -17
rect -2130 -119 -2096 -85
rect -2130 -187 -2096 -153
rect -2130 -255 -2096 -221
rect 2096 221 2130 255
rect 2096 153 2130 187
rect 2096 85 2130 119
rect 2096 17 2130 51
rect 2096 -51 2130 -17
rect 2096 -119 2130 -85
rect 2096 -187 2130 -153
rect 2096 -255 2130 -221
rect -2023 -368 -1989 -334
rect -1955 -368 -1921 -334
rect -1887 -368 -1853 -334
rect -1819 -368 -1785 -334
rect -1751 -368 -1717 -334
rect -1683 -368 -1649 -334
rect -1615 -368 -1581 -334
rect -1547 -368 -1513 -334
rect -1479 -368 -1445 -334
rect -1411 -368 -1377 -334
rect -1343 -368 -1309 -334
rect -1275 -368 -1241 -334
rect -1207 -368 -1173 -334
rect -1139 -368 -1105 -334
rect -1071 -368 -1037 -334
rect -1003 -368 -969 -334
rect -935 -368 -901 -334
rect -867 -368 -833 -334
rect -799 -368 -765 -334
rect -731 -368 -697 -334
rect -663 -368 -629 -334
rect -595 -368 -561 -334
rect -527 -368 -493 -334
rect -459 -368 -425 -334
rect -391 -368 -357 -334
rect -323 -368 -289 -334
rect -255 -368 -221 -334
rect -187 -368 -153 -334
rect -119 -368 -85 -334
rect -51 -368 -17 -334
rect 17 -368 51 -334
rect 85 -368 119 -334
rect 153 -368 187 -334
rect 221 -368 255 -334
rect 289 -368 323 -334
rect 357 -368 391 -334
rect 425 -368 459 -334
rect 493 -368 527 -334
rect 561 -368 595 -334
rect 629 -368 663 -334
rect 697 -368 731 -334
rect 765 -368 799 -334
rect 833 -368 867 -334
rect 901 -368 935 -334
rect 969 -368 1003 -334
rect 1037 -368 1071 -334
rect 1105 -368 1139 -334
rect 1173 -368 1207 -334
rect 1241 -368 1275 -334
rect 1309 -368 1343 -334
rect 1377 -368 1411 -334
rect 1445 -368 1479 -334
rect 1513 -368 1547 -334
rect 1581 -368 1615 -334
rect 1649 -368 1683 -334
rect 1717 -368 1751 -334
rect 1785 -368 1819 -334
rect 1853 -368 1887 -334
rect 1921 -368 1955 -334
rect 1989 -368 2023 -334
<< poly >>
rect -2000 222 2000 238
rect -2000 188 -1955 222
rect -1921 188 -1887 222
rect -1853 188 -1819 222
rect -1785 188 -1751 222
rect -1717 188 -1683 222
rect -1649 188 -1615 222
rect -1581 188 -1547 222
rect -1513 188 -1479 222
rect -1445 188 -1411 222
rect -1377 188 -1343 222
rect -1309 188 -1275 222
rect -1241 188 -1207 222
rect -1173 188 -1139 222
rect -1105 188 -1071 222
rect -1037 188 -1003 222
rect -969 188 -935 222
rect -901 188 -867 222
rect -833 188 -799 222
rect -765 188 -731 222
rect -697 188 -663 222
rect -629 188 -595 222
rect -561 188 -527 222
rect -493 188 -459 222
rect -425 188 -391 222
rect -357 188 -323 222
rect -289 188 -255 222
rect -221 188 -187 222
rect -153 188 -119 222
rect -85 188 -51 222
rect -17 188 17 222
rect 51 188 85 222
rect 119 188 153 222
rect 187 188 221 222
rect 255 188 289 222
rect 323 188 357 222
rect 391 188 425 222
rect 459 188 493 222
rect 527 188 561 222
rect 595 188 629 222
rect 663 188 697 222
rect 731 188 765 222
rect 799 188 833 222
rect 867 188 901 222
rect 935 188 969 222
rect 1003 188 1037 222
rect 1071 188 1105 222
rect 1139 188 1173 222
rect 1207 188 1241 222
rect 1275 188 1309 222
rect 1343 188 1377 222
rect 1411 188 1445 222
rect 1479 188 1513 222
rect 1547 188 1581 222
rect 1615 188 1649 222
rect 1683 188 1717 222
rect 1751 188 1785 222
rect 1819 188 1853 222
rect 1887 188 1921 222
rect 1955 188 2000 222
rect -2000 165 2000 188
rect -2000 -188 2000 -165
rect -2000 -222 -1955 -188
rect -1921 -222 -1887 -188
rect -1853 -222 -1819 -188
rect -1785 -222 -1751 -188
rect -1717 -222 -1683 -188
rect -1649 -222 -1615 -188
rect -1581 -222 -1547 -188
rect -1513 -222 -1479 -188
rect -1445 -222 -1411 -188
rect -1377 -222 -1343 -188
rect -1309 -222 -1275 -188
rect -1241 -222 -1207 -188
rect -1173 -222 -1139 -188
rect -1105 -222 -1071 -188
rect -1037 -222 -1003 -188
rect -969 -222 -935 -188
rect -901 -222 -867 -188
rect -833 -222 -799 -188
rect -765 -222 -731 -188
rect -697 -222 -663 -188
rect -629 -222 -595 -188
rect -561 -222 -527 -188
rect -493 -222 -459 -188
rect -425 -222 -391 -188
rect -357 -222 -323 -188
rect -289 -222 -255 -188
rect -221 -222 -187 -188
rect -153 -222 -119 -188
rect -85 -222 -51 -188
rect -17 -222 17 -188
rect 51 -222 85 -188
rect 119 -222 153 -188
rect 187 -222 221 -188
rect 255 -222 289 -188
rect 323 -222 357 -188
rect 391 -222 425 -188
rect 459 -222 493 -188
rect 527 -222 561 -188
rect 595 -222 629 -188
rect 663 -222 697 -188
rect 731 -222 765 -188
rect 799 -222 833 -188
rect 867 -222 901 -188
rect 935 -222 969 -188
rect 1003 -222 1037 -188
rect 1071 -222 1105 -188
rect 1139 -222 1173 -188
rect 1207 -222 1241 -188
rect 1275 -222 1309 -188
rect 1343 -222 1377 -188
rect 1411 -222 1445 -188
rect 1479 -222 1513 -188
rect 1547 -222 1581 -188
rect 1615 -222 1649 -188
rect 1683 -222 1717 -188
rect 1751 -222 1785 -188
rect 1819 -222 1853 -188
rect 1887 -222 1921 -188
rect 1955 -222 2000 -188
rect -2000 -238 2000 -222
<< polycont >>
rect -1955 188 -1921 222
rect -1887 188 -1853 222
rect -1819 188 -1785 222
rect -1751 188 -1717 222
rect -1683 188 -1649 222
rect -1615 188 -1581 222
rect -1547 188 -1513 222
rect -1479 188 -1445 222
rect -1411 188 -1377 222
rect -1343 188 -1309 222
rect -1275 188 -1241 222
rect -1207 188 -1173 222
rect -1139 188 -1105 222
rect -1071 188 -1037 222
rect -1003 188 -969 222
rect -935 188 -901 222
rect -867 188 -833 222
rect -799 188 -765 222
rect -731 188 -697 222
rect -663 188 -629 222
rect -595 188 -561 222
rect -527 188 -493 222
rect -459 188 -425 222
rect -391 188 -357 222
rect -323 188 -289 222
rect -255 188 -221 222
rect -187 188 -153 222
rect -119 188 -85 222
rect -51 188 -17 222
rect 17 188 51 222
rect 85 188 119 222
rect 153 188 187 222
rect 221 188 255 222
rect 289 188 323 222
rect 357 188 391 222
rect 425 188 459 222
rect 493 188 527 222
rect 561 188 595 222
rect 629 188 663 222
rect 697 188 731 222
rect 765 188 799 222
rect 833 188 867 222
rect 901 188 935 222
rect 969 188 1003 222
rect 1037 188 1071 222
rect 1105 188 1139 222
rect 1173 188 1207 222
rect 1241 188 1275 222
rect 1309 188 1343 222
rect 1377 188 1411 222
rect 1445 188 1479 222
rect 1513 188 1547 222
rect 1581 188 1615 222
rect 1649 188 1683 222
rect 1717 188 1751 222
rect 1785 188 1819 222
rect 1853 188 1887 222
rect 1921 188 1955 222
rect -1955 -222 -1921 -188
rect -1887 -222 -1853 -188
rect -1819 -222 -1785 -188
rect -1751 -222 -1717 -188
rect -1683 -222 -1649 -188
rect -1615 -222 -1581 -188
rect -1547 -222 -1513 -188
rect -1479 -222 -1445 -188
rect -1411 -222 -1377 -188
rect -1343 -222 -1309 -188
rect -1275 -222 -1241 -188
rect -1207 -222 -1173 -188
rect -1139 -222 -1105 -188
rect -1071 -222 -1037 -188
rect -1003 -222 -969 -188
rect -935 -222 -901 -188
rect -867 -222 -833 -188
rect -799 -222 -765 -188
rect -731 -222 -697 -188
rect -663 -222 -629 -188
rect -595 -222 -561 -188
rect -527 -222 -493 -188
rect -459 -222 -425 -188
rect -391 -222 -357 -188
rect -323 -222 -289 -188
rect -255 -222 -221 -188
rect -187 -222 -153 -188
rect -119 -222 -85 -188
rect -51 -222 -17 -188
rect 17 -222 51 -188
rect 85 -222 119 -188
rect 153 -222 187 -188
rect 221 -222 255 -188
rect 289 -222 323 -188
rect 357 -222 391 -188
rect 425 -222 459 -188
rect 493 -222 527 -188
rect 561 -222 595 -188
rect 629 -222 663 -188
rect 697 -222 731 -188
rect 765 -222 799 -188
rect 833 -222 867 -188
rect 901 -222 935 -188
rect 969 -222 1003 -188
rect 1037 -222 1071 -188
rect 1105 -222 1139 -188
rect 1173 -222 1207 -188
rect 1241 -222 1275 -188
rect 1309 -222 1343 -188
rect 1377 -222 1411 -188
rect 1445 -222 1479 -188
rect 1513 -222 1547 -188
rect 1581 -222 1615 -188
rect 1649 -222 1683 -188
rect 1717 -222 1751 -188
rect 1785 -222 1819 -188
rect 1853 -222 1887 -188
rect 1921 -222 1955 -188
<< npolyres >>
rect -2000 -165 2000 165
<< locali >>
rect -2130 334 -2023 368
rect -1989 334 -1955 368
rect -1921 334 -1887 368
rect -1853 334 -1819 368
rect -1785 334 -1751 368
rect -1717 334 -1683 368
rect -1649 334 -1615 368
rect -1581 334 -1547 368
rect -1513 334 -1479 368
rect -1445 334 -1411 368
rect -1377 334 -1343 368
rect -1309 334 -1275 368
rect -1241 334 -1207 368
rect -1173 334 -1139 368
rect -1105 334 -1071 368
rect -1037 334 -1003 368
rect -969 334 -935 368
rect -901 334 -867 368
rect -833 334 -799 368
rect -765 334 -731 368
rect -697 334 -663 368
rect -629 334 -595 368
rect -561 334 -527 368
rect -493 334 -459 368
rect -425 334 -391 368
rect -357 334 -323 368
rect -289 334 -255 368
rect -221 334 -187 368
rect -153 334 -119 368
rect -85 334 -51 368
rect -17 334 17 368
rect 51 334 85 368
rect 119 334 153 368
rect 187 334 221 368
rect 255 334 289 368
rect 323 334 357 368
rect 391 334 425 368
rect 459 334 493 368
rect 527 334 561 368
rect 595 334 629 368
rect 663 334 697 368
rect 731 334 765 368
rect 799 334 833 368
rect 867 334 901 368
rect 935 334 969 368
rect 1003 334 1037 368
rect 1071 334 1105 368
rect 1139 334 1173 368
rect 1207 334 1241 368
rect 1275 334 1309 368
rect 1343 334 1377 368
rect 1411 334 1445 368
rect 1479 334 1513 368
rect 1547 334 1581 368
rect 1615 334 1649 368
rect 1683 334 1717 368
rect 1751 334 1785 368
rect 1819 334 1853 368
rect 1887 334 1921 368
rect 1955 334 1989 368
rect 2023 334 2130 368
rect -2130 255 -2096 334
rect 2096 255 2130 334
rect -2130 187 -2096 221
rect -2000 188 -1955 222
rect -1921 188 -1887 222
rect -1853 188 -1819 222
rect -1785 188 -1751 222
rect -1717 188 -1683 222
rect -1649 188 -1615 222
rect -1581 188 -1547 222
rect -1513 188 -1479 222
rect -1445 188 -1411 222
rect -1377 188 -1343 222
rect -1309 188 -1275 222
rect -1241 188 -1207 222
rect -1173 188 -1139 222
rect -1105 188 -1071 222
rect -1037 188 -1003 222
rect -969 188 -935 222
rect -901 188 -867 222
rect -833 188 -799 222
rect -765 188 -731 222
rect -697 188 -663 222
rect -629 188 -595 222
rect -561 188 -527 222
rect -493 188 -459 222
rect -425 188 -391 222
rect -357 188 -323 222
rect -289 188 -255 222
rect -221 188 -187 222
rect -153 188 -119 222
rect -85 188 -51 222
rect -17 188 17 222
rect 51 188 85 222
rect 119 188 153 222
rect 187 188 221 222
rect 255 188 289 222
rect 323 188 357 222
rect 391 188 425 222
rect 459 188 493 222
rect 527 188 561 222
rect 595 188 629 222
rect 663 188 697 222
rect 731 188 765 222
rect 799 188 833 222
rect 867 188 901 222
rect 935 188 969 222
rect 1003 188 1037 222
rect 1071 188 1105 222
rect 1139 188 1173 222
rect 1207 188 1241 222
rect 1275 188 1309 222
rect 1343 188 1377 222
rect 1411 188 1445 222
rect 1479 188 1513 222
rect 1547 188 1581 222
rect 1615 188 1649 222
rect 1683 188 1717 222
rect 1751 188 1785 222
rect 1819 188 1853 222
rect 1887 188 1921 222
rect 1955 188 2000 222
rect -2130 119 -2096 153
rect -2130 51 -2096 85
rect -2130 -17 -2096 17
rect -2130 -85 -2096 -51
rect -2130 -153 -2096 -119
rect -2130 -221 -2096 -187
rect 2096 187 2130 221
rect 2096 119 2130 153
rect 2096 51 2130 85
rect 2096 -17 2130 17
rect 2096 -85 2130 -51
rect 2096 -153 2130 -119
rect -2000 -222 -1955 -188
rect -1921 -222 -1887 -188
rect -1853 -222 -1819 -188
rect -1785 -222 -1751 -188
rect -1717 -222 -1683 -188
rect -1649 -222 -1615 -188
rect -1581 -222 -1547 -188
rect -1513 -222 -1479 -188
rect -1445 -222 -1411 -188
rect -1377 -222 -1343 -188
rect -1309 -222 -1275 -188
rect -1241 -222 -1207 -188
rect -1173 -222 -1139 -188
rect -1105 -222 -1071 -188
rect -1037 -222 -1003 -188
rect -969 -222 -935 -188
rect -901 -222 -867 -188
rect -833 -222 -799 -188
rect -765 -222 -731 -188
rect -697 -222 -663 -188
rect -629 -222 -595 -188
rect -561 -222 -527 -188
rect -493 -222 -459 -188
rect -425 -222 -391 -188
rect -357 -222 -323 -188
rect -289 -222 -255 -188
rect -221 -222 -187 -188
rect -153 -222 -119 -188
rect -85 -222 -51 -188
rect -17 -222 17 -188
rect 51 -222 85 -188
rect 119 -222 153 -188
rect 187 -222 221 -188
rect 255 -222 289 -188
rect 323 -222 357 -188
rect 391 -222 425 -188
rect 459 -222 493 -188
rect 527 -222 561 -188
rect 595 -222 629 -188
rect 663 -222 697 -188
rect 731 -222 765 -188
rect 799 -222 833 -188
rect 867 -222 901 -188
rect 935 -222 969 -188
rect 1003 -222 1037 -188
rect 1071 -222 1105 -188
rect 1139 -222 1173 -188
rect 1207 -222 1241 -188
rect 1275 -222 1309 -188
rect 1343 -222 1377 -188
rect 1411 -222 1445 -188
rect 1479 -222 1513 -188
rect 1547 -222 1581 -188
rect 1615 -222 1649 -188
rect 1683 -222 1717 -188
rect 1751 -222 1785 -188
rect 1819 -222 1853 -188
rect 1887 -222 1921 -188
rect 1955 -222 2000 -188
rect 2096 -221 2130 -187
rect -2130 -334 -2096 -255
rect 2096 -334 2130 -255
rect -2130 -368 -2023 -334
rect -1989 -368 -1955 -334
rect -1921 -368 -1887 -334
rect -1853 -368 -1819 -334
rect -1785 -368 -1751 -334
rect -1717 -368 -1683 -334
rect -1649 -368 -1615 -334
rect -1581 -368 -1547 -334
rect -1513 -368 -1479 -334
rect -1445 -368 -1411 -334
rect -1377 -368 -1343 -334
rect -1309 -368 -1275 -334
rect -1241 -368 -1207 -334
rect -1173 -368 -1139 -334
rect -1105 -368 -1071 -334
rect -1037 -368 -1003 -334
rect -969 -368 -935 -334
rect -901 -368 -867 -334
rect -833 -368 -799 -334
rect -765 -368 -731 -334
rect -697 -368 -663 -334
rect -629 -368 -595 -334
rect -561 -368 -527 -334
rect -493 -368 -459 -334
rect -425 -368 -391 -334
rect -357 -368 -323 -334
rect -289 -368 -255 -334
rect -221 -368 -187 -334
rect -153 -368 -119 -334
rect -85 -368 -51 -334
rect -17 -368 17 -334
rect 51 -368 85 -334
rect 119 -368 153 -334
rect 187 -368 221 -334
rect 255 -368 289 -334
rect 323 -368 357 -334
rect 391 -368 425 -334
rect 459 -368 493 -334
rect 527 -368 561 -334
rect 595 -368 629 -334
rect 663 -368 697 -334
rect 731 -368 765 -334
rect 799 -368 833 -334
rect 867 -368 901 -334
rect 935 -368 969 -334
rect 1003 -368 1037 -334
rect 1071 -368 1105 -334
rect 1139 -368 1173 -334
rect 1207 -368 1241 -334
rect 1275 -368 1309 -334
rect 1343 -368 1377 -334
rect 1411 -368 1445 -334
rect 1479 -368 1513 -334
rect 1547 -368 1581 -334
rect 1615 -368 1649 -334
rect 1683 -368 1717 -334
rect 1751 -368 1785 -334
rect 1819 -368 1853 -334
rect 1887 -368 1921 -334
rect 1955 -368 1989 -334
rect 2023 -368 2130 -334
<< properties >>
string FIXED_BBOX -2113 -351 2113 351
<< end >>
