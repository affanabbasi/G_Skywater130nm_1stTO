magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -2421 1460 2421 1494
rect -2421 -1460 -2387 1460
rect 2387 -1460 2421 1460
rect -2421 -1494 2421 -1460
<< nmoslvt >>
rect -2261 -1320 -1861 1320
rect -1803 -1320 -1403 1320
rect -1345 -1320 -945 1320
rect -887 -1320 -487 1320
rect -429 -1320 -29 1320
rect 29 -1320 429 1320
rect 487 -1320 887 1320
rect 945 -1320 1345 1320
rect 1403 -1320 1803 1320
rect 1861 -1320 2261 1320
<< ndiff >>
rect -2319 1275 -2261 1320
rect -2319 1241 -2307 1275
rect -2273 1241 -2261 1275
rect -2319 1207 -2261 1241
rect -2319 1173 -2307 1207
rect -2273 1173 -2261 1207
rect -2319 1139 -2261 1173
rect -2319 1105 -2307 1139
rect -2273 1105 -2261 1139
rect -2319 1071 -2261 1105
rect -2319 1037 -2307 1071
rect -2273 1037 -2261 1071
rect -2319 1003 -2261 1037
rect -2319 969 -2307 1003
rect -2273 969 -2261 1003
rect -2319 935 -2261 969
rect -2319 901 -2307 935
rect -2273 901 -2261 935
rect -2319 867 -2261 901
rect -2319 833 -2307 867
rect -2273 833 -2261 867
rect -2319 799 -2261 833
rect -2319 765 -2307 799
rect -2273 765 -2261 799
rect -2319 731 -2261 765
rect -2319 697 -2307 731
rect -2273 697 -2261 731
rect -2319 663 -2261 697
rect -2319 629 -2307 663
rect -2273 629 -2261 663
rect -2319 595 -2261 629
rect -2319 561 -2307 595
rect -2273 561 -2261 595
rect -2319 527 -2261 561
rect -2319 493 -2307 527
rect -2273 493 -2261 527
rect -2319 459 -2261 493
rect -2319 425 -2307 459
rect -2273 425 -2261 459
rect -2319 391 -2261 425
rect -2319 357 -2307 391
rect -2273 357 -2261 391
rect -2319 323 -2261 357
rect -2319 289 -2307 323
rect -2273 289 -2261 323
rect -2319 255 -2261 289
rect -2319 221 -2307 255
rect -2273 221 -2261 255
rect -2319 187 -2261 221
rect -2319 153 -2307 187
rect -2273 153 -2261 187
rect -2319 119 -2261 153
rect -2319 85 -2307 119
rect -2273 85 -2261 119
rect -2319 51 -2261 85
rect -2319 17 -2307 51
rect -2273 17 -2261 51
rect -2319 -17 -2261 17
rect -2319 -51 -2307 -17
rect -2273 -51 -2261 -17
rect -2319 -85 -2261 -51
rect -2319 -119 -2307 -85
rect -2273 -119 -2261 -85
rect -2319 -153 -2261 -119
rect -2319 -187 -2307 -153
rect -2273 -187 -2261 -153
rect -2319 -221 -2261 -187
rect -2319 -255 -2307 -221
rect -2273 -255 -2261 -221
rect -2319 -289 -2261 -255
rect -2319 -323 -2307 -289
rect -2273 -323 -2261 -289
rect -2319 -357 -2261 -323
rect -2319 -391 -2307 -357
rect -2273 -391 -2261 -357
rect -2319 -425 -2261 -391
rect -2319 -459 -2307 -425
rect -2273 -459 -2261 -425
rect -2319 -493 -2261 -459
rect -2319 -527 -2307 -493
rect -2273 -527 -2261 -493
rect -2319 -561 -2261 -527
rect -2319 -595 -2307 -561
rect -2273 -595 -2261 -561
rect -2319 -629 -2261 -595
rect -2319 -663 -2307 -629
rect -2273 -663 -2261 -629
rect -2319 -697 -2261 -663
rect -2319 -731 -2307 -697
rect -2273 -731 -2261 -697
rect -2319 -765 -2261 -731
rect -2319 -799 -2307 -765
rect -2273 -799 -2261 -765
rect -2319 -833 -2261 -799
rect -2319 -867 -2307 -833
rect -2273 -867 -2261 -833
rect -2319 -901 -2261 -867
rect -2319 -935 -2307 -901
rect -2273 -935 -2261 -901
rect -2319 -969 -2261 -935
rect -2319 -1003 -2307 -969
rect -2273 -1003 -2261 -969
rect -2319 -1037 -2261 -1003
rect -2319 -1071 -2307 -1037
rect -2273 -1071 -2261 -1037
rect -2319 -1105 -2261 -1071
rect -2319 -1139 -2307 -1105
rect -2273 -1139 -2261 -1105
rect -2319 -1173 -2261 -1139
rect -2319 -1207 -2307 -1173
rect -2273 -1207 -2261 -1173
rect -2319 -1241 -2261 -1207
rect -2319 -1275 -2307 -1241
rect -2273 -1275 -2261 -1241
rect -2319 -1320 -2261 -1275
rect -1861 1275 -1803 1320
rect -1861 1241 -1849 1275
rect -1815 1241 -1803 1275
rect -1861 1207 -1803 1241
rect -1861 1173 -1849 1207
rect -1815 1173 -1803 1207
rect -1861 1139 -1803 1173
rect -1861 1105 -1849 1139
rect -1815 1105 -1803 1139
rect -1861 1071 -1803 1105
rect -1861 1037 -1849 1071
rect -1815 1037 -1803 1071
rect -1861 1003 -1803 1037
rect -1861 969 -1849 1003
rect -1815 969 -1803 1003
rect -1861 935 -1803 969
rect -1861 901 -1849 935
rect -1815 901 -1803 935
rect -1861 867 -1803 901
rect -1861 833 -1849 867
rect -1815 833 -1803 867
rect -1861 799 -1803 833
rect -1861 765 -1849 799
rect -1815 765 -1803 799
rect -1861 731 -1803 765
rect -1861 697 -1849 731
rect -1815 697 -1803 731
rect -1861 663 -1803 697
rect -1861 629 -1849 663
rect -1815 629 -1803 663
rect -1861 595 -1803 629
rect -1861 561 -1849 595
rect -1815 561 -1803 595
rect -1861 527 -1803 561
rect -1861 493 -1849 527
rect -1815 493 -1803 527
rect -1861 459 -1803 493
rect -1861 425 -1849 459
rect -1815 425 -1803 459
rect -1861 391 -1803 425
rect -1861 357 -1849 391
rect -1815 357 -1803 391
rect -1861 323 -1803 357
rect -1861 289 -1849 323
rect -1815 289 -1803 323
rect -1861 255 -1803 289
rect -1861 221 -1849 255
rect -1815 221 -1803 255
rect -1861 187 -1803 221
rect -1861 153 -1849 187
rect -1815 153 -1803 187
rect -1861 119 -1803 153
rect -1861 85 -1849 119
rect -1815 85 -1803 119
rect -1861 51 -1803 85
rect -1861 17 -1849 51
rect -1815 17 -1803 51
rect -1861 -17 -1803 17
rect -1861 -51 -1849 -17
rect -1815 -51 -1803 -17
rect -1861 -85 -1803 -51
rect -1861 -119 -1849 -85
rect -1815 -119 -1803 -85
rect -1861 -153 -1803 -119
rect -1861 -187 -1849 -153
rect -1815 -187 -1803 -153
rect -1861 -221 -1803 -187
rect -1861 -255 -1849 -221
rect -1815 -255 -1803 -221
rect -1861 -289 -1803 -255
rect -1861 -323 -1849 -289
rect -1815 -323 -1803 -289
rect -1861 -357 -1803 -323
rect -1861 -391 -1849 -357
rect -1815 -391 -1803 -357
rect -1861 -425 -1803 -391
rect -1861 -459 -1849 -425
rect -1815 -459 -1803 -425
rect -1861 -493 -1803 -459
rect -1861 -527 -1849 -493
rect -1815 -527 -1803 -493
rect -1861 -561 -1803 -527
rect -1861 -595 -1849 -561
rect -1815 -595 -1803 -561
rect -1861 -629 -1803 -595
rect -1861 -663 -1849 -629
rect -1815 -663 -1803 -629
rect -1861 -697 -1803 -663
rect -1861 -731 -1849 -697
rect -1815 -731 -1803 -697
rect -1861 -765 -1803 -731
rect -1861 -799 -1849 -765
rect -1815 -799 -1803 -765
rect -1861 -833 -1803 -799
rect -1861 -867 -1849 -833
rect -1815 -867 -1803 -833
rect -1861 -901 -1803 -867
rect -1861 -935 -1849 -901
rect -1815 -935 -1803 -901
rect -1861 -969 -1803 -935
rect -1861 -1003 -1849 -969
rect -1815 -1003 -1803 -969
rect -1861 -1037 -1803 -1003
rect -1861 -1071 -1849 -1037
rect -1815 -1071 -1803 -1037
rect -1861 -1105 -1803 -1071
rect -1861 -1139 -1849 -1105
rect -1815 -1139 -1803 -1105
rect -1861 -1173 -1803 -1139
rect -1861 -1207 -1849 -1173
rect -1815 -1207 -1803 -1173
rect -1861 -1241 -1803 -1207
rect -1861 -1275 -1849 -1241
rect -1815 -1275 -1803 -1241
rect -1861 -1320 -1803 -1275
rect -1403 1275 -1345 1320
rect -1403 1241 -1391 1275
rect -1357 1241 -1345 1275
rect -1403 1207 -1345 1241
rect -1403 1173 -1391 1207
rect -1357 1173 -1345 1207
rect -1403 1139 -1345 1173
rect -1403 1105 -1391 1139
rect -1357 1105 -1345 1139
rect -1403 1071 -1345 1105
rect -1403 1037 -1391 1071
rect -1357 1037 -1345 1071
rect -1403 1003 -1345 1037
rect -1403 969 -1391 1003
rect -1357 969 -1345 1003
rect -1403 935 -1345 969
rect -1403 901 -1391 935
rect -1357 901 -1345 935
rect -1403 867 -1345 901
rect -1403 833 -1391 867
rect -1357 833 -1345 867
rect -1403 799 -1345 833
rect -1403 765 -1391 799
rect -1357 765 -1345 799
rect -1403 731 -1345 765
rect -1403 697 -1391 731
rect -1357 697 -1345 731
rect -1403 663 -1345 697
rect -1403 629 -1391 663
rect -1357 629 -1345 663
rect -1403 595 -1345 629
rect -1403 561 -1391 595
rect -1357 561 -1345 595
rect -1403 527 -1345 561
rect -1403 493 -1391 527
rect -1357 493 -1345 527
rect -1403 459 -1345 493
rect -1403 425 -1391 459
rect -1357 425 -1345 459
rect -1403 391 -1345 425
rect -1403 357 -1391 391
rect -1357 357 -1345 391
rect -1403 323 -1345 357
rect -1403 289 -1391 323
rect -1357 289 -1345 323
rect -1403 255 -1345 289
rect -1403 221 -1391 255
rect -1357 221 -1345 255
rect -1403 187 -1345 221
rect -1403 153 -1391 187
rect -1357 153 -1345 187
rect -1403 119 -1345 153
rect -1403 85 -1391 119
rect -1357 85 -1345 119
rect -1403 51 -1345 85
rect -1403 17 -1391 51
rect -1357 17 -1345 51
rect -1403 -17 -1345 17
rect -1403 -51 -1391 -17
rect -1357 -51 -1345 -17
rect -1403 -85 -1345 -51
rect -1403 -119 -1391 -85
rect -1357 -119 -1345 -85
rect -1403 -153 -1345 -119
rect -1403 -187 -1391 -153
rect -1357 -187 -1345 -153
rect -1403 -221 -1345 -187
rect -1403 -255 -1391 -221
rect -1357 -255 -1345 -221
rect -1403 -289 -1345 -255
rect -1403 -323 -1391 -289
rect -1357 -323 -1345 -289
rect -1403 -357 -1345 -323
rect -1403 -391 -1391 -357
rect -1357 -391 -1345 -357
rect -1403 -425 -1345 -391
rect -1403 -459 -1391 -425
rect -1357 -459 -1345 -425
rect -1403 -493 -1345 -459
rect -1403 -527 -1391 -493
rect -1357 -527 -1345 -493
rect -1403 -561 -1345 -527
rect -1403 -595 -1391 -561
rect -1357 -595 -1345 -561
rect -1403 -629 -1345 -595
rect -1403 -663 -1391 -629
rect -1357 -663 -1345 -629
rect -1403 -697 -1345 -663
rect -1403 -731 -1391 -697
rect -1357 -731 -1345 -697
rect -1403 -765 -1345 -731
rect -1403 -799 -1391 -765
rect -1357 -799 -1345 -765
rect -1403 -833 -1345 -799
rect -1403 -867 -1391 -833
rect -1357 -867 -1345 -833
rect -1403 -901 -1345 -867
rect -1403 -935 -1391 -901
rect -1357 -935 -1345 -901
rect -1403 -969 -1345 -935
rect -1403 -1003 -1391 -969
rect -1357 -1003 -1345 -969
rect -1403 -1037 -1345 -1003
rect -1403 -1071 -1391 -1037
rect -1357 -1071 -1345 -1037
rect -1403 -1105 -1345 -1071
rect -1403 -1139 -1391 -1105
rect -1357 -1139 -1345 -1105
rect -1403 -1173 -1345 -1139
rect -1403 -1207 -1391 -1173
rect -1357 -1207 -1345 -1173
rect -1403 -1241 -1345 -1207
rect -1403 -1275 -1391 -1241
rect -1357 -1275 -1345 -1241
rect -1403 -1320 -1345 -1275
rect -945 1275 -887 1320
rect -945 1241 -933 1275
rect -899 1241 -887 1275
rect -945 1207 -887 1241
rect -945 1173 -933 1207
rect -899 1173 -887 1207
rect -945 1139 -887 1173
rect -945 1105 -933 1139
rect -899 1105 -887 1139
rect -945 1071 -887 1105
rect -945 1037 -933 1071
rect -899 1037 -887 1071
rect -945 1003 -887 1037
rect -945 969 -933 1003
rect -899 969 -887 1003
rect -945 935 -887 969
rect -945 901 -933 935
rect -899 901 -887 935
rect -945 867 -887 901
rect -945 833 -933 867
rect -899 833 -887 867
rect -945 799 -887 833
rect -945 765 -933 799
rect -899 765 -887 799
rect -945 731 -887 765
rect -945 697 -933 731
rect -899 697 -887 731
rect -945 663 -887 697
rect -945 629 -933 663
rect -899 629 -887 663
rect -945 595 -887 629
rect -945 561 -933 595
rect -899 561 -887 595
rect -945 527 -887 561
rect -945 493 -933 527
rect -899 493 -887 527
rect -945 459 -887 493
rect -945 425 -933 459
rect -899 425 -887 459
rect -945 391 -887 425
rect -945 357 -933 391
rect -899 357 -887 391
rect -945 323 -887 357
rect -945 289 -933 323
rect -899 289 -887 323
rect -945 255 -887 289
rect -945 221 -933 255
rect -899 221 -887 255
rect -945 187 -887 221
rect -945 153 -933 187
rect -899 153 -887 187
rect -945 119 -887 153
rect -945 85 -933 119
rect -899 85 -887 119
rect -945 51 -887 85
rect -945 17 -933 51
rect -899 17 -887 51
rect -945 -17 -887 17
rect -945 -51 -933 -17
rect -899 -51 -887 -17
rect -945 -85 -887 -51
rect -945 -119 -933 -85
rect -899 -119 -887 -85
rect -945 -153 -887 -119
rect -945 -187 -933 -153
rect -899 -187 -887 -153
rect -945 -221 -887 -187
rect -945 -255 -933 -221
rect -899 -255 -887 -221
rect -945 -289 -887 -255
rect -945 -323 -933 -289
rect -899 -323 -887 -289
rect -945 -357 -887 -323
rect -945 -391 -933 -357
rect -899 -391 -887 -357
rect -945 -425 -887 -391
rect -945 -459 -933 -425
rect -899 -459 -887 -425
rect -945 -493 -887 -459
rect -945 -527 -933 -493
rect -899 -527 -887 -493
rect -945 -561 -887 -527
rect -945 -595 -933 -561
rect -899 -595 -887 -561
rect -945 -629 -887 -595
rect -945 -663 -933 -629
rect -899 -663 -887 -629
rect -945 -697 -887 -663
rect -945 -731 -933 -697
rect -899 -731 -887 -697
rect -945 -765 -887 -731
rect -945 -799 -933 -765
rect -899 -799 -887 -765
rect -945 -833 -887 -799
rect -945 -867 -933 -833
rect -899 -867 -887 -833
rect -945 -901 -887 -867
rect -945 -935 -933 -901
rect -899 -935 -887 -901
rect -945 -969 -887 -935
rect -945 -1003 -933 -969
rect -899 -1003 -887 -969
rect -945 -1037 -887 -1003
rect -945 -1071 -933 -1037
rect -899 -1071 -887 -1037
rect -945 -1105 -887 -1071
rect -945 -1139 -933 -1105
rect -899 -1139 -887 -1105
rect -945 -1173 -887 -1139
rect -945 -1207 -933 -1173
rect -899 -1207 -887 -1173
rect -945 -1241 -887 -1207
rect -945 -1275 -933 -1241
rect -899 -1275 -887 -1241
rect -945 -1320 -887 -1275
rect -487 1275 -429 1320
rect -487 1241 -475 1275
rect -441 1241 -429 1275
rect -487 1207 -429 1241
rect -487 1173 -475 1207
rect -441 1173 -429 1207
rect -487 1139 -429 1173
rect -487 1105 -475 1139
rect -441 1105 -429 1139
rect -487 1071 -429 1105
rect -487 1037 -475 1071
rect -441 1037 -429 1071
rect -487 1003 -429 1037
rect -487 969 -475 1003
rect -441 969 -429 1003
rect -487 935 -429 969
rect -487 901 -475 935
rect -441 901 -429 935
rect -487 867 -429 901
rect -487 833 -475 867
rect -441 833 -429 867
rect -487 799 -429 833
rect -487 765 -475 799
rect -441 765 -429 799
rect -487 731 -429 765
rect -487 697 -475 731
rect -441 697 -429 731
rect -487 663 -429 697
rect -487 629 -475 663
rect -441 629 -429 663
rect -487 595 -429 629
rect -487 561 -475 595
rect -441 561 -429 595
rect -487 527 -429 561
rect -487 493 -475 527
rect -441 493 -429 527
rect -487 459 -429 493
rect -487 425 -475 459
rect -441 425 -429 459
rect -487 391 -429 425
rect -487 357 -475 391
rect -441 357 -429 391
rect -487 323 -429 357
rect -487 289 -475 323
rect -441 289 -429 323
rect -487 255 -429 289
rect -487 221 -475 255
rect -441 221 -429 255
rect -487 187 -429 221
rect -487 153 -475 187
rect -441 153 -429 187
rect -487 119 -429 153
rect -487 85 -475 119
rect -441 85 -429 119
rect -487 51 -429 85
rect -487 17 -475 51
rect -441 17 -429 51
rect -487 -17 -429 17
rect -487 -51 -475 -17
rect -441 -51 -429 -17
rect -487 -85 -429 -51
rect -487 -119 -475 -85
rect -441 -119 -429 -85
rect -487 -153 -429 -119
rect -487 -187 -475 -153
rect -441 -187 -429 -153
rect -487 -221 -429 -187
rect -487 -255 -475 -221
rect -441 -255 -429 -221
rect -487 -289 -429 -255
rect -487 -323 -475 -289
rect -441 -323 -429 -289
rect -487 -357 -429 -323
rect -487 -391 -475 -357
rect -441 -391 -429 -357
rect -487 -425 -429 -391
rect -487 -459 -475 -425
rect -441 -459 -429 -425
rect -487 -493 -429 -459
rect -487 -527 -475 -493
rect -441 -527 -429 -493
rect -487 -561 -429 -527
rect -487 -595 -475 -561
rect -441 -595 -429 -561
rect -487 -629 -429 -595
rect -487 -663 -475 -629
rect -441 -663 -429 -629
rect -487 -697 -429 -663
rect -487 -731 -475 -697
rect -441 -731 -429 -697
rect -487 -765 -429 -731
rect -487 -799 -475 -765
rect -441 -799 -429 -765
rect -487 -833 -429 -799
rect -487 -867 -475 -833
rect -441 -867 -429 -833
rect -487 -901 -429 -867
rect -487 -935 -475 -901
rect -441 -935 -429 -901
rect -487 -969 -429 -935
rect -487 -1003 -475 -969
rect -441 -1003 -429 -969
rect -487 -1037 -429 -1003
rect -487 -1071 -475 -1037
rect -441 -1071 -429 -1037
rect -487 -1105 -429 -1071
rect -487 -1139 -475 -1105
rect -441 -1139 -429 -1105
rect -487 -1173 -429 -1139
rect -487 -1207 -475 -1173
rect -441 -1207 -429 -1173
rect -487 -1241 -429 -1207
rect -487 -1275 -475 -1241
rect -441 -1275 -429 -1241
rect -487 -1320 -429 -1275
rect -29 1275 29 1320
rect -29 1241 -17 1275
rect 17 1241 29 1275
rect -29 1207 29 1241
rect -29 1173 -17 1207
rect 17 1173 29 1207
rect -29 1139 29 1173
rect -29 1105 -17 1139
rect 17 1105 29 1139
rect -29 1071 29 1105
rect -29 1037 -17 1071
rect 17 1037 29 1071
rect -29 1003 29 1037
rect -29 969 -17 1003
rect 17 969 29 1003
rect -29 935 29 969
rect -29 901 -17 935
rect 17 901 29 935
rect -29 867 29 901
rect -29 833 -17 867
rect 17 833 29 867
rect -29 799 29 833
rect -29 765 -17 799
rect 17 765 29 799
rect -29 731 29 765
rect -29 697 -17 731
rect 17 697 29 731
rect -29 663 29 697
rect -29 629 -17 663
rect 17 629 29 663
rect -29 595 29 629
rect -29 561 -17 595
rect 17 561 29 595
rect -29 527 29 561
rect -29 493 -17 527
rect 17 493 29 527
rect -29 459 29 493
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -493 29 -459
rect -29 -527 -17 -493
rect 17 -527 29 -493
rect -29 -561 29 -527
rect -29 -595 -17 -561
rect 17 -595 29 -561
rect -29 -629 29 -595
rect -29 -663 -17 -629
rect 17 -663 29 -629
rect -29 -697 29 -663
rect -29 -731 -17 -697
rect 17 -731 29 -697
rect -29 -765 29 -731
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -833 29 -799
rect -29 -867 -17 -833
rect 17 -867 29 -833
rect -29 -901 29 -867
rect -29 -935 -17 -901
rect 17 -935 29 -901
rect -29 -969 29 -935
rect -29 -1003 -17 -969
rect 17 -1003 29 -969
rect -29 -1037 29 -1003
rect -29 -1071 -17 -1037
rect 17 -1071 29 -1037
rect -29 -1105 29 -1071
rect -29 -1139 -17 -1105
rect 17 -1139 29 -1105
rect -29 -1173 29 -1139
rect -29 -1207 -17 -1173
rect 17 -1207 29 -1173
rect -29 -1241 29 -1207
rect -29 -1275 -17 -1241
rect 17 -1275 29 -1241
rect -29 -1320 29 -1275
rect 429 1275 487 1320
rect 429 1241 441 1275
rect 475 1241 487 1275
rect 429 1207 487 1241
rect 429 1173 441 1207
rect 475 1173 487 1207
rect 429 1139 487 1173
rect 429 1105 441 1139
rect 475 1105 487 1139
rect 429 1071 487 1105
rect 429 1037 441 1071
rect 475 1037 487 1071
rect 429 1003 487 1037
rect 429 969 441 1003
rect 475 969 487 1003
rect 429 935 487 969
rect 429 901 441 935
rect 475 901 487 935
rect 429 867 487 901
rect 429 833 441 867
rect 475 833 487 867
rect 429 799 487 833
rect 429 765 441 799
rect 475 765 487 799
rect 429 731 487 765
rect 429 697 441 731
rect 475 697 487 731
rect 429 663 487 697
rect 429 629 441 663
rect 475 629 487 663
rect 429 595 487 629
rect 429 561 441 595
rect 475 561 487 595
rect 429 527 487 561
rect 429 493 441 527
rect 475 493 487 527
rect 429 459 487 493
rect 429 425 441 459
rect 475 425 487 459
rect 429 391 487 425
rect 429 357 441 391
rect 475 357 487 391
rect 429 323 487 357
rect 429 289 441 323
rect 475 289 487 323
rect 429 255 487 289
rect 429 221 441 255
rect 475 221 487 255
rect 429 187 487 221
rect 429 153 441 187
rect 475 153 487 187
rect 429 119 487 153
rect 429 85 441 119
rect 475 85 487 119
rect 429 51 487 85
rect 429 17 441 51
rect 475 17 487 51
rect 429 -17 487 17
rect 429 -51 441 -17
rect 475 -51 487 -17
rect 429 -85 487 -51
rect 429 -119 441 -85
rect 475 -119 487 -85
rect 429 -153 487 -119
rect 429 -187 441 -153
rect 475 -187 487 -153
rect 429 -221 487 -187
rect 429 -255 441 -221
rect 475 -255 487 -221
rect 429 -289 487 -255
rect 429 -323 441 -289
rect 475 -323 487 -289
rect 429 -357 487 -323
rect 429 -391 441 -357
rect 475 -391 487 -357
rect 429 -425 487 -391
rect 429 -459 441 -425
rect 475 -459 487 -425
rect 429 -493 487 -459
rect 429 -527 441 -493
rect 475 -527 487 -493
rect 429 -561 487 -527
rect 429 -595 441 -561
rect 475 -595 487 -561
rect 429 -629 487 -595
rect 429 -663 441 -629
rect 475 -663 487 -629
rect 429 -697 487 -663
rect 429 -731 441 -697
rect 475 -731 487 -697
rect 429 -765 487 -731
rect 429 -799 441 -765
rect 475 -799 487 -765
rect 429 -833 487 -799
rect 429 -867 441 -833
rect 475 -867 487 -833
rect 429 -901 487 -867
rect 429 -935 441 -901
rect 475 -935 487 -901
rect 429 -969 487 -935
rect 429 -1003 441 -969
rect 475 -1003 487 -969
rect 429 -1037 487 -1003
rect 429 -1071 441 -1037
rect 475 -1071 487 -1037
rect 429 -1105 487 -1071
rect 429 -1139 441 -1105
rect 475 -1139 487 -1105
rect 429 -1173 487 -1139
rect 429 -1207 441 -1173
rect 475 -1207 487 -1173
rect 429 -1241 487 -1207
rect 429 -1275 441 -1241
rect 475 -1275 487 -1241
rect 429 -1320 487 -1275
rect 887 1275 945 1320
rect 887 1241 899 1275
rect 933 1241 945 1275
rect 887 1207 945 1241
rect 887 1173 899 1207
rect 933 1173 945 1207
rect 887 1139 945 1173
rect 887 1105 899 1139
rect 933 1105 945 1139
rect 887 1071 945 1105
rect 887 1037 899 1071
rect 933 1037 945 1071
rect 887 1003 945 1037
rect 887 969 899 1003
rect 933 969 945 1003
rect 887 935 945 969
rect 887 901 899 935
rect 933 901 945 935
rect 887 867 945 901
rect 887 833 899 867
rect 933 833 945 867
rect 887 799 945 833
rect 887 765 899 799
rect 933 765 945 799
rect 887 731 945 765
rect 887 697 899 731
rect 933 697 945 731
rect 887 663 945 697
rect 887 629 899 663
rect 933 629 945 663
rect 887 595 945 629
rect 887 561 899 595
rect 933 561 945 595
rect 887 527 945 561
rect 887 493 899 527
rect 933 493 945 527
rect 887 459 945 493
rect 887 425 899 459
rect 933 425 945 459
rect 887 391 945 425
rect 887 357 899 391
rect 933 357 945 391
rect 887 323 945 357
rect 887 289 899 323
rect 933 289 945 323
rect 887 255 945 289
rect 887 221 899 255
rect 933 221 945 255
rect 887 187 945 221
rect 887 153 899 187
rect 933 153 945 187
rect 887 119 945 153
rect 887 85 899 119
rect 933 85 945 119
rect 887 51 945 85
rect 887 17 899 51
rect 933 17 945 51
rect 887 -17 945 17
rect 887 -51 899 -17
rect 933 -51 945 -17
rect 887 -85 945 -51
rect 887 -119 899 -85
rect 933 -119 945 -85
rect 887 -153 945 -119
rect 887 -187 899 -153
rect 933 -187 945 -153
rect 887 -221 945 -187
rect 887 -255 899 -221
rect 933 -255 945 -221
rect 887 -289 945 -255
rect 887 -323 899 -289
rect 933 -323 945 -289
rect 887 -357 945 -323
rect 887 -391 899 -357
rect 933 -391 945 -357
rect 887 -425 945 -391
rect 887 -459 899 -425
rect 933 -459 945 -425
rect 887 -493 945 -459
rect 887 -527 899 -493
rect 933 -527 945 -493
rect 887 -561 945 -527
rect 887 -595 899 -561
rect 933 -595 945 -561
rect 887 -629 945 -595
rect 887 -663 899 -629
rect 933 -663 945 -629
rect 887 -697 945 -663
rect 887 -731 899 -697
rect 933 -731 945 -697
rect 887 -765 945 -731
rect 887 -799 899 -765
rect 933 -799 945 -765
rect 887 -833 945 -799
rect 887 -867 899 -833
rect 933 -867 945 -833
rect 887 -901 945 -867
rect 887 -935 899 -901
rect 933 -935 945 -901
rect 887 -969 945 -935
rect 887 -1003 899 -969
rect 933 -1003 945 -969
rect 887 -1037 945 -1003
rect 887 -1071 899 -1037
rect 933 -1071 945 -1037
rect 887 -1105 945 -1071
rect 887 -1139 899 -1105
rect 933 -1139 945 -1105
rect 887 -1173 945 -1139
rect 887 -1207 899 -1173
rect 933 -1207 945 -1173
rect 887 -1241 945 -1207
rect 887 -1275 899 -1241
rect 933 -1275 945 -1241
rect 887 -1320 945 -1275
rect 1345 1275 1403 1320
rect 1345 1241 1357 1275
rect 1391 1241 1403 1275
rect 1345 1207 1403 1241
rect 1345 1173 1357 1207
rect 1391 1173 1403 1207
rect 1345 1139 1403 1173
rect 1345 1105 1357 1139
rect 1391 1105 1403 1139
rect 1345 1071 1403 1105
rect 1345 1037 1357 1071
rect 1391 1037 1403 1071
rect 1345 1003 1403 1037
rect 1345 969 1357 1003
rect 1391 969 1403 1003
rect 1345 935 1403 969
rect 1345 901 1357 935
rect 1391 901 1403 935
rect 1345 867 1403 901
rect 1345 833 1357 867
rect 1391 833 1403 867
rect 1345 799 1403 833
rect 1345 765 1357 799
rect 1391 765 1403 799
rect 1345 731 1403 765
rect 1345 697 1357 731
rect 1391 697 1403 731
rect 1345 663 1403 697
rect 1345 629 1357 663
rect 1391 629 1403 663
rect 1345 595 1403 629
rect 1345 561 1357 595
rect 1391 561 1403 595
rect 1345 527 1403 561
rect 1345 493 1357 527
rect 1391 493 1403 527
rect 1345 459 1403 493
rect 1345 425 1357 459
rect 1391 425 1403 459
rect 1345 391 1403 425
rect 1345 357 1357 391
rect 1391 357 1403 391
rect 1345 323 1403 357
rect 1345 289 1357 323
rect 1391 289 1403 323
rect 1345 255 1403 289
rect 1345 221 1357 255
rect 1391 221 1403 255
rect 1345 187 1403 221
rect 1345 153 1357 187
rect 1391 153 1403 187
rect 1345 119 1403 153
rect 1345 85 1357 119
rect 1391 85 1403 119
rect 1345 51 1403 85
rect 1345 17 1357 51
rect 1391 17 1403 51
rect 1345 -17 1403 17
rect 1345 -51 1357 -17
rect 1391 -51 1403 -17
rect 1345 -85 1403 -51
rect 1345 -119 1357 -85
rect 1391 -119 1403 -85
rect 1345 -153 1403 -119
rect 1345 -187 1357 -153
rect 1391 -187 1403 -153
rect 1345 -221 1403 -187
rect 1345 -255 1357 -221
rect 1391 -255 1403 -221
rect 1345 -289 1403 -255
rect 1345 -323 1357 -289
rect 1391 -323 1403 -289
rect 1345 -357 1403 -323
rect 1345 -391 1357 -357
rect 1391 -391 1403 -357
rect 1345 -425 1403 -391
rect 1345 -459 1357 -425
rect 1391 -459 1403 -425
rect 1345 -493 1403 -459
rect 1345 -527 1357 -493
rect 1391 -527 1403 -493
rect 1345 -561 1403 -527
rect 1345 -595 1357 -561
rect 1391 -595 1403 -561
rect 1345 -629 1403 -595
rect 1345 -663 1357 -629
rect 1391 -663 1403 -629
rect 1345 -697 1403 -663
rect 1345 -731 1357 -697
rect 1391 -731 1403 -697
rect 1345 -765 1403 -731
rect 1345 -799 1357 -765
rect 1391 -799 1403 -765
rect 1345 -833 1403 -799
rect 1345 -867 1357 -833
rect 1391 -867 1403 -833
rect 1345 -901 1403 -867
rect 1345 -935 1357 -901
rect 1391 -935 1403 -901
rect 1345 -969 1403 -935
rect 1345 -1003 1357 -969
rect 1391 -1003 1403 -969
rect 1345 -1037 1403 -1003
rect 1345 -1071 1357 -1037
rect 1391 -1071 1403 -1037
rect 1345 -1105 1403 -1071
rect 1345 -1139 1357 -1105
rect 1391 -1139 1403 -1105
rect 1345 -1173 1403 -1139
rect 1345 -1207 1357 -1173
rect 1391 -1207 1403 -1173
rect 1345 -1241 1403 -1207
rect 1345 -1275 1357 -1241
rect 1391 -1275 1403 -1241
rect 1345 -1320 1403 -1275
rect 1803 1275 1861 1320
rect 1803 1241 1815 1275
rect 1849 1241 1861 1275
rect 1803 1207 1861 1241
rect 1803 1173 1815 1207
rect 1849 1173 1861 1207
rect 1803 1139 1861 1173
rect 1803 1105 1815 1139
rect 1849 1105 1861 1139
rect 1803 1071 1861 1105
rect 1803 1037 1815 1071
rect 1849 1037 1861 1071
rect 1803 1003 1861 1037
rect 1803 969 1815 1003
rect 1849 969 1861 1003
rect 1803 935 1861 969
rect 1803 901 1815 935
rect 1849 901 1861 935
rect 1803 867 1861 901
rect 1803 833 1815 867
rect 1849 833 1861 867
rect 1803 799 1861 833
rect 1803 765 1815 799
rect 1849 765 1861 799
rect 1803 731 1861 765
rect 1803 697 1815 731
rect 1849 697 1861 731
rect 1803 663 1861 697
rect 1803 629 1815 663
rect 1849 629 1861 663
rect 1803 595 1861 629
rect 1803 561 1815 595
rect 1849 561 1861 595
rect 1803 527 1861 561
rect 1803 493 1815 527
rect 1849 493 1861 527
rect 1803 459 1861 493
rect 1803 425 1815 459
rect 1849 425 1861 459
rect 1803 391 1861 425
rect 1803 357 1815 391
rect 1849 357 1861 391
rect 1803 323 1861 357
rect 1803 289 1815 323
rect 1849 289 1861 323
rect 1803 255 1861 289
rect 1803 221 1815 255
rect 1849 221 1861 255
rect 1803 187 1861 221
rect 1803 153 1815 187
rect 1849 153 1861 187
rect 1803 119 1861 153
rect 1803 85 1815 119
rect 1849 85 1861 119
rect 1803 51 1861 85
rect 1803 17 1815 51
rect 1849 17 1861 51
rect 1803 -17 1861 17
rect 1803 -51 1815 -17
rect 1849 -51 1861 -17
rect 1803 -85 1861 -51
rect 1803 -119 1815 -85
rect 1849 -119 1861 -85
rect 1803 -153 1861 -119
rect 1803 -187 1815 -153
rect 1849 -187 1861 -153
rect 1803 -221 1861 -187
rect 1803 -255 1815 -221
rect 1849 -255 1861 -221
rect 1803 -289 1861 -255
rect 1803 -323 1815 -289
rect 1849 -323 1861 -289
rect 1803 -357 1861 -323
rect 1803 -391 1815 -357
rect 1849 -391 1861 -357
rect 1803 -425 1861 -391
rect 1803 -459 1815 -425
rect 1849 -459 1861 -425
rect 1803 -493 1861 -459
rect 1803 -527 1815 -493
rect 1849 -527 1861 -493
rect 1803 -561 1861 -527
rect 1803 -595 1815 -561
rect 1849 -595 1861 -561
rect 1803 -629 1861 -595
rect 1803 -663 1815 -629
rect 1849 -663 1861 -629
rect 1803 -697 1861 -663
rect 1803 -731 1815 -697
rect 1849 -731 1861 -697
rect 1803 -765 1861 -731
rect 1803 -799 1815 -765
rect 1849 -799 1861 -765
rect 1803 -833 1861 -799
rect 1803 -867 1815 -833
rect 1849 -867 1861 -833
rect 1803 -901 1861 -867
rect 1803 -935 1815 -901
rect 1849 -935 1861 -901
rect 1803 -969 1861 -935
rect 1803 -1003 1815 -969
rect 1849 -1003 1861 -969
rect 1803 -1037 1861 -1003
rect 1803 -1071 1815 -1037
rect 1849 -1071 1861 -1037
rect 1803 -1105 1861 -1071
rect 1803 -1139 1815 -1105
rect 1849 -1139 1861 -1105
rect 1803 -1173 1861 -1139
rect 1803 -1207 1815 -1173
rect 1849 -1207 1861 -1173
rect 1803 -1241 1861 -1207
rect 1803 -1275 1815 -1241
rect 1849 -1275 1861 -1241
rect 1803 -1320 1861 -1275
rect 2261 1275 2319 1320
rect 2261 1241 2273 1275
rect 2307 1241 2319 1275
rect 2261 1207 2319 1241
rect 2261 1173 2273 1207
rect 2307 1173 2319 1207
rect 2261 1139 2319 1173
rect 2261 1105 2273 1139
rect 2307 1105 2319 1139
rect 2261 1071 2319 1105
rect 2261 1037 2273 1071
rect 2307 1037 2319 1071
rect 2261 1003 2319 1037
rect 2261 969 2273 1003
rect 2307 969 2319 1003
rect 2261 935 2319 969
rect 2261 901 2273 935
rect 2307 901 2319 935
rect 2261 867 2319 901
rect 2261 833 2273 867
rect 2307 833 2319 867
rect 2261 799 2319 833
rect 2261 765 2273 799
rect 2307 765 2319 799
rect 2261 731 2319 765
rect 2261 697 2273 731
rect 2307 697 2319 731
rect 2261 663 2319 697
rect 2261 629 2273 663
rect 2307 629 2319 663
rect 2261 595 2319 629
rect 2261 561 2273 595
rect 2307 561 2319 595
rect 2261 527 2319 561
rect 2261 493 2273 527
rect 2307 493 2319 527
rect 2261 459 2319 493
rect 2261 425 2273 459
rect 2307 425 2319 459
rect 2261 391 2319 425
rect 2261 357 2273 391
rect 2307 357 2319 391
rect 2261 323 2319 357
rect 2261 289 2273 323
rect 2307 289 2319 323
rect 2261 255 2319 289
rect 2261 221 2273 255
rect 2307 221 2319 255
rect 2261 187 2319 221
rect 2261 153 2273 187
rect 2307 153 2319 187
rect 2261 119 2319 153
rect 2261 85 2273 119
rect 2307 85 2319 119
rect 2261 51 2319 85
rect 2261 17 2273 51
rect 2307 17 2319 51
rect 2261 -17 2319 17
rect 2261 -51 2273 -17
rect 2307 -51 2319 -17
rect 2261 -85 2319 -51
rect 2261 -119 2273 -85
rect 2307 -119 2319 -85
rect 2261 -153 2319 -119
rect 2261 -187 2273 -153
rect 2307 -187 2319 -153
rect 2261 -221 2319 -187
rect 2261 -255 2273 -221
rect 2307 -255 2319 -221
rect 2261 -289 2319 -255
rect 2261 -323 2273 -289
rect 2307 -323 2319 -289
rect 2261 -357 2319 -323
rect 2261 -391 2273 -357
rect 2307 -391 2319 -357
rect 2261 -425 2319 -391
rect 2261 -459 2273 -425
rect 2307 -459 2319 -425
rect 2261 -493 2319 -459
rect 2261 -527 2273 -493
rect 2307 -527 2319 -493
rect 2261 -561 2319 -527
rect 2261 -595 2273 -561
rect 2307 -595 2319 -561
rect 2261 -629 2319 -595
rect 2261 -663 2273 -629
rect 2307 -663 2319 -629
rect 2261 -697 2319 -663
rect 2261 -731 2273 -697
rect 2307 -731 2319 -697
rect 2261 -765 2319 -731
rect 2261 -799 2273 -765
rect 2307 -799 2319 -765
rect 2261 -833 2319 -799
rect 2261 -867 2273 -833
rect 2307 -867 2319 -833
rect 2261 -901 2319 -867
rect 2261 -935 2273 -901
rect 2307 -935 2319 -901
rect 2261 -969 2319 -935
rect 2261 -1003 2273 -969
rect 2307 -1003 2319 -969
rect 2261 -1037 2319 -1003
rect 2261 -1071 2273 -1037
rect 2307 -1071 2319 -1037
rect 2261 -1105 2319 -1071
rect 2261 -1139 2273 -1105
rect 2307 -1139 2319 -1105
rect 2261 -1173 2319 -1139
rect 2261 -1207 2273 -1173
rect 2307 -1207 2319 -1173
rect 2261 -1241 2319 -1207
rect 2261 -1275 2273 -1241
rect 2307 -1275 2319 -1241
rect 2261 -1320 2319 -1275
<< ndiffc >>
rect -2307 1241 -2273 1275
rect -2307 1173 -2273 1207
rect -2307 1105 -2273 1139
rect -2307 1037 -2273 1071
rect -2307 969 -2273 1003
rect -2307 901 -2273 935
rect -2307 833 -2273 867
rect -2307 765 -2273 799
rect -2307 697 -2273 731
rect -2307 629 -2273 663
rect -2307 561 -2273 595
rect -2307 493 -2273 527
rect -2307 425 -2273 459
rect -2307 357 -2273 391
rect -2307 289 -2273 323
rect -2307 221 -2273 255
rect -2307 153 -2273 187
rect -2307 85 -2273 119
rect -2307 17 -2273 51
rect -2307 -51 -2273 -17
rect -2307 -119 -2273 -85
rect -2307 -187 -2273 -153
rect -2307 -255 -2273 -221
rect -2307 -323 -2273 -289
rect -2307 -391 -2273 -357
rect -2307 -459 -2273 -425
rect -2307 -527 -2273 -493
rect -2307 -595 -2273 -561
rect -2307 -663 -2273 -629
rect -2307 -731 -2273 -697
rect -2307 -799 -2273 -765
rect -2307 -867 -2273 -833
rect -2307 -935 -2273 -901
rect -2307 -1003 -2273 -969
rect -2307 -1071 -2273 -1037
rect -2307 -1139 -2273 -1105
rect -2307 -1207 -2273 -1173
rect -2307 -1275 -2273 -1241
rect -1849 1241 -1815 1275
rect -1849 1173 -1815 1207
rect -1849 1105 -1815 1139
rect -1849 1037 -1815 1071
rect -1849 969 -1815 1003
rect -1849 901 -1815 935
rect -1849 833 -1815 867
rect -1849 765 -1815 799
rect -1849 697 -1815 731
rect -1849 629 -1815 663
rect -1849 561 -1815 595
rect -1849 493 -1815 527
rect -1849 425 -1815 459
rect -1849 357 -1815 391
rect -1849 289 -1815 323
rect -1849 221 -1815 255
rect -1849 153 -1815 187
rect -1849 85 -1815 119
rect -1849 17 -1815 51
rect -1849 -51 -1815 -17
rect -1849 -119 -1815 -85
rect -1849 -187 -1815 -153
rect -1849 -255 -1815 -221
rect -1849 -323 -1815 -289
rect -1849 -391 -1815 -357
rect -1849 -459 -1815 -425
rect -1849 -527 -1815 -493
rect -1849 -595 -1815 -561
rect -1849 -663 -1815 -629
rect -1849 -731 -1815 -697
rect -1849 -799 -1815 -765
rect -1849 -867 -1815 -833
rect -1849 -935 -1815 -901
rect -1849 -1003 -1815 -969
rect -1849 -1071 -1815 -1037
rect -1849 -1139 -1815 -1105
rect -1849 -1207 -1815 -1173
rect -1849 -1275 -1815 -1241
rect -1391 1241 -1357 1275
rect -1391 1173 -1357 1207
rect -1391 1105 -1357 1139
rect -1391 1037 -1357 1071
rect -1391 969 -1357 1003
rect -1391 901 -1357 935
rect -1391 833 -1357 867
rect -1391 765 -1357 799
rect -1391 697 -1357 731
rect -1391 629 -1357 663
rect -1391 561 -1357 595
rect -1391 493 -1357 527
rect -1391 425 -1357 459
rect -1391 357 -1357 391
rect -1391 289 -1357 323
rect -1391 221 -1357 255
rect -1391 153 -1357 187
rect -1391 85 -1357 119
rect -1391 17 -1357 51
rect -1391 -51 -1357 -17
rect -1391 -119 -1357 -85
rect -1391 -187 -1357 -153
rect -1391 -255 -1357 -221
rect -1391 -323 -1357 -289
rect -1391 -391 -1357 -357
rect -1391 -459 -1357 -425
rect -1391 -527 -1357 -493
rect -1391 -595 -1357 -561
rect -1391 -663 -1357 -629
rect -1391 -731 -1357 -697
rect -1391 -799 -1357 -765
rect -1391 -867 -1357 -833
rect -1391 -935 -1357 -901
rect -1391 -1003 -1357 -969
rect -1391 -1071 -1357 -1037
rect -1391 -1139 -1357 -1105
rect -1391 -1207 -1357 -1173
rect -1391 -1275 -1357 -1241
rect -933 1241 -899 1275
rect -933 1173 -899 1207
rect -933 1105 -899 1139
rect -933 1037 -899 1071
rect -933 969 -899 1003
rect -933 901 -899 935
rect -933 833 -899 867
rect -933 765 -899 799
rect -933 697 -899 731
rect -933 629 -899 663
rect -933 561 -899 595
rect -933 493 -899 527
rect -933 425 -899 459
rect -933 357 -899 391
rect -933 289 -899 323
rect -933 221 -899 255
rect -933 153 -899 187
rect -933 85 -899 119
rect -933 17 -899 51
rect -933 -51 -899 -17
rect -933 -119 -899 -85
rect -933 -187 -899 -153
rect -933 -255 -899 -221
rect -933 -323 -899 -289
rect -933 -391 -899 -357
rect -933 -459 -899 -425
rect -933 -527 -899 -493
rect -933 -595 -899 -561
rect -933 -663 -899 -629
rect -933 -731 -899 -697
rect -933 -799 -899 -765
rect -933 -867 -899 -833
rect -933 -935 -899 -901
rect -933 -1003 -899 -969
rect -933 -1071 -899 -1037
rect -933 -1139 -899 -1105
rect -933 -1207 -899 -1173
rect -933 -1275 -899 -1241
rect -475 1241 -441 1275
rect -475 1173 -441 1207
rect -475 1105 -441 1139
rect -475 1037 -441 1071
rect -475 969 -441 1003
rect -475 901 -441 935
rect -475 833 -441 867
rect -475 765 -441 799
rect -475 697 -441 731
rect -475 629 -441 663
rect -475 561 -441 595
rect -475 493 -441 527
rect -475 425 -441 459
rect -475 357 -441 391
rect -475 289 -441 323
rect -475 221 -441 255
rect -475 153 -441 187
rect -475 85 -441 119
rect -475 17 -441 51
rect -475 -51 -441 -17
rect -475 -119 -441 -85
rect -475 -187 -441 -153
rect -475 -255 -441 -221
rect -475 -323 -441 -289
rect -475 -391 -441 -357
rect -475 -459 -441 -425
rect -475 -527 -441 -493
rect -475 -595 -441 -561
rect -475 -663 -441 -629
rect -475 -731 -441 -697
rect -475 -799 -441 -765
rect -475 -867 -441 -833
rect -475 -935 -441 -901
rect -475 -1003 -441 -969
rect -475 -1071 -441 -1037
rect -475 -1139 -441 -1105
rect -475 -1207 -441 -1173
rect -475 -1275 -441 -1241
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1139
rect -17 1037 17 1071
rect -17 969 17 1003
rect -17 901 17 935
rect -17 833 17 867
rect -17 765 17 799
rect -17 697 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -697
rect -17 -799 17 -765
rect -17 -867 17 -833
rect -17 -935 17 -901
rect -17 -1003 17 -969
rect -17 -1071 17 -1037
rect -17 -1139 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect 441 1241 475 1275
rect 441 1173 475 1207
rect 441 1105 475 1139
rect 441 1037 475 1071
rect 441 969 475 1003
rect 441 901 475 935
rect 441 833 475 867
rect 441 765 475 799
rect 441 697 475 731
rect 441 629 475 663
rect 441 561 475 595
rect 441 493 475 527
rect 441 425 475 459
rect 441 357 475 391
rect 441 289 475 323
rect 441 221 475 255
rect 441 153 475 187
rect 441 85 475 119
rect 441 17 475 51
rect 441 -51 475 -17
rect 441 -119 475 -85
rect 441 -187 475 -153
rect 441 -255 475 -221
rect 441 -323 475 -289
rect 441 -391 475 -357
rect 441 -459 475 -425
rect 441 -527 475 -493
rect 441 -595 475 -561
rect 441 -663 475 -629
rect 441 -731 475 -697
rect 441 -799 475 -765
rect 441 -867 475 -833
rect 441 -935 475 -901
rect 441 -1003 475 -969
rect 441 -1071 475 -1037
rect 441 -1139 475 -1105
rect 441 -1207 475 -1173
rect 441 -1275 475 -1241
rect 899 1241 933 1275
rect 899 1173 933 1207
rect 899 1105 933 1139
rect 899 1037 933 1071
rect 899 969 933 1003
rect 899 901 933 935
rect 899 833 933 867
rect 899 765 933 799
rect 899 697 933 731
rect 899 629 933 663
rect 899 561 933 595
rect 899 493 933 527
rect 899 425 933 459
rect 899 357 933 391
rect 899 289 933 323
rect 899 221 933 255
rect 899 153 933 187
rect 899 85 933 119
rect 899 17 933 51
rect 899 -51 933 -17
rect 899 -119 933 -85
rect 899 -187 933 -153
rect 899 -255 933 -221
rect 899 -323 933 -289
rect 899 -391 933 -357
rect 899 -459 933 -425
rect 899 -527 933 -493
rect 899 -595 933 -561
rect 899 -663 933 -629
rect 899 -731 933 -697
rect 899 -799 933 -765
rect 899 -867 933 -833
rect 899 -935 933 -901
rect 899 -1003 933 -969
rect 899 -1071 933 -1037
rect 899 -1139 933 -1105
rect 899 -1207 933 -1173
rect 899 -1275 933 -1241
rect 1357 1241 1391 1275
rect 1357 1173 1391 1207
rect 1357 1105 1391 1139
rect 1357 1037 1391 1071
rect 1357 969 1391 1003
rect 1357 901 1391 935
rect 1357 833 1391 867
rect 1357 765 1391 799
rect 1357 697 1391 731
rect 1357 629 1391 663
rect 1357 561 1391 595
rect 1357 493 1391 527
rect 1357 425 1391 459
rect 1357 357 1391 391
rect 1357 289 1391 323
rect 1357 221 1391 255
rect 1357 153 1391 187
rect 1357 85 1391 119
rect 1357 17 1391 51
rect 1357 -51 1391 -17
rect 1357 -119 1391 -85
rect 1357 -187 1391 -153
rect 1357 -255 1391 -221
rect 1357 -323 1391 -289
rect 1357 -391 1391 -357
rect 1357 -459 1391 -425
rect 1357 -527 1391 -493
rect 1357 -595 1391 -561
rect 1357 -663 1391 -629
rect 1357 -731 1391 -697
rect 1357 -799 1391 -765
rect 1357 -867 1391 -833
rect 1357 -935 1391 -901
rect 1357 -1003 1391 -969
rect 1357 -1071 1391 -1037
rect 1357 -1139 1391 -1105
rect 1357 -1207 1391 -1173
rect 1357 -1275 1391 -1241
rect 1815 1241 1849 1275
rect 1815 1173 1849 1207
rect 1815 1105 1849 1139
rect 1815 1037 1849 1071
rect 1815 969 1849 1003
rect 1815 901 1849 935
rect 1815 833 1849 867
rect 1815 765 1849 799
rect 1815 697 1849 731
rect 1815 629 1849 663
rect 1815 561 1849 595
rect 1815 493 1849 527
rect 1815 425 1849 459
rect 1815 357 1849 391
rect 1815 289 1849 323
rect 1815 221 1849 255
rect 1815 153 1849 187
rect 1815 85 1849 119
rect 1815 17 1849 51
rect 1815 -51 1849 -17
rect 1815 -119 1849 -85
rect 1815 -187 1849 -153
rect 1815 -255 1849 -221
rect 1815 -323 1849 -289
rect 1815 -391 1849 -357
rect 1815 -459 1849 -425
rect 1815 -527 1849 -493
rect 1815 -595 1849 -561
rect 1815 -663 1849 -629
rect 1815 -731 1849 -697
rect 1815 -799 1849 -765
rect 1815 -867 1849 -833
rect 1815 -935 1849 -901
rect 1815 -1003 1849 -969
rect 1815 -1071 1849 -1037
rect 1815 -1139 1849 -1105
rect 1815 -1207 1849 -1173
rect 1815 -1275 1849 -1241
rect 2273 1241 2307 1275
rect 2273 1173 2307 1207
rect 2273 1105 2307 1139
rect 2273 1037 2307 1071
rect 2273 969 2307 1003
rect 2273 901 2307 935
rect 2273 833 2307 867
rect 2273 765 2307 799
rect 2273 697 2307 731
rect 2273 629 2307 663
rect 2273 561 2307 595
rect 2273 493 2307 527
rect 2273 425 2307 459
rect 2273 357 2307 391
rect 2273 289 2307 323
rect 2273 221 2307 255
rect 2273 153 2307 187
rect 2273 85 2307 119
rect 2273 17 2307 51
rect 2273 -51 2307 -17
rect 2273 -119 2307 -85
rect 2273 -187 2307 -153
rect 2273 -255 2307 -221
rect 2273 -323 2307 -289
rect 2273 -391 2307 -357
rect 2273 -459 2307 -425
rect 2273 -527 2307 -493
rect 2273 -595 2307 -561
rect 2273 -663 2307 -629
rect 2273 -731 2307 -697
rect 2273 -799 2307 -765
rect 2273 -867 2307 -833
rect 2273 -935 2307 -901
rect 2273 -1003 2307 -969
rect 2273 -1071 2307 -1037
rect 2273 -1139 2307 -1105
rect 2273 -1207 2307 -1173
rect 2273 -1275 2307 -1241
<< psubdiff >>
rect -2421 1460 -2295 1494
rect -2261 1460 -2227 1494
rect -2193 1460 -2159 1494
rect -2125 1460 -2091 1494
rect -2057 1460 -2023 1494
rect -1989 1460 -1955 1494
rect -1921 1460 -1887 1494
rect -1853 1460 -1819 1494
rect -1785 1460 -1751 1494
rect -1717 1460 -1683 1494
rect -1649 1460 -1615 1494
rect -1581 1460 -1547 1494
rect -1513 1460 -1479 1494
rect -1445 1460 -1411 1494
rect -1377 1460 -1343 1494
rect -1309 1460 -1275 1494
rect -1241 1460 -1207 1494
rect -1173 1460 -1139 1494
rect -1105 1460 -1071 1494
rect -1037 1460 -1003 1494
rect -969 1460 -935 1494
rect -901 1460 -867 1494
rect -833 1460 -799 1494
rect -765 1460 -731 1494
rect -697 1460 -663 1494
rect -629 1460 -595 1494
rect -561 1460 -527 1494
rect -493 1460 -459 1494
rect -425 1460 -391 1494
rect -357 1460 -323 1494
rect -289 1460 -255 1494
rect -221 1460 -187 1494
rect -153 1460 -119 1494
rect -85 1460 -51 1494
rect -17 1460 17 1494
rect 51 1460 85 1494
rect 119 1460 153 1494
rect 187 1460 221 1494
rect 255 1460 289 1494
rect 323 1460 357 1494
rect 391 1460 425 1494
rect 459 1460 493 1494
rect 527 1460 561 1494
rect 595 1460 629 1494
rect 663 1460 697 1494
rect 731 1460 765 1494
rect 799 1460 833 1494
rect 867 1460 901 1494
rect 935 1460 969 1494
rect 1003 1460 1037 1494
rect 1071 1460 1105 1494
rect 1139 1460 1173 1494
rect 1207 1460 1241 1494
rect 1275 1460 1309 1494
rect 1343 1460 1377 1494
rect 1411 1460 1445 1494
rect 1479 1460 1513 1494
rect 1547 1460 1581 1494
rect 1615 1460 1649 1494
rect 1683 1460 1717 1494
rect 1751 1460 1785 1494
rect 1819 1460 1853 1494
rect 1887 1460 1921 1494
rect 1955 1460 1989 1494
rect 2023 1460 2057 1494
rect 2091 1460 2125 1494
rect 2159 1460 2193 1494
rect 2227 1460 2261 1494
rect 2295 1460 2421 1494
rect -2421 1377 -2387 1460
rect -2421 1309 -2387 1343
rect 2387 1377 2421 1460
rect -2421 1241 -2387 1275
rect -2421 1173 -2387 1207
rect -2421 1105 -2387 1139
rect -2421 1037 -2387 1071
rect -2421 969 -2387 1003
rect -2421 901 -2387 935
rect -2421 833 -2387 867
rect -2421 765 -2387 799
rect -2421 697 -2387 731
rect -2421 629 -2387 663
rect -2421 561 -2387 595
rect -2421 493 -2387 527
rect -2421 425 -2387 459
rect -2421 357 -2387 391
rect -2421 289 -2387 323
rect -2421 221 -2387 255
rect -2421 153 -2387 187
rect -2421 85 -2387 119
rect -2421 17 -2387 51
rect -2421 -51 -2387 -17
rect -2421 -119 -2387 -85
rect -2421 -187 -2387 -153
rect -2421 -255 -2387 -221
rect -2421 -323 -2387 -289
rect -2421 -391 -2387 -357
rect -2421 -459 -2387 -425
rect -2421 -527 -2387 -493
rect -2421 -595 -2387 -561
rect -2421 -663 -2387 -629
rect -2421 -731 -2387 -697
rect -2421 -799 -2387 -765
rect -2421 -867 -2387 -833
rect -2421 -935 -2387 -901
rect -2421 -1003 -2387 -969
rect -2421 -1071 -2387 -1037
rect -2421 -1139 -2387 -1105
rect -2421 -1207 -2387 -1173
rect -2421 -1275 -2387 -1241
rect -2421 -1343 -2387 -1309
rect 2387 1309 2421 1343
rect 2387 1241 2421 1275
rect 2387 1173 2421 1207
rect 2387 1105 2421 1139
rect 2387 1037 2421 1071
rect 2387 969 2421 1003
rect 2387 901 2421 935
rect 2387 833 2421 867
rect 2387 765 2421 799
rect 2387 697 2421 731
rect 2387 629 2421 663
rect 2387 561 2421 595
rect 2387 493 2421 527
rect 2387 425 2421 459
rect 2387 357 2421 391
rect 2387 289 2421 323
rect 2387 221 2421 255
rect 2387 153 2421 187
rect 2387 85 2421 119
rect 2387 17 2421 51
rect 2387 -51 2421 -17
rect 2387 -119 2421 -85
rect 2387 -187 2421 -153
rect 2387 -255 2421 -221
rect 2387 -323 2421 -289
rect 2387 -391 2421 -357
rect 2387 -459 2421 -425
rect 2387 -527 2421 -493
rect 2387 -595 2421 -561
rect 2387 -663 2421 -629
rect 2387 -731 2421 -697
rect 2387 -799 2421 -765
rect 2387 -867 2421 -833
rect 2387 -935 2421 -901
rect 2387 -1003 2421 -969
rect 2387 -1071 2421 -1037
rect 2387 -1139 2421 -1105
rect 2387 -1207 2421 -1173
rect 2387 -1275 2421 -1241
rect -2421 -1460 -2387 -1377
rect 2387 -1343 2421 -1309
rect 2387 -1460 2421 -1377
rect -2421 -1494 -2295 -1460
rect -2261 -1494 -2227 -1460
rect -2193 -1494 -2159 -1460
rect -2125 -1494 -2091 -1460
rect -2057 -1494 -2023 -1460
rect -1989 -1494 -1955 -1460
rect -1921 -1494 -1887 -1460
rect -1853 -1494 -1819 -1460
rect -1785 -1494 -1751 -1460
rect -1717 -1494 -1683 -1460
rect -1649 -1494 -1615 -1460
rect -1581 -1494 -1547 -1460
rect -1513 -1494 -1479 -1460
rect -1445 -1494 -1411 -1460
rect -1377 -1494 -1343 -1460
rect -1309 -1494 -1275 -1460
rect -1241 -1494 -1207 -1460
rect -1173 -1494 -1139 -1460
rect -1105 -1494 -1071 -1460
rect -1037 -1494 -1003 -1460
rect -969 -1494 -935 -1460
rect -901 -1494 -867 -1460
rect -833 -1494 -799 -1460
rect -765 -1494 -731 -1460
rect -697 -1494 -663 -1460
rect -629 -1494 -595 -1460
rect -561 -1494 -527 -1460
rect -493 -1494 -459 -1460
rect -425 -1494 -391 -1460
rect -357 -1494 -323 -1460
rect -289 -1494 -255 -1460
rect -221 -1494 -187 -1460
rect -153 -1494 -119 -1460
rect -85 -1494 -51 -1460
rect -17 -1494 17 -1460
rect 51 -1494 85 -1460
rect 119 -1494 153 -1460
rect 187 -1494 221 -1460
rect 255 -1494 289 -1460
rect 323 -1494 357 -1460
rect 391 -1494 425 -1460
rect 459 -1494 493 -1460
rect 527 -1494 561 -1460
rect 595 -1494 629 -1460
rect 663 -1494 697 -1460
rect 731 -1494 765 -1460
rect 799 -1494 833 -1460
rect 867 -1494 901 -1460
rect 935 -1494 969 -1460
rect 1003 -1494 1037 -1460
rect 1071 -1494 1105 -1460
rect 1139 -1494 1173 -1460
rect 1207 -1494 1241 -1460
rect 1275 -1494 1309 -1460
rect 1343 -1494 1377 -1460
rect 1411 -1494 1445 -1460
rect 1479 -1494 1513 -1460
rect 1547 -1494 1581 -1460
rect 1615 -1494 1649 -1460
rect 1683 -1494 1717 -1460
rect 1751 -1494 1785 -1460
rect 1819 -1494 1853 -1460
rect 1887 -1494 1921 -1460
rect 1955 -1494 1989 -1460
rect 2023 -1494 2057 -1460
rect 2091 -1494 2125 -1460
rect 2159 -1494 2193 -1460
rect 2227 -1494 2261 -1460
rect 2295 -1494 2421 -1460
<< psubdiffcont >>
rect -2295 1460 -2261 1494
rect -2227 1460 -2193 1494
rect -2159 1460 -2125 1494
rect -2091 1460 -2057 1494
rect -2023 1460 -1989 1494
rect -1955 1460 -1921 1494
rect -1887 1460 -1853 1494
rect -1819 1460 -1785 1494
rect -1751 1460 -1717 1494
rect -1683 1460 -1649 1494
rect -1615 1460 -1581 1494
rect -1547 1460 -1513 1494
rect -1479 1460 -1445 1494
rect -1411 1460 -1377 1494
rect -1343 1460 -1309 1494
rect -1275 1460 -1241 1494
rect -1207 1460 -1173 1494
rect -1139 1460 -1105 1494
rect -1071 1460 -1037 1494
rect -1003 1460 -969 1494
rect -935 1460 -901 1494
rect -867 1460 -833 1494
rect -799 1460 -765 1494
rect -731 1460 -697 1494
rect -663 1460 -629 1494
rect -595 1460 -561 1494
rect -527 1460 -493 1494
rect -459 1460 -425 1494
rect -391 1460 -357 1494
rect -323 1460 -289 1494
rect -255 1460 -221 1494
rect -187 1460 -153 1494
rect -119 1460 -85 1494
rect -51 1460 -17 1494
rect 17 1460 51 1494
rect 85 1460 119 1494
rect 153 1460 187 1494
rect 221 1460 255 1494
rect 289 1460 323 1494
rect 357 1460 391 1494
rect 425 1460 459 1494
rect 493 1460 527 1494
rect 561 1460 595 1494
rect 629 1460 663 1494
rect 697 1460 731 1494
rect 765 1460 799 1494
rect 833 1460 867 1494
rect 901 1460 935 1494
rect 969 1460 1003 1494
rect 1037 1460 1071 1494
rect 1105 1460 1139 1494
rect 1173 1460 1207 1494
rect 1241 1460 1275 1494
rect 1309 1460 1343 1494
rect 1377 1460 1411 1494
rect 1445 1460 1479 1494
rect 1513 1460 1547 1494
rect 1581 1460 1615 1494
rect 1649 1460 1683 1494
rect 1717 1460 1751 1494
rect 1785 1460 1819 1494
rect 1853 1460 1887 1494
rect 1921 1460 1955 1494
rect 1989 1460 2023 1494
rect 2057 1460 2091 1494
rect 2125 1460 2159 1494
rect 2193 1460 2227 1494
rect 2261 1460 2295 1494
rect -2421 1343 -2387 1377
rect 2387 1343 2421 1377
rect -2421 1275 -2387 1309
rect -2421 1207 -2387 1241
rect -2421 1139 -2387 1173
rect -2421 1071 -2387 1105
rect -2421 1003 -2387 1037
rect -2421 935 -2387 969
rect -2421 867 -2387 901
rect -2421 799 -2387 833
rect -2421 731 -2387 765
rect -2421 663 -2387 697
rect -2421 595 -2387 629
rect -2421 527 -2387 561
rect -2421 459 -2387 493
rect -2421 391 -2387 425
rect -2421 323 -2387 357
rect -2421 255 -2387 289
rect -2421 187 -2387 221
rect -2421 119 -2387 153
rect -2421 51 -2387 85
rect -2421 -17 -2387 17
rect -2421 -85 -2387 -51
rect -2421 -153 -2387 -119
rect -2421 -221 -2387 -187
rect -2421 -289 -2387 -255
rect -2421 -357 -2387 -323
rect -2421 -425 -2387 -391
rect -2421 -493 -2387 -459
rect -2421 -561 -2387 -527
rect -2421 -629 -2387 -595
rect -2421 -697 -2387 -663
rect -2421 -765 -2387 -731
rect -2421 -833 -2387 -799
rect -2421 -901 -2387 -867
rect -2421 -969 -2387 -935
rect -2421 -1037 -2387 -1003
rect -2421 -1105 -2387 -1071
rect -2421 -1173 -2387 -1139
rect -2421 -1241 -2387 -1207
rect -2421 -1309 -2387 -1275
rect 2387 1275 2421 1309
rect 2387 1207 2421 1241
rect 2387 1139 2421 1173
rect 2387 1071 2421 1105
rect 2387 1003 2421 1037
rect 2387 935 2421 969
rect 2387 867 2421 901
rect 2387 799 2421 833
rect 2387 731 2421 765
rect 2387 663 2421 697
rect 2387 595 2421 629
rect 2387 527 2421 561
rect 2387 459 2421 493
rect 2387 391 2421 425
rect 2387 323 2421 357
rect 2387 255 2421 289
rect 2387 187 2421 221
rect 2387 119 2421 153
rect 2387 51 2421 85
rect 2387 -17 2421 17
rect 2387 -85 2421 -51
rect 2387 -153 2421 -119
rect 2387 -221 2421 -187
rect 2387 -289 2421 -255
rect 2387 -357 2421 -323
rect 2387 -425 2421 -391
rect 2387 -493 2421 -459
rect 2387 -561 2421 -527
rect 2387 -629 2421 -595
rect 2387 -697 2421 -663
rect 2387 -765 2421 -731
rect 2387 -833 2421 -799
rect 2387 -901 2421 -867
rect 2387 -969 2421 -935
rect 2387 -1037 2421 -1003
rect 2387 -1105 2421 -1071
rect 2387 -1173 2421 -1139
rect 2387 -1241 2421 -1207
rect 2387 -1309 2421 -1275
rect -2421 -1377 -2387 -1343
rect 2387 -1377 2421 -1343
rect -2295 -1494 -2261 -1460
rect -2227 -1494 -2193 -1460
rect -2159 -1494 -2125 -1460
rect -2091 -1494 -2057 -1460
rect -2023 -1494 -1989 -1460
rect -1955 -1494 -1921 -1460
rect -1887 -1494 -1853 -1460
rect -1819 -1494 -1785 -1460
rect -1751 -1494 -1717 -1460
rect -1683 -1494 -1649 -1460
rect -1615 -1494 -1581 -1460
rect -1547 -1494 -1513 -1460
rect -1479 -1494 -1445 -1460
rect -1411 -1494 -1377 -1460
rect -1343 -1494 -1309 -1460
rect -1275 -1494 -1241 -1460
rect -1207 -1494 -1173 -1460
rect -1139 -1494 -1105 -1460
rect -1071 -1494 -1037 -1460
rect -1003 -1494 -969 -1460
rect -935 -1494 -901 -1460
rect -867 -1494 -833 -1460
rect -799 -1494 -765 -1460
rect -731 -1494 -697 -1460
rect -663 -1494 -629 -1460
rect -595 -1494 -561 -1460
rect -527 -1494 -493 -1460
rect -459 -1494 -425 -1460
rect -391 -1494 -357 -1460
rect -323 -1494 -289 -1460
rect -255 -1494 -221 -1460
rect -187 -1494 -153 -1460
rect -119 -1494 -85 -1460
rect -51 -1494 -17 -1460
rect 17 -1494 51 -1460
rect 85 -1494 119 -1460
rect 153 -1494 187 -1460
rect 221 -1494 255 -1460
rect 289 -1494 323 -1460
rect 357 -1494 391 -1460
rect 425 -1494 459 -1460
rect 493 -1494 527 -1460
rect 561 -1494 595 -1460
rect 629 -1494 663 -1460
rect 697 -1494 731 -1460
rect 765 -1494 799 -1460
rect 833 -1494 867 -1460
rect 901 -1494 935 -1460
rect 969 -1494 1003 -1460
rect 1037 -1494 1071 -1460
rect 1105 -1494 1139 -1460
rect 1173 -1494 1207 -1460
rect 1241 -1494 1275 -1460
rect 1309 -1494 1343 -1460
rect 1377 -1494 1411 -1460
rect 1445 -1494 1479 -1460
rect 1513 -1494 1547 -1460
rect 1581 -1494 1615 -1460
rect 1649 -1494 1683 -1460
rect 1717 -1494 1751 -1460
rect 1785 -1494 1819 -1460
rect 1853 -1494 1887 -1460
rect 1921 -1494 1955 -1460
rect 1989 -1494 2023 -1460
rect 2057 -1494 2091 -1460
rect 2125 -1494 2159 -1460
rect 2193 -1494 2227 -1460
rect 2261 -1494 2295 -1460
<< poly >>
rect -2114 1392 -2008 1408
rect -2114 1375 -2078 1392
rect -2261 1358 -2078 1375
rect -2044 1375 -2008 1392
rect -1656 1392 -1550 1408
rect -1656 1375 -1620 1392
rect -2044 1358 -1861 1375
rect -2261 1320 -1861 1358
rect -1803 1358 -1620 1375
rect -1586 1375 -1550 1392
rect -1198 1392 -1092 1408
rect -1198 1375 -1162 1392
rect -1586 1358 -1403 1375
rect -1803 1320 -1403 1358
rect -1345 1358 -1162 1375
rect -1128 1375 -1092 1392
rect -740 1392 -634 1408
rect -740 1375 -704 1392
rect -1128 1358 -945 1375
rect -1345 1320 -945 1358
rect -887 1358 -704 1375
rect -670 1375 -634 1392
rect -282 1392 -176 1408
rect -282 1375 -246 1392
rect -670 1358 -487 1375
rect -887 1320 -487 1358
rect -429 1358 -246 1375
rect -212 1375 -176 1392
rect 176 1392 282 1408
rect 176 1375 212 1392
rect -212 1358 -29 1375
rect -429 1320 -29 1358
rect 29 1358 212 1375
rect 246 1375 282 1392
rect 634 1392 740 1408
rect 634 1375 670 1392
rect 246 1358 429 1375
rect 29 1320 429 1358
rect 487 1358 670 1375
rect 704 1375 740 1392
rect 1092 1392 1198 1408
rect 1092 1375 1128 1392
rect 704 1358 887 1375
rect 487 1320 887 1358
rect 945 1358 1128 1375
rect 1162 1375 1198 1392
rect 1550 1392 1656 1408
rect 1550 1375 1586 1392
rect 1162 1358 1345 1375
rect 945 1320 1345 1358
rect 1403 1358 1586 1375
rect 1620 1375 1656 1392
rect 2008 1392 2114 1408
rect 2008 1375 2044 1392
rect 1620 1358 1803 1375
rect 1403 1320 1803 1358
rect 1861 1358 2044 1375
rect 2078 1375 2114 1392
rect 2078 1358 2261 1375
rect 1861 1320 2261 1358
rect -2261 -1358 -1861 -1320
rect -2261 -1375 -2078 -1358
rect -2114 -1392 -2078 -1375
rect -2044 -1375 -1861 -1358
rect -1803 -1358 -1403 -1320
rect -1803 -1375 -1620 -1358
rect -2044 -1392 -2008 -1375
rect -2114 -1408 -2008 -1392
rect -1656 -1392 -1620 -1375
rect -1586 -1375 -1403 -1358
rect -1345 -1358 -945 -1320
rect -1345 -1375 -1162 -1358
rect -1586 -1392 -1550 -1375
rect -1656 -1408 -1550 -1392
rect -1198 -1392 -1162 -1375
rect -1128 -1375 -945 -1358
rect -887 -1358 -487 -1320
rect -887 -1375 -704 -1358
rect -1128 -1392 -1092 -1375
rect -1198 -1408 -1092 -1392
rect -740 -1392 -704 -1375
rect -670 -1375 -487 -1358
rect -429 -1358 -29 -1320
rect -429 -1375 -246 -1358
rect -670 -1392 -634 -1375
rect -740 -1408 -634 -1392
rect -282 -1392 -246 -1375
rect -212 -1375 -29 -1358
rect 29 -1358 429 -1320
rect 29 -1375 212 -1358
rect -212 -1392 -176 -1375
rect -282 -1408 -176 -1392
rect 176 -1392 212 -1375
rect 246 -1375 429 -1358
rect 487 -1358 887 -1320
rect 487 -1375 670 -1358
rect 246 -1392 282 -1375
rect 176 -1408 282 -1392
rect 634 -1392 670 -1375
rect 704 -1375 887 -1358
rect 945 -1358 1345 -1320
rect 945 -1375 1128 -1358
rect 704 -1392 740 -1375
rect 634 -1408 740 -1392
rect 1092 -1392 1128 -1375
rect 1162 -1375 1345 -1358
rect 1403 -1358 1803 -1320
rect 1403 -1375 1586 -1358
rect 1162 -1392 1198 -1375
rect 1092 -1408 1198 -1392
rect 1550 -1392 1586 -1375
rect 1620 -1375 1803 -1358
rect 1861 -1358 2261 -1320
rect 1861 -1375 2044 -1358
rect 1620 -1392 1656 -1375
rect 1550 -1408 1656 -1392
rect 2008 -1392 2044 -1375
rect 2078 -1375 2261 -1358
rect 2078 -1392 2114 -1375
rect 2008 -1408 2114 -1392
<< polycont >>
rect -2078 1358 -2044 1392
rect -1620 1358 -1586 1392
rect -1162 1358 -1128 1392
rect -704 1358 -670 1392
rect -246 1358 -212 1392
rect 212 1358 246 1392
rect 670 1358 704 1392
rect 1128 1358 1162 1392
rect 1586 1358 1620 1392
rect 2044 1358 2078 1392
rect -2078 -1392 -2044 -1358
rect -1620 -1392 -1586 -1358
rect -1162 -1392 -1128 -1358
rect -704 -1392 -670 -1358
rect -246 -1392 -212 -1358
rect 212 -1392 246 -1358
rect 670 -1392 704 -1358
rect 1128 -1392 1162 -1358
rect 1586 -1392 1620 -1358
rect 2044 -1392 2078 -1358
<< locali >>
rect -2421 1460 -2295 1494
rect -2261 1460 -2227 1494
rect -2193 1460 -2159 1494
rect -2125 1460 -2091 1494
rect -2057 1460 -2023 1494
rect -1989 1460 -1955 1494
rect -1921 1460 -1887 1494
rect -1853 1460 -1819 1494
rect -1785 1460 -1751 1494
rect -1717 1460 -1683 1494
rect -1649 1460 -1615 1494
rect -1581 1460 -1547 1494
rect -1513 1460 -1479 1494
rect -1445 1460 -1411 1494
rect -1377 1460 -1343 1494
rect -1309 1460 -1275 1494
rect -1241 1460 -1207 1494
rect -1173 1460 -1139 1494
rect -1105 1460 -1071 1494
rect -1037 1460 -1003 1494
rect -969 1460 -935 1494
rect -901 1460 -867 1494
rect -833 1460 -799 1494
rect -765 1460 -731 1494
rect -697 1460 -663 1494
rect -629 1460 -595 1494
rect -561 1460 -527 1494
rect -493 1460 -459 1494
rect -425 1460 -391 1494
rect -357 1460 -323 1494
rect -289 1460 -255 1494
rect -221 1460 -187 1494
rect -153 1460 -119 1494
rect -85 1460 -51 1494
rect -17 1460 17 1494
rect 51 1460 85 1494
rect 119 1460 153 1494
rect 187 1460 221 1494
rect 255 1460 289 1494
rect 323 1460 357 1494
rect 391 1460 425 1494
rect 459 1460 493 1494
rect 527 1460 561 1494
rect 595 1460 629 1494
rect 663 1460 697 1494
rect 731 1460 765 1494
rect 799 1460 833 1494
rect 867 1460 901 1494
rect 935 1460 969 1494
rect 1003 1460 1037 1494
rect 1071 1460 1105 1494
rect 1139 1460 1173 1494
rect 1207 1460 1241 1494
rect 1275 1460 1309 1494
rect 1343 1460 1377 1494
rect 1411 1460 1445 1494
rect 1479 1460 1513 1494
rect 1547 1460 1581 1494
rect 1615 1460 1649 1494
rect 1683 1460 1717 1494
rect 1751 1460 1785 1494
rect 1819 1460 1853 1494
rect 1887 1460 1921 1494
rect 1955 1460 1989 1494
rect 2023 1460 2057 1494
rect 2091 1460 2125 1494
rect 2159 1460 2193 1494
rect 2227 1460 2261 1494
rect 2295 1460 2421 1494
rect -2421 1377 -2387 1460
rect -2114 1358 -2078 1392
rect -2044 1358 -2008 1392
rect -1656 1358 -1620 1392
rect -1586 1358 -1550 1392
rect -1198 1358 -1162 1392
rect -1128 1358 -1092 1392
rect -740 1358 -704 1392
rect -670 1358 -634 1392
rect -282 1358 -246 1392
rect -212 1358 -176 1392
rect 176 1358 212 1392
rect 246 1358 282 1392
rect 634 1358 670 1392
rect 704 1358 740 1392
rect 1092 1358 1128 1392
rect 1162 1358 1198 1392
rect 1550 1358 1586 1392
rect 1620 1358 1656 1392
rect 2008 1358 2044 1392
rect 2078 1358 2114 1392
rect 2387 1377 2421 1460
rect -2421 1309 -2387 1343
rect -2421 1241 -2387 1275
rect -2421 1173 -2387 1207
rect -2421 1105 -2387 1139
rect -2421 1037 -2387 1071
rect -2421 969 -2387 1003
rect -2421 901 -2387 935
rect -2421 833 -2387 867
rect -2421 765 -2387 799
rect -2421 697 -2387 731
rect -2421 629 -2387 663
rect -2421 561 -2387 595
rect -2421 493 -2387 527
rect -2421 425 -2387 459
rect -2421 357 -2387 391
rect -2421 289 -2387 323
rect -2421 221 -2387 255
rect -2421 153 -2387 187
rect -2421 85 -2387 119
rect -2421 17 -2387 51
rect -2421 -51 -2387 -17
rect -2421 -119 -2387 -85
rect -2421 -187 -2387 -153
rect -2421 -255 -2387 -221
rect -2421 -323 -2387 -289
rect -2421 -391 -2387 -357
rect -2421 -459 -2387 -425
rect -2421 -527 -2387 -493
rect -2421 -595 -2387 -561
rect -2421 -663 -2387 -629
rect -2421 -731 -2387 -697
rect -2421 -799 -2387 -765
rect -2421 -867 -2387 -833
rect -2421 -935 -2387 -901
rect -2421 -1003 -2387 -969
rect -2421 -1071 -2387 -1037
rect -2421 -1139 -2387 -1105
rect -2421 -1207 -2387 -1173
rect -2421 -1275 -2387 -1241
rect -2421 -1343 -2387 -1309
rect -2307 1277 -2273 1324
rect -2307 1207 -2273 1241
rect -2307 1139 -2273 1171
rect -2307 1071 -2273 1099
rect -2307 1003 -2273 1027
rect -2307 935 -2273 955
rect -2307 867 -2273 883
rect -2307 799 -2273 811
rect -2307 731 -2273 739
rect -2307 663 -2273 667
rect -2307 557 -2273 561
rect -2307 485 -2273 493
rect -2307 413 -2273 425
rect -2307 341 -2273 357
rect -2307 269 -2273 289
rect -2307 197 -2273 221
rect -2307 125 -2273 153
rect -2307 53 -2273 85
rect -2307 -17 -2273 17
rect -2307 -85 -2273 -53
rect -2307 -153 -2273 -125
rect -2307 -221 -2273 -197
rect -2307 -289 -2273 -269
rect -2307 -357 -2273 -341
rect -2307 -425 -2273 -413
rect -2307 -493 -2273 -485
rect -2307 -561 -2273 -557
rect -2307 -667 -2273 -663
rect -2307 -739 -2273 -731
rect -2307 -811 -2273 -799
rect -2307 -883 -2273 -867
rect -2307 -955 -2273 -935
rect -2307 -1027 -2273 -1003
rect -2307 -1099 -2273 -1071
rect -2307 -1171 -2273 -1139
rect -2307 -1241 -2273 -1207
rect -2307 -1324 -2273 -1277
rect -1849 1277 -1815 1324
rect -1849 1207 -1815 1241
rect -1849 1139 -1815 1171
rect -1849 1071 -1815 1099
rect -1849 1003 -1815 1027
rect -1849 935 -1815 955
rect -1849 867 -1815 883
rect -1849 799 -1815 811
rect -1849 731 -1815 739
rect -1849 663 -1815 667
rect -1849 557 -1815 561
rect -1849 485 -1815 493
rect -1849 413 -1815 425
rect -1849 341 -1815 357
rect -1849 269 -1815 289
rect -1849 197 -1815 221
rect -1849 125 -1815 153
rect -1849 53 -1815 85
rect -1849 -17 -1815 17
rect -1849 -85 -1815 -53
rect -1849 -153 -1815 -125
rect -1849 -221 -1815 -197
rect -1849 -289 -1815 -269
rect -1849 -357 -1815 -341
rect -1849 -425 -1815 -413
rect -1849 -493 -1815 -485
rect -1849 -561 -1815 -557
rect -1849 -667 -1815 -663
rect -1849 -739 -1815 -731
rect -1849 -811 -1815 -799
rect -1849 -883 -1815 -867
rect -1849 -955 -1815 -935
rect -1849 -1027 -1815 -1003
rect -1849 -1099 -1815 -1071
rect -1849 -1171 -1815 -1139
rect -1849 -1241 -1815 -1207
rect -1849 -1324 -1815 -1277
rect -1391 1277 -1357 1324
rect -1391 1207 -1357 1241
rect -1391 1139 -1357 1171
rect -1391 1071 -1357 1099
rect -1391 1003 -1357 1027
rect -1391 935 -1357 955
rect -1391 867 -1357 883
rect -1391 799 -1357 811
rect -1391 731 -1357 739
rect -1391 663 -1357 667
rect -1391 557 -1357 561
rect -1391 485 -1357 493
rect -1391 413 -1357 425
rect -1391 341 -1357 357
rect -1391 269 -1357 289
rect -1391 197 -1357 221
rect -1391 125 -1357 153
rect -1391 53 -1357 85
rect -1391 -17 -1357 17
rect -1391 -85 -1357 -53
rect -1391 -153 -1357 -125
rect -1391 -221 -1357 -197
rect -1391 -289 -1357 -269
rect -1391 -357 -1357 -341
rect -1391 -425 -1357 -413
rect -1391 -493 -1357 -485
rect -1391 -561 -1357 -557
rect -1391 -667 -1357 -663
rect -1391 -739 -1357 -731
rect -1391 -811 -1357 -799
rect -1391 -883 -1357 -867
rect -1391 -955 -1357 -935
rect -1391 -1027 -1357 -1003
rect -1391 -1099 -1357 -1071
rect -1391 -1171 -1357 -1139
rect -1391 -1241 -1357 -1207
rect -1391 -1324 -1357 -1277
rect -933 1277 -899 1324
rect -933 1207 -899 1241
rect -933 1139 -899 1171
rect -933 1071 -899 1099
rect -933 1003 -899 1027
rect -933 935 -899 955
rect -933 867 -899 883
rect -933 799 -899 811
rect -933 731 -899 739
rect -933 663 -899 667
rect -933 557 -899 561
rect -933 485 -899 493
rect -933 413 -899 425
rect -933 341 -899 357
rect -933 269 -899 289
rect -933 197 -899 221
rect -933 125 -899 153
rect -933 53 -899 85
rect -933 -17 -899 17
rect -933 -85 -899 -53
rect -933 -153 -899 -125
rect -933 -221 -899 -197
rect -933 -289 -899 -269
rect -933 -357 -899 -341
rect -933 -425 -899 -413
rect -933 -493 -899 -485
rect -933 -561 -899 -557
rect -933 -667 -899 -663
rect -933 -739 -899 -731
rect -933 -811 -899 -799
rect -933 -883 -899 -867
rect -933 -955 -899 -935
rect -933 -1027 -899 -1003
rect -933 -1099 -899 -1071
rect -933 -1171 -899 -1139
rect -933 -1241 -899 -1207
rect -933 -1324 -899 -1277
rect -475 1277 -441 1324
rect -475 1207 -441 1241
rect -475 1139 -441 1171
rect -475 1071 -441 1099
rect -475 1003 -441 1027
rect -475 935 -441 955
rect -475 867 -441 883
rect -475 799 -441 811
rect -475 731 -441 739
rect -475 663 -441 667
rect -475 557 -441 561
rect -475 485 -441 493
rect -475 413 -441 425
rect -475 341 -441 357
rect -475 269 -441 289
rect -475 197 -441 221
rect -475 125 -441 153
rect -475 53 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -53
rect -475 -153 -441 -125
rect -475 -221 -441 -197
rect -475 -289 -441 -269
rect -475 -357 -441 -341
rect -475 -425 -441 -413
rect -475 -493 -441 -485
rect -475 -561 -441 -557
rect -475 -667 -441 -663
rect -475 -739 -441 -731
rect -475 -811 -441 -799
rect -475 -883 -441 -867
rect -475 -955 -441 -935
rect -475 -1027 -441 -1003
rect -475 -1099 -441 -1071
rect -475 -1171 -441 -1139
rect -475 -1241 -441 -1207
rect -475 -1324 -441 -1277
rect -17 1277 17 1324
rect -17 1207 17 1241
rect -17 1139 17 1171
rect -17 1071 17 1099
rect -17 1003 17 1027
rect -17 935 17 955
rect -17 867 17 883
rect -17 799 17 811
rect -17 731 17 739
rect -17 663 17 667
rect -17 557 17 561
rect -17 485 17 493
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -493 17 -485
rect -17 -561 17 -557
rect -17 -667 17 -663
rect -17 -739 17 -731
rect -17 -811 17 -799
rect -17 -883 17 -867
rect -17 -955 17 -935
rect -17 -1027 17 -1003
rect -17 -1099 17 -1071
rect -17 -1171 17 -1139
rect -17 -1241 17 -1207
rect -17 -1324 17 -1277
rect 441 1277 475 1324
rect 441 1207 475 1241
rect 441 1139 475 1171
rect 441 1071 475 1099
rect 441 1003 475 1027
rect 441 935 475 955
rect 441 867 475 883
rect 441 799 475 811
rect 441 731 475 739
rect 441 663 475 667
rect 441 557 475 561
rect 441 485 475 493
rect 441 413 475 425
rect 441 341 475 357
rect 441 269 475 289
rect 441 197 475 221
rect 441 125 475 153
rect 441 53 475 85
rect 441 -17 475 17
rect 441 -85 475 -53
rect 441 -153 475 -125
rect 441 -221 475 -197
rect 441 -289 475 -269
rect 441 -357 475 -341
rect 441 -425 475 -413
rect 441 -493 475 -485
rect 441 -561 475 -557
rect 441 -667 475 -663
rect 441 -739 475 -731
rect 441 -811 475 -799
rect 441 -883 475 -867
rect 441 -955 475 -935
rect 441 -1027 475 -1003
rect 441 -1099 475 -1071
rect 441 -1171 475 -1139
rect 441 -1241 475 -1207
rect 441 -1324 475 -1277
rect 899 1277 933 1324
rect 899 1207 933 1241
rect 899 1139 933 1171
rect 899 1071 933 1099
rect 899 1003 933 1027
rect 899 935 933 955
rect 899 867 933 883
rect 899 799 933 811
rect 899 731 933 739
rect 899 663 933 667
rect 899 557 933 561
rect 899 485 933 493
rect 899 413 933 425
rect 899 341 933 357
rect 899 269 933 289
rect 899 197 933 221
rect 899 125 933 153
rect 899 53 933 85
rect 899 -17 933 17
rect 899 -85 933 -53
rect 899 -153 933 -125
rect 899 -221 933 -197
rect 899 -289 933 -269
rect 899 -357 933 -341
rect 899 -425 933 -413
rect 899 -493 933 -485
rect 899 -561 933 -557
rect 899 -667 933 -663
rect 899 -739 933 -731
rect 899 -811 933 -799
rect 899 -883 933 -867
rect 899 -955 933 -935
rect 899 -1027 933 -1003
rect 899 -1099 933 -1071
rect 899 -1171 933 -1139
rect 899 -1241 933 -1207
rect 899 -1324 933 -1277
rect 1357 1277 1391 1324
rect 1357 1207 1391 1241
rect 1357 1139 1391 1171
rect 1357 1071 1391 1099
rect 1357 1003 1391 1027
rect 1357 935 1391 955
rect 1357 867 1391 883
rect 1357 799 1391 811
rect 1357 731 1391 739
rect 1357 663 1391 667
rect 1357 557 1391 561
rect 1357 485 1391 493
rect 1357 413 1391 425
rect 1357 341 1391 357
rect 1357 269 1391 289
rect 1357 197 1391 221
rect 1357 125 1391 153
rect 1357 53 1391 85
rect 1357 -17 1391 17
rect 1357 -85 1391 -53
rect 1357 -153 1391 -125
rect 1357 -221 1391 -197
rect 1357 -289 1391 -269
rect 1357 -357 1391 -341
rect 1357 -425 1391 -413
rect 1357 -493 1391 -485
rect 1357 -561 1391 -557
rect 1357 -667 1391 -663
rect 1357 -739 1391 -731
rect 1357 -811 1391 -799
rect 1357 -883 1391 -867
rect 1357 -955 1391 -935
rect 1357 -1027 1391 -1003
rect 1357 -1099 1391 -1071
rect 1357 -1171 1391 -1139
rect 1357 -1241 1391 -1207
rect 1357 -1324 1391 -1277
rect 1815 1277 1849 1324
rect 1815 1207 1849 1241
rect 1815 1139 1849 1171
rect 1815 1071 1849 1099
rect 1815 1003 1849 1027
rect 1815 935 1849 955
rect 1815 867 1849 883
rect 1815 799 1849 811
rect 1815 731 1849 739
rect 1815 663 1849 667
rect 1815 557 1849 561
rect 1815 485 1849 493
rect 1815 413 1849 425
rect 1815 341 1849 357
rect 1815 269 1849 289
rect 1815 197 1849 221
rect 1815 125 1849 153
rect 1815 53 1849 85
rect 1815 -17 1849 17
rect 1815 -85 1849 -53
rect 1815 -153 1849 -125
rect 1815 -221 1849 -197
rect 1815 -289 1849 -269
rect 1815 -357 1849 -341
rect 1815 -425 1849 -413
rect 1815 -493 1849 -485
rect 1815 -561 1849 -557
rect 1815 -667 1849 -663
rect 1815 -739 1849 -731
rect 1815 -811 1849 -799
rect 1815 -883 1849 -867
rect 1815 -955 1849 -935
rect 1815 -1027 1849 -1003
rect 1815 -1099 1849 -1071
rect 1815 -1171 1849 -1139
rect 1815 -1241 1849 -1207
rect 1815 -1324 1849 -1277
rect 2273 1277 2307 1324
rect 2273 1207 2307 1241
rect 2273 1139 2307 1171
rect 2273 1071 2307 1099
rect 2273 1003 2307 1027
rect 2273 935 2307 955
rect 2273 867 2307 883
rect 2273 799 2307 811
rect 2273 731 2307 739
rect 2273 663 2307 667
rect 2273 557 2307 561
rect 2273 485 2307 493
rect 2273 413 2307 425
rect 2273 341 2307 357
rect 2273 269 2307 289
rect 2273 197 2307 221
rect 2273 125 2307 153
rect 2273 53 2307 85
rect 2273 -17 2307 17
rect 2273 -85 2307 -53
rect 2273 -153 2307 -125
rect 2273 -221 2307 -197
rect 2273 -289 2307 -269
rect 2273 -357 2307 -341
rect 2273 -425 2307 -413
rect 2273 -493 2307 -485
rect 2273 -561 2307 -557
rect 2273 -667 2307 -663
rect 2273 -739 2307 -731
rect 2273 -811 2307 -799
rect 2273 -883 2307 -867
rect 2273 -955 2307 -935
rect 2273 -1027 2307 -1003
rect 2273 -1099 2307 -1071
rect 2273 -1171 2307 -1139
rect 2273 -1241 2307 -1207
rect 2273 -1324 2307 -1277
rect 2387 1309 2421 1343
rect 2387 1241 2421 1275
rect 2387 1173 2421 1207
rect 2387 1105 2421 1139
rect 2387 1037 2421 1071
rect 2387 969 2421 1003
rect 2387 901 2421 935
rect 2387 833 2421 867
rect 2387 765 2421 799
rect 2387 697 2421 731
rect 2387 629 2421 663
rect 2387 561 2421 595
rect 2387 493 2421 527
rect 2387 425 2421 459
rect 2387 357 2421 391
rect 2387 289 2421 323
rect 2387 221 2421 255
rect 2387 153 2421 187
rect 2387 85 2421 119
rect 2387 17 2421 51
rect 2387 -51 2421 -17
rect 2387 -119 2421 -85
rect 2387 -187 2421 -153
rect 2387 -255 2421 -221
rect 2387 -323 2421 -289
rect 2387 -391 2421 -357
rect 2387 -459 2421 -425
rect 2387 -527 2421 -493
rect 2387 -595 2421 -561
rect 2387 -663 2421 -629
rect 2387 -731 2421 -697
rect 2387 -799 2421 -765
rect 2387 -867 2421 -833
rect 2387 -935 2421 -901
rect 2387 -1003 2421 -969
rect 2387 -1071 2421 -1037
rect 2387 -1139 2421 -1105
rect 2387 -1207 2421 -1173
rect 2387 -1275 2421 -1241
rect 2387 -1343 2421 -1309
rect -2421 -1460 -2387 -1377
rect -2114 -1392 -2078 -1358
rect -2044 -1392 -2008 -1358
rect -1656 -1392 -1620 -1358
rect -1586 -1392 -1550 -1358
rect -1198 -1392 -1162 -1358
rect -1128 -1392 -1092 -1358
rect -740 -1392 -704 -1358
rect -670 -1392 -634 -1358
rect -282 -1392 -246 -1358
rect -212 -1392 -176 -1358
rect 176 -1392 212 -1358
rect 246 -1392 282 -1358
rect 634 -1392 670 -1358
rect 704 -1392 740 -1358
rect 1092 -1392 1128 -1358
rect 1162 -1392 1198 -1358
rect 1550 -1392 1586 -1358
rect 1620 -1392 1656 -1358
rect 2008 -1392 2044 -1358
rect 2078 -1392 2114 -1358
rect 2387 -1460 2421 -1377
rect -2421 -1494 -2357 -1460
rect -2323 -1494 -2295 -1460
rect -2251 -1494 -2227 -1460
rect -2179 -1494 -2159 -1460
rect -2107 -1494 -2091 -1460
rect -2035 -1494 -2023 -1460
rect -1963 -1494 -1955 -1460
rect -1891 -1494 -1887 -1460
rect -1785 -1494 -1781 -1460
rect -1717 -1494 -1709 -1460
rect -1649 -1494 -1637 -1460
rect -1581 -1494 -1565 -1460
rect -1513 -1494 -1493 -1460
rect -1445 -1494 -1421 -1460
rect -1377 -1494 -1349 -1460
rect -1309 -1494 -1277 -1460
rect -1241 -1494 -1207 -1460
rect -1171 -1494 -1139 -1460
rect -1099 -1494 -1071 -1460
rect -1027 -1494 -1003 -1460
rect -955 -1494 -935 -1460
rect -883 -1494 -867 -1460
rect -811 -1494 -799 -1460
rect -739 -1494 -731 -1460
rect -667 -1494 -663 -1460
rect -561 -1494 -557 -1460
rect -493 -1494 -485 -1460
rect -425 -1494 -413 -1460
rect -357 -1494 -341 -1460
rect -289 -1494 -269 -1460
rect -221 -1494 -197 -1460
rect -153 -1494 -125 -1460
rect -85 -1494 -53 -1460
rect -17 -1494 17 -1460
rect 53 -1494 85 -1460
rect 125 -1494 153 -1460
rect 197 -1494 221 -1460
rect 269 -1494 289 -1460
rect 341 -1494 357 -1460
rect 413 -1494 425 -1460
rect 485 -1494 493 -1460
rect 557 -1494 561 -1460
rect 663 -1494 667 -1460
rect 731 -1494 739 -1460
rect 799 -1494 811 -1460
rect 867 -1494 883 -1460
rect 935 -1494 955 -1460
rect 1003 -1494 1027 -1460
rect 1071 -1494 1099 -1460
rect 1139 -1494 1171 -1460
rect 1207 -1494 1241 -1460
rect 1277 -1494 1309 -1460
rect 1349 -1494 1377 -1460
rect 1421 -1494 1445 -1460
rect 1493 -1494 1513 -1460
rect 1565 -1494 1581 -1460
rect 1637 -1494 1649 -1460
rect 1709 -1494 1717 -1460
rect 1781 -1494 1785 -1460
rect 1887 -1494 1891 -1460
rect 1955 -1494 1963 -1460
rect 2023 -1494 2035 -1460
rect 2091 -1494 2107 -1460
rect 2159 -1494 2179 -1460
rect 2227 -1494 2251 -1460
rect 2295 -1494 2323 -1460
rect 2357 -1494 2421 -1460
<< viali >>
rect -2307 1275 -2273 1277
rect -2307 1243 -2273 1275
rect -2307 1173 -2273 1205
rect -2307 1171 -2273 1173
rect -2307 1105 -2273 1133
rect -2307 1099 -2273 1105
rect -2307 1037 -2273 1061
rect -2307 1027 -2273 1037
rect -2307 969 -2273 989
rect -2307 955 -2273 969
rect -2307 901 -2273 917
rect -2307 883 -2273 901
rect -2307 833 -2273 845
rect -2307 811 -2273 833
rect -2307 765 -2273 773
rect -2307 739 -2273 765
rect -2307 697 -2273 701
rect -2307 667 -2273 697
rect -2307 595 -2273 629
rect -2307 527 -2273 557
rect -2307 523 -2273 527
rect -2307 459 -2273 485
rect -2307 451 -2273 459
rect -2307 391 -2273 413
rect -2307 379 -2273 391
rect -2307 323 -2273 341
rect -2307 307 -2273 323
rect -2307 255 -2273 269
rect -2307 235 -2273 255
rect -2307 187 -2273 197
rect -2307 163 -2273 187
rect -2307 119 -2273 125
rect -2307 91 -2273 119
rect -2307 51 -2273 53
rect -2307 19 -2273 51
rect -2307 -51 -2273 -19
rect -2307 -53 -2273 -51
rect -2307 -119 -2273 -91
rect -2307 -125 -2273 -119
rect -2307 -187 -2273 -163
rect -2307 -197 -2273 -187
rect -2307 -255 -2273 -235
rect -2307 -269 -2273 -255
rect -2307 -323 -2273 -307
rect -2307 -341 -2273 -323
rect -2307 -391 -2273 -379
rect -2307 -413 -2273 -391
rect -2307 -459 -2273 -451
rect -2307 -485 -2273 -459
rect -2307 -527 -2273 -523
rect -2307 -557 -2273 -527
rect -2307 -629 -2273 -595
rect -2307 -697 -2273 -667
rect -2307 -701 -2273 -697
rect -2307 -765 -2273 -739
rect -2307 -773 -2273 -765
rect -2307 -833 -2273 -811
rect -2307 -845 -2273 -833
rect -2307 -901 -2273 -883
rect -2307 -917 -2273 -901
rect -2307 -969 -2273 -955
rect -2307 -989 -2273 -969
rect -2307 -1037 -2273 -1027
rect -2307 -1061 -2273 -1037
rect -2307 -1105 -2273 -1099
rect -2307 -1133 -2273 -1105
rect -2307 -1173 -2273 -1171
rect -2307 -1205 -2273 -1173
rect -2307 -1275 -2273 -1243
rect -2307 -1277 -2273 -1275
rect -1849 1275 -1815 1277
rect -1849 1243 -1815 1275
rect -1849 1173 -1815 1205
rect -1849 1171 -1815 1173
rect -1849 1105 -1815 1133
rect -1849 1099 -1815 1105
rect -1849 1037 -1815 1061
rect -1849 1027 -1815 1037
rect -1849 969 -1815 989
rect -1849 955 -1815 969
rect -1849 901 -1815 917
rect -1849 883 -1815 901
rect -1849 833 -1815 845
rect -1849 811 -1815 833
rect -1849 765 -1815 773
rect -1849 739 -1815 765
rect -1849 697 -1815 701
rect -1849 667 -1815 697
rect -1849 595 -1815 629
rect -1849 527 -1815 557
rect -1849 523 -1815 527
rect -1849 459 -1815 485
rect -1849 451 -1815 459
rect -1849 391 -1815 413
rect -1849 379 -1815 391
rect -1849 323 -1815 341
rect -1849 307 -1815 323
rect -1849 255 -1815 269
rect -1849 235 -1815 255
rect -1849 187 -1815 197
rect -1849 163 -1815 187
rect -1849 119 -1815 125
rect -1849 91 -1815 119
rect -1849 51 -1815 53
rect -1849 19 -1815 51
rect -1849 -51 -1815 -19
rect -1849 -53 -1815 -51
rect -1849 -119 -1815 -91
rect -1849 -125 -1815 -119
rect -1849 -187 -1815 -163
rect -1849 -197 -1815 -187
rect -1849 -255 -1815 -235
rect -1849 -269 -1815 -255
rect -1849 -323 -1815 -307
rect -1849 -341 -1815 -323
rect -1849 -391 -1815 -379
rect -1849 -413 -1815 -391
rect -1849 -459 -1815 -451
rect -1849 -485 -1815 -459
rect -1849 -527 -1815 -523
rect -1849 -557 -1815 -527
rect -1849 -629 -1815 -595
rect -1849 -697 -1815 -667
rect -1849 -701 -1815 -697
rect -1849 -765 -1815 -739
rect -1849 -773 -1815 -765
rect -1849 -833 -1815 -811
rect -1849 -845 -1815 -833
rect -1849 -901 -1815 -883
rect -1849 -917 -1815 -901
rect -1849 -969 -1815 -955
rect -1849 -989 -1815 -969
rect -1849 -1037 -1815 -1027
rect -1849 -1061 -1815 -1037
rect -1849 -1105 -1815 -1099
rect -1849 -1133 -1815 -1105
rect -1849 -1173 -1815 -1171
rect -1849 -1205 -1815 -1173
rect -1849 -1275 -1815 -1243
rect -1849 -1277 -1815 -1275
rect -1391 1275 -1357 1277
rect -1391 1243 -1357 1275
rect -1391 1173 -1357 1205
rect -1391 1171 -1357 1173
rect -1391 1105 -1357 1133
rect -1391 1099 -1357 1105
rect -1391 1037 -1357 1061
rect -1391 1027 -1357 1037
rect -1391 969 -1357 989
rect -1391 955 -1357 969
rect -1391 901 -1357 917
rect -1391 883 -1357 901
rect -1391 833 -1357 845
rect -1391 811 -1357 833
rect -1391 765 -1357 773
rect -1391 739 -1357 765
rect -1391 697 -1357 701
rect -1391 667 -1357 697
rect -1391 595 -1357 629
rect -1391 527 -1357 557
rect -1391 523 -1357 527
rect -1391 459 -1357 485
rect -1391 451 -1357 459
rect -1391 391 -1357 413
rect -1391 379 -1357 391
rect -1391 323 -1357 341
rect -1391 307 -1357 323
rect -1391 255 -1357 269
rect -1391 235 -1357 255
rect -1391 187 -1357 197
rect -1391 163 -1357 187
rect -1391 119 -1357 125
rect -1391 91 -1357 119
rect -1391 51 -1357 53
rect -1391 19 -1357 51
rect -1391 -51 -1357 -19
rect -1391 -53 -1357 -51
rect -1391 -119 -1357 -91
rect -1391 -125 -1357 -119
rect -1391 -187 -1357 -163
rect -1391 -197 -1357 -187
rect -1391 -255 -1357 -235
rect -1391 -269 -1357 -255
rect -1391 -323 -1357 -307
rect -1391 -341 -1357 -323
rect -1391 -391 -1357 -379
rect -1391 -413 -1357 -391
rect -1391 -459 -1357 -451
rect -1391 -485 -1357 -459
rect -1391 -527 -1357 -523
rect -1391 -557 -1357 -527
rect -1391 -629 -1357 -595
rect -1391 -697 -1357 -667
rect -1391 -701 -1357 -697
rect -1391 -765 -1357 -739
rect -1391 -773 -1357 -765
rect -1391 -833 -1357 -811
rect -1391 -845 -1357 -833
rect -1391 -901 -1357 -883
rect -1391 -917 -1357 -901
rect -1391 -969 -1357 -955
rect -1391 -989 -1357 -969
rect -1391 -1037 -1357 -1027
rect -1391 -1061 -1357 -1037
rect -1391 -1105 -1357 -1099
rect -1391 -1133 -1357 -1105
rect -1391 -1173 -1357 -1171
rect -1391 -1205 -1357 -1173
rect -1391 -1275 -1357 -1243
rect -1391 -1277 -1357 -1275
rect -933 1275 -899 1277
rect -933 1243 -899 1275
rect -933 1173 -899 1205
rect -933 1171 -899 1173
rect -933 1105 -899 1133
rect -933 1099 -899 1105
rect -933 1037 -899 1061
rect -933 1027 -899 1037
rect -933 969 -899 989
rect -933 955 -899 969
rect -933 901 -899 917
rect -933 883 -899 901
rect -933 833 -899 845
rect -933 811 -899 833
rect -933 765 -899 773
rect -933 739 -899 765
rect -933 697 -899 701
rect -933 667 -899 697
rect -933 595 -899 629
rect -933 527 -899 557
rect -933 523 -899 527
rect -933 459 -899 485
rect -933 451 -899 459
rect -933 391 -899 413
rect -933 379 -899 391
rect -933 323 -899 341
rect -933 307 -899 323
rect -933 255 -899 269
rect -933 235 -899 255
rect -933 187 -899 197
rect -933 163 -899 187
rect -933 119 -899 125
rect -933 91 -899 119
rect -933 51 -899 53
rect -933 19 -899 51
rect -933 -51 -899 -19
rect -933 -53 -899 -51
rect -933 -119 -899 -91
rect -933 -125 -899 -119
rect -933 -187 -899 -163
rect -933 -197 -899 -187
rect -933 -255 -899 -235
rect -933 -269 -899 -255
rect -933 -323 -899 -307
rect -933 -341 -899 -323
rect -933 -391 -899 -379
rect -933 -413 -899 -391
rect -933 -459 -899 -451
rect -933 -485 -899 -459
rect -933 -527 -899 -523
rect -933 -557 -899 -527
rect -933 -629 -899 -595
rect -933 -697 -899 -667
rect -933 -701 -899 -697
rect -933 -765 -899 -739
rect -933 -773 -899 -765
rect -933 -833 -899 -811
rect -933 -845 -899 -833
rect -933 -901 -899 -883
rect -933 -917 -899 -901
rect -933 -969 -899 -955
rect -933 -989 -899 -969
rect -933 -1037 -899 -1027
rect -933 -1061 -899 -1037
rect -933 -1105 -899 -1099
rect -933 -1133 -899 -1105
rect -933 -1173 -899 -1171
rect -933 -1205 -899 -1173
rect -933 -1275 -899 -1243
rect -933 -1277 -899 -1275
rect -475 1275 -441 1277
rect -475 1243 -441 1275
rect -475 1173 -441 1205
rect -475 1171 -441 1173
rect -475 1105 -441 1133
rect -475 1099 -441 1105
rect -475 1037 -441 1061
rect -475 1027 -441 1037
rect -475 969 -441 989
rect -475 955 -441 969
rect -475 901 -441 917
rect -475 883 -441 901
rect -475 833 -441 845
rect -475 811 -441 833
rect -475 765 -441 773
rect -475 739 -441 765
rect -475 697 -441 701
rect -475 667 -441 697
rect -475 595 -441 629
rect -475 527 -441 557
rect -475 523 -441 527
rect -475 459 -441 485
rect -475 451 -441 459
rect -475 391 -441 413
rect -475 379 -441 391
rect -475 323 -441 341
rect -475 307 -441 323
rect -475 255 -441 269
rect -475 235 -441 255
rect -475 187 -441 197
rect -475 163 -441 187
rect -475 119 -441 125
rect -475 91 -441 119
rect -475 51 -441 53
rect -475 19 -441 51
rect -475 -51 -441 -19
rect -475 -53 -441 -51
rect -475 -119 -441 -91
rect -475 -125 -441 -119
rect -475 -187 -441 -163
rect -475 -197 -441 -187
rect -475 -255 -441 -235
rect -475 -269 -441 -255
rect -475 -323 -441 -307
rect -475 -341 -441 -323
rect -475 -391 -441 -379
rect -475 -413 -441 -391
rect -475 -459 -441 -451
rect -475 -485 -441 -459
rect -475 -527 -441 -523
rect -475 -557 -441 -527
rect -475 -629 -441 -595
rect -475 -697 -441 -667
rect -475 -701 -441 -697
rect -475 -765 -441 -739
rect -475 -773 -441 -765
rect -475 -833 -441 -811
rect -475 -845 -441 -833
rect -475 -901 -441 -883
rect -475 -917 -441 -901
rect -475 -969 -441 -955
rect -475 -989 -441 -969
rect -475 -1037 -441 -1027
rect -475 -1061 -441 -1037
rect -475 -1105 -441 -1099
rect -475 -1133 -441 -1105
rect -475 -1173 -441 -1171
rect -475 -1205 -441 -1173
rect -475 -1275 -441 -1243
rect -475 -1277 -441 -1275
rect -17 1275 17 1277
rect -17 1243 17 1275
rect -17 1173 17 1205
rect -17 1171 17 1173
rect -17 1105 17 1133
rect -17 1099 17 1105
rect -17 1037 17 1061
rect -17 1027 17 1037
rect -17 969 17 989
rect -17 955 17 969
rect -17 901 17 917
rect -17 883 17 901
rect -17 833 17 845
rect -17 811 17 833
rect -17 765 17 773
rect -17 739 17 765
rect -17 697 17 701
rect -17 667 17 697
rect -17 595 17 629
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -667
rect -17 -701 17 -697
rect -17 -765 17 -739
rect -17 -773 17 -765
rect -17 -833 17 -811
rect -17 -845 17 -833
rect -17 -901 17 -883
rect -17 -917 17 -901
rect -17 -969 17 -955
rect -17 -989 17 -969
rect -17 -1037 17 -1027
rect -17 -1061 17 -1037
rect -17 -1105 17 -1099
rect -17 -1133 17 -1105
rect -17 -1173 17 -1171
rect -17 -1205 17 -1173
rect -17 -1275 17 -1243
rect -17 -1277 17 -1275
rect 441 1275 475 1277
rect 441 1243 475 1275
rect 441 1173 475 1205
rect 441 1171 475 1173
rect 441 1105 475 1133
rect 441 1099 475 1105
rect 441 1037 475 1061
rect 441 1027 475 1037
rect 441 969 475 989
rect 441 955 475 969
rect 441 901 475 917
rect 441 883 475 901
rect 441 833 475 845
rect 441 811 475 833
rect 441 765 475 773
rect 441 739 475 765
rect 441 697 475 701
rect 441 667 475 697
rect 441 595 475 629
rect 441 527 475 557
rect 441 523 475 527
rect 441 459 475 485
rect 441 451 475 459
rect 441 391 475 413
rect 441 379 475 391
rect 441 323 475 341
rect 441 307 475 323
rect 441 255 475 269
rect 441 235 475 255
rect 441 187 475 197
rect 441 163 475 187
rect 441 119 475 125
rect 441 91 475 119
rect 441 51 475 53
rect 441 19 475 51
rect 441 -51 475 -19
rect 441 -53 475 -51
rect 441 -119 475 -91
rect 441 -125 475 -119
rect 441 -187 475 -163
rect 441 -197 475 -187
rect 441 -255 475 -235
rect 441 -269 475 -255
rect 441 -323 475 -307
rect 441 -341 475 -323
rect 441 -391 475 -379
rect 441 -413 475 -391
rect 441 -459 475 -451
rect 441 -485 475 -459
rect 441 -527 475 -523
rect 441 -557 475 -527
rect 441 -629 475 -595
rect 441 -697 475 -667
rect 441 -701 475 -697
rect 441 -765 475 -739
rect 441 -773 475 -765
rect 441 -833 475 -811
rect 441 -845 475 -833
rect 441 -901 475 -883
rect 441 -917 475 -901
rect 441 -969 475 -955
rect 441 -989 475 -969
rect 441 -1037 475 -1027
rect 441 -1061 475 -1037
rect 441 -1105 475 -1099
rect 441 -1133 475 -1105
rect 441 -1173 475 -1171
rect 441 -1205 475 -1173
rect 441 -1275 475 -1243
rect 441 -1277 475 -1275
rect 899 1275 933 1277
rect 899 1243 933 1275
rect 899 1173 933 1205
rect 899 1171 933 1173
rect 899 1105 933 1133
rect 899 1099 933 1105
rect 899 1037 933 1061
rect 899 1027 933 1037
rect 899 969 933 989
rect 899 955 933 969
rect 899 901 933 917
rect 899 883 933 901
rect 899 833 933 845
rect 899 811 933 833
rect 899 765 933 773
rect 899 739 933 765
rect 899 697 933 701
rect 899 667 933 697
rect 899 595 933 629
rect 899 527 933 557
rect 899 523 933 527
rect 899 459 933 485
rect 899 451 933 459
rect 899 391 933 413
rect 899 379 933 391
rect 899 323 933 341
rect 899 307 933 323
rect 899 255 933 269
rect 899 235 933 255
rect 899 187 933 197
rect 899 163 933 187
rect 899 119 933 125
rect 899 91 933 119
rect 899 51 933 53
rect 899 19 933 51
rect 899 -51 933 -19
rect 899 -53 933 -51
rect 899 -119 933 -91
rect 899 -125 933 -119
rect 899 -187 933 -163
rect 899 -197 933 -187
rect 899 -255 933 -235
rect 899 -269 933 -255
rect 899 -323 933 -307
rect 899 -341 933 -323
rect 899 -391 933 -379
rect 899 -413 933 -391
rect 899 -459 933 -451
rect 899 -485 933 -459
rect 899 -527 933 -523
rect 899 -557 933 -527
rect 899 -629 933 -595
rect 899 -697 933 -667
rect 899 -701 933 -697
rect 899 -765 933 -739
rect 899 -773 933 -765
rect 899 -833 933 -811
rect 899 -845 933 -833
rect 899 -901 933 -883
rect 899 -917 933 -901
rect 899 -969 933 -955
rect 899 -989 933 -969
rect 899 -1037 933 -1027
rect 899 -1061 933 -1037
rect 899 -1105 933 -1099
rect 899 -1133 933 -1105
rect 899 -1173 933 -1171
rect 899 -1205 933 -1173
rect 899 -1275 933 -1243
rect 899 -1277 933 -1275
rect 1357 1275 1391 1277
rect 1357 1243 1391 1275
rect 1357 1173 1391 1205
rect 1357 1171 1391 1173
rect 1357 1105 1391 1133
rect 1357 1099 1391 1105
rect 1357 1037 1391 1061
rect 1357 1027 1391 1037
rect 1357 969 1391 989
rect 1357 955 1391 969
rect 1357 901 1391 917
rect 1357 883 1391 901
rect 1357 833 1391 845
rect 1357 811 1391 833
rect 1357 765 1391 773
rect 1357 739 1391 765
rect 1357 697 1391 701
rect 1357 667 1391 697
rect 1357 595 1391 629
rect 1357 527 1391 557
rect 1357 523 1391 527
rect 1357 459 1391 485
rect 1357 451 1391 459
rect 1357 391 1391 413
rect 1357 379 1391 391
rect 1357 323 1391 341
rect 1357 307 1391 323
rect 1357 255 1391 269
rect 1357 235 1391 255
rect 1357 187 1391 197
rect 1357 163 1391 187
rect 1357 119 1391 125
rect 1357 91 1391 119
rect 1357 51 1391 53
rect 1357 19 1391 51
rect 1357 -51 1391 -19
rect 1357 -53 1391 -51
rect 1357 -119 1391 -91
rect 1357 -125 1391 -119
rect 1357 -187 1391 -163
rect 1357 -197 1391 -187
rect 1357 -255 1391 -235
rect 1357 -269 1391 -255
rect 1357 -323 1391 -307
rect 1357 -341 1391 -323
rect 1357 -391 1391 -379
rect 1357 -413 1391 -391
rect 1357 -459 1391 -451
rect 1357 -485 1391 -459
rect 1357 -527 1391 -523
rect 1357 -557 1391 -527
rect 1357 -629 1391 -595
rect 1357 -697 1391 -667
rect 1357 -701 1391 -697
rect 1357 -765 1391 -739
rect 1357 -773 1391 -765
rect 1357 -833 1391 -811
rect 1357 -845 1391 -833
rect 1357 -901 1391 -883
rect 1357 -917 1391 -901
rect 1357 -969 1391 -955
rect 1357 -989 1391 -969
rect 1357 -1037 1391 -1027
rect 1357 -1061 1391 -1037
rect 1357 -1105 1391 -1099
rect 1357 -1133 1391 -1105
rect 1357 -1173 1391 -1171
rect 1357 -1205 1391 -1173
rect 1357 -1275 1391 -1243
rect 1357 -1277 1391 -1275
rect 1815 1275 1849 1277
rect 1815 1243 1849 1275
rect 1815 1173 1849 1205
rect 1815 1171 1849 1173
rect 1815 1105 1849 1133
rect 1815 1099 1849 1105
rect 1815 1037 1849 1061
rect 1815 1027 1849 1037
rect 1815 969 1849 989
rect 1815 955 1849 969
rect 1815 901 1849 917
rect 1815 883 1849 901
rect 1815 833 1849 845
rect 1815 811 1849 833
rect 1815 765 1849 773
rect 1815 739 1849 765
rect 1815 697 1849 701
rect 1815 667 1849 697
rect 1815 595 1849 629
rect 1815 527 1849 557
rect 1815 523 1849 527
rect 1815 459 1849 485
rect 1815 451 1849 459
rect 1815 391 1849 413
rect 1815 379 1849 391
rect 1815 323 1849 341
rect 1815 307 1849 323
rect 1815 255 1849 269
rect 1815 235 1849 255
rect 1815 187 1849 197
rect 1815 163 1849 187
rect 1815 119 1849 125
rect 1815 91 1849 119
rect 1815 51 1849 53
rect 1815 19 1849 51
rect 1815 -51 1849 -19
rect 1815 -53 1849 -51
rect 1815 -119 1849 -91
rect 1815 -125 1849 -119
rect 1815 -187 1849 -163
rect 1815 -197 1849 -187
rect 1815 -255 1849 -235
rect 1815 -269 1849 -255
rect 1815 -323 1849 -307
rect 1815 -341 1849 -323
rect 1815 -391 1849 -379
rect 1815 -413 1849 -391
rect 1815 -459 1849 -451
rect 1815 -485 1849 -459
rect 1815 -527 1849 -523
rect 1815 -557 1849 -527
rect 1815 -629 1849 -595
rect 1815 -697 1849 -667
rect 1815 -701 1849 -697
rect 1815 -765 1849 -739
rect 1815 -773 1849 -765
rect 1815 -833 1849 -811
rect 1815 -845 1849 -833
rect 1815 -901 1849 -883
rect 1815 -917 1849 -901
rect 1815 -969 1849 -955
rect 1815 -989 1849 -969
rect 1815 -1037 1849 -1027
rect 1815 -1061 1849 -1037
rect 1815 -1105 1849 -1099
rect 1815 -1133 1849 -1105
rect 1815 -1173 1849 -1171
rect 1815 -1205 1849 -1173
rect 1815 -1275 1849 -1243
rect 1815 -1277 1849 -1275
rect 2273 1275 2307 1277
rect 2273 1243 2307 1275
rect 2273 1173 2307 1205
rect 2273 1171 2307 1173
rect 2273 1105 2307 1133
rect 2273 1099 2307 1105
rect 2273 1037 2307 1061
rect 2273 1027 2307 1037
rect 2273 969 2307 989
rect 2273 955 2307 969
rect 2273 901 2307 917
rect 2273 883 2307 901
rect 2273 833 2307 845
rect 2273 811 2307 833
rect 2273 765 2307 773
rect 2273 739 2307 765
rect 2273 697 2307 701
rect 2273 667 2307 697
rect 2273 595 2307 629
rect 2273 527 2307 557
rect 2273 523 2307 527
rect 2273 459 2307 485
rect 2273 451 2307 459
rect 2273 391 2307 413
rect 2273 379 2307 391
rect 2273 323 2307 341
rect 2273 307 2307 323
rect 2273 255 2307 269
rect 2273 235 2307 255
rect 2273 187 2307 197
rect 2273 163 2307 187
rect 2273 119 2307 125
rect 2273 91 2307 119
rect 2273 51 2307 53
rect 2273 19 2307 51
rect 2273 -51 2307 -19
rect 2273 -53 2307 -51
rect 2273 -119 2307 -91
rect 2273 -125 2307 -119
rect 2273 -187 2307 -163
rect 2273 -197 2307 -187
rect 2273 -255 2307 -235
rect 2273 -269 2307 -255
rect 2273 -323 2307 -307
rect 2273 -341 2307 -323
rect 2273 -391 2307 -379
rect 2273 -413 2307 -391
rect 2273 -459 2307 -451
rect 2273 -485 2307 -459
rect 2273 -527 2307 -523
rect 2273 -557 2307 -527
rect 2273 -629 2307 -595
rect 2273 -697 2307 -667
rect 2273 -701 2307 -697
rect 2273 -765 2307 -739
rect 2273 -773 2307 -765
rect 2273 -833 2307 -811
rect 2273 -845 2307 -833
rect 2273 -901 2307 -883
rect 2273 -917 2307 -901
rect 2273 -969 2307 -955
rect 2273 -989 2307 -969
rect 2273 -1037 2307 -1027
rect 2273 -1061 2307 -1037
rect 2273 -1105 2307 -1099
rect 2273 -1133 2307 -1105
rect 2273 -1173 2307 -1171
rect 2273 -1205 2307 -1173
rect 2273 -1275 2307 -1243
rect 2273 -1277 2307 -1275
rect -2357 -1494 -2323 -1460
rect -2285 -1494 -2261 -1460
rect -2261 -1494 -2251 -1460
rect -2213 -1494 -2193 -1460
rect -2193 -1494 -2179 -1460
rect -2141 -1494 -2125 -1460
rect -2125 -1494 -2107 -1460
rect -2069 -1494 -2057 -1460
rect -2057 -1494 -2035 -1460
rect -1997 -1494 -1989 -1460
rect -1989 -1494 -1963 -1460
rect -1925 -1494 -1921 -1460
rect -1921 -1494 -1891 -1460
rect -1853 -1494 -1819 -1460
rect -1781 -1494 -1751 -1460
rect -1751 -1494 -1747 -1460
rect -1709 -1494 -1683 -1460
rect -1683 -1494 -1675 -1460
rect -1637 -1494 -1615 -1460
rect -1615 -1494 -1603 -1460
rect -1565 -1494 -1547 -1460
rect -1547 -1494 -1531 -1460
rect -1493 -1494 -1479 -1460
rect -1479 -1494 -1459 -1460
rect -1421 -1494 -1411 -1460
rect -1411 -1494 -1387 -1460
rect -1349 -1494 -1343 -1460
rect -1343 -1494 -1315 -1460
rect -1277 -1494 -1275 -1460
rect -1275 -1494 -1243 -1460
rect -1205 -1494 -1173 -1460
rect -1173 -1494 -1171 -1460
rect -1133 -1494 -1105 -1460
rect -1105 -1494 -1099 -1460
rect -1061 -1494 -1037 -1460
rect -1037 -1494 -1027 -1460
rect -989 -1494 -969 -1460
rect -969 -1494 -955 -1460
rect -917 -1494 -901 -1460
rect -901 -1494 -883 -1460
rect -845 -1494 -833 -1460
rect -833 -1494 -811 -1460
rect -773 -1494 -765 -1460
rect -765 -1494 -739 -1460
rect -701 -1494 -697 -1460
rect -697 -1494 -667 -1460
rect -629 -1494 -595 -1460
rect -557 -1494 -527 -1460
rect -527 -1494 -523 -1460
rect -485 -1494 -459 -1460
rect -459 -1494 -451 -1460
rect -413 -1494 -391 -1460
rect -391 -1494 -379 -1460
rect -341 -1494 -323 -1460
rect -323 -1494 -307 -1460
rect -269 -1494 -255 -1460
rect -255 -1494 -235 -1460
rect -197 -1494 -187 -1460
rect -187 -1494 -163 -1460
rect -125 -1494 -119 -1460
rect -119 -1494 -91 -1460
rect -53 -1494 -51 -1460
rect -51 -1494 -19 -1460
rect 19 -1494 51 -1460
rect 51 -1494 53 -1460
rect 91 -1494 119 -1460
rect 119 -1494 125 -1460
rect 163 -1494 187 -1460
rect 187 -1494 197 -1460
rect 235 -1494 255 -1460
rect 255 -1494 269 -1460
rect 307 -1494 323 -1460
rect 323 -1494 341 -1460
rect 379 -1494 391 -1460
rect 391 -1494 413 -1460
rect 451 -1494 459 -1460
rect 459 -1494 485 -1460
rect 523 -1494 527 -1460
rect 527 -1494 557 -1460
rect 595 -1494 629 -1460
rect 667 -1494 697 -1460
rect 697 -1494 701 -1460
rect 739 -1494 765 -1460
rect 765 -1494 773 -1460
rect 811 -1494 833 -1460
rect 833 -1494 845 -1460
rect 883 -1494 901 -1460
rect 901 -1494 917 -1460
rect 955 -1494 969 -1460
rect 969 -1494 989 -1460
rect 1027 -1494 1037 -1460
rect 1037 -1494 1061 -1460
rect 1099 -1494 1105 -1460
rect 1105 -1494 1133 -1460
rect 1171 -1494 1173 -1460
rect 1173 -1494 1205 -1460
rect 1243 -1494 1275 -1460
rect 1275 -1494 1277 -1460
rect 1315 -1494 1343 -1460
rect 1343 -1494 1349 -1460
rect 1387 -1494 1411 -1460
rect 1411 -1494 1421 -1460
rect 1459 -1494 1479 -1460
rect 1479 -1494 1493 -1460
rect 1531 -1494 1547 -1460
rect 1547 -1494 1565 -1460
rect 1603 -1494 1615 -1460
rect 1615 -1494 1637 -1460
rect 1675 -1494 1683 -1460
rect 1683 -1494 1709 -1460
rect 1747 -1494 1751 -1460
rect 1751 -1494 1781 -1460
rect 1819 -1494 1853 -1460
rect 1891 -1494 1921 -1460
rect 1921 -1494 1925 -1460
rect 1963 -1494 1989 -1460
rect 1989 -1494 1997 -1460
rect 2035 -1494 2057 -1460
rect 2057 -1494 2069 -1460
rect 2107 -1494 2125 -1460
rect 2125 -1494 2141 -1460
rect 2179 -1494 2193 -1460
rect 2193 -1494 2213 -1460
rect 2251 -1494 2261 -1460
rect 2261 -1494 2285 -1460
rect 2323 -1494 2357 -1460
<< metal1 >>
rect -2313 1277 -2267 1320
rect -2313 1243 -2307 1277
rect -2273 1243 -2267 1277
rect -2313 1205 -2267 1243
rect -2313 1171 -2307 1205
rect -2273 1171 -2267 1205
rect -2313 1133 -2267 1171
rect -2313 1099 -2307 1133
rect -2273 1099 -2267 1133
rect -2313 1061 -2267 1099
rect -2313 1027 -2307 1061
rect -2273 1027 -2267 1061
rect -2313 989 -2267 1027
rect -2313 955 -2307 989
rect -2273 955 -2267 989
rect -2313 917 -2267 955
rect -2313 883 -2307 917
rect -2273 883 -2267 917
rect -2313 845 -2267 883
rect -2313 811 -2307 845
rect -2273 811 -2267 845
rect -2313 773 -2267 811
rect -2313 739 -2307 773
rect -2273 739 -2267 773
rect -2313 701 -2267 739
rect -2313 667 -2307 701
rect -2273 667 -2267 701
rect -2313 629 -2267 667
rect -2313 595 -2307 629
rect -2273 595 -2267 629
rect -2313 557 -2267 595
rect -2313 523 -2307 557
rect -2273 523 -2267 557
rect -2313 485 -2267 523
rect -2313 451 -2307 485
rect -2273 451 -2267 485
rect -2313 413 -2267 451
rect -2313 379 -2307 413
rect -2273 379 -2267 413
rect -2313 341 -2267 379
rect -2313 307 -2307 341
rect -2273 307 -2267 341
rect -2313 269 -2267 307
rect -2313 235 -2307 269
rect -2273 235 -2267 269
rect -2313 197 -2267 235
rect -2313 163 -2307 197
rect -2273 163 -2267 197
rect -2313 125 -2267 163
rect -2313 91 -2307 125
rect -2273 91 -2267 125
rect -2313 53 -2267 91
rect -2313 19 -2307 53
rect -2273 19 -2267 53
rect -2313 -19 -2267 19
rect -2313 -53 -2307 -19
rect -2273 -53 -2267 -19
rect -2313 -91 -2267 -53
rect -2313 -125 -2307 -91
rect -2273 -125 -2267 -91
rect -2313 -163 -2267 -125
rect -2313 -197 -2307 -163
rect -2273 -197 -2267 -163
rect -2313 -235 -2267 -197
rect -2313 -269 -2307 -235
rect -2273 -269 -2267 -235
rect -2313 -307 -2267 -269
rect -2313 -341 -2307 -307
rect -2273 -341 -2267 -307
rect -2313 -379 -2267 -341
rect -2313 -413 -2307 -379
rect -2273 -413 -2267 -379
rect -2313 -451 -2267 -413
rect -2313 -485 -2307 -451
rect -2273 -485 -2267 -451
rect -2313 -523 -2267 -485
rect -2313 -557 -2307 -523
rect -2273 -557 -2267 -523
rect -2313 -595 -2267 -557
rect -2313 -629 -2307 -595
rect -2273 -629 -2267 -595
rect -2313 -667 -2267 -629
rect -2313 -701 -2307 -667
rect -2273 -701 -2267 -667
rect -2313 -739 -2267 -701
rect -2313 -773 -2307 -739
rect -2273 -773 -2267 -739
rect -2313 -811 -2267 -773
rect -2313 -845 -2307 -811
rect -2273 -845 -2267 -811
rect -2313 -883 -2267 -845
rect -2313 -917 -2307 -883
rect -2273 -917 -2267 -883
rect -2313 -955 -2267 -917
rect -2313 -989 -2307 -955
rect -2273 -989 -2267 -955
rect -2313 -1027 -2267 -989
rect -2313 -1061 -2307 -1027
rect -2273 -1061 -2267 -1027
rect -2313 -1099 -2267 -1061
rect -2313 -1133 -2307 -1099
rect -2273 -1133 -2267 -1099
rect -2313 -1171 -2267 -1133
rect -2313 -1205 -2307 -1171
rect -2273 -1205 -2267 -1171
rect -2313 -1243 -2267 -1205
rect -2313 -1277 -2307 -1243
rect -2273 -1277 -2267 -1243
rect -2313 -1320 -2267 -1277
rect -1855 1277 -1809 1320
rect -1855 1243 -1849 1277
rect -1815 1243 -1809 1277
rect -1855 1205 -1809 1243
rect -1855 1171 -1849 1205
rect -1815 1171 -1809 1205
rect -1855 1133 -1809 1171
rect -1855 1099 -1849 1133
rect -1815 1099 -1809 1133
rect -1855 1061 -1809 1099
rect -1855 1027 -1849 1061
rect -1815 1027 -1809 1061
rect -1855 989 -1809 1027
rect -1855 955 -1849 989
rect -1815 955 -1809 989
rect -1855 917 -1809 955
rect -1855 883 -1849 917
rect -1815 883 -1809 917
rect -1855 845 -1809 883
rect -1855 811 -1849 845
rect -1815 811 -1809 845
rect -1855 773 -1809 811
rect -1855 739 -1849 773
rect -1815 739 -1809 773
rect -1855 701 -1809 739
rect -1855 667 -1849 701
rect -1815 667 -1809 701
rect -1855 629 -1809 667
rect -1855 595 -1849 629
rect -1815 595 -1809 629
rect -1855 557 -1809 595
rect -1855 523 -1849 557
rect -1815 523 -1809 557
rect -1855 485 -1809 523
rect -1855 451 -1849 485
rect -1815 451 -1809 485
rect -1855 413 -1809 451
rect -1855 379 -1849 413
rect -1815 379 -1809 413
rect -1855 341 -1809 379
rect -1855 307 -1849 341
rect -1815 307 -1809 341
rect -1855 269 -1809 307
rect -1855 235 -1849 269
rect -1815 235 -1809 269
rect -1855 197 -1809 235
rect -1855 163 -1849 197
rect -1815 163 -1809 197
rect -1855 125 -1809 163
rect -1855 91 -1849 125
rect -1815 91 -1809 125
rect -1855 53 -1809 91
rect -1855 19 -1849 53
rect -1815 19 -1809 53
rect -1855 -19 -1809 19
rect -1855 -53 -1849 -19
rect -1815 -53 -1809 -19
rect -1855 -91 -1809 -53
rect -1855 -125 -1849 -91
rect -1815 -125 -1809 -91
rect -1855 -163 -1809 -125
rect -1855 -197 -1849 -163
rect -1815 -197 -1809 -163
rect -1855 -235 -1809 -197
rect -1855 -269 -1849 -235
rect -1815 -269 -1809 -235
rect -1855 -307 -1809 -269
rect -1855 -341 -1849 -307
rect -1815 -341 -1809 -307
rect -1855 -379 -1809 -341
rect -1855 -413 -1849 -379
rect -1815 -413 -1809 -379
rect -1855 -451 -1809 -413
rect -1855 -485 -1849 -451
rect -1815 -485 -1809 -451
rect -1855 -523 -1809 -485
rect -1855 -557 -1849 -523
rect -1815 -557 -1809 -523
rect -1855 -595 -1809 -557
rect -1855 -629 -1849 -595
rect -1815 -629 -1809 -595
rect -1855 -667 -1809 -629
rect -1855 -701 -1849 -667
rect -1815 -701 -1809 -667
rect -1855 -739 -1809 -701
rect -1855 -773 -1849 -739
rect -1815 -773 -1809 -739
rect -1855 -811 -1809 -773
rect -1855 -845 -1849 -811
rect -1815 -845 -1809 -811
rect -1855 -883 -1809 -845
rect -1855 -917 -1849 -883
rect -1815 -917 -1809 -883
rect -1855 -955 -1809 -917
rect -1855 -989 -1849 -955
rect -1815 -989 -1809 -955
rect -1855 -1027 -1809 -989
rect -1855 -1061 -1849 -1027
rect -1815 -1061 -1809 -1027
rect -1855 -1099 -1809 -1061
rect -1855 -1133 -1849 -1099
rect -1815 -1133 -1809 -1099
rect -1855 -1171 -1809 -1133
rect -1855 -1205 -1849 -1171
rect -1815 -1205 -1809 -1171
rect -1855 -1243 -1809 -1205
rect -1855 -1277 -1849 -1243
rect -1815 -1277 -1809 -1243
rect -1855 -1320 -1809 -1277
rect -1397 1277 -1351 1320
rect -1397 1243 -1391 1277
rect -1357 1243 -1351 1277
rect -1397 1205 -1351 1243
rect -1397 1171 -1391 1205
rect -1357 1171 -1351 1205
rect -1397 1133 -1351 1171
rect -1397 1099 -1391 1133
rect -1357 1099 -1351 1133
rect -1397 1061 -1351 1099
rect -1397 1027 -1391 1061
rect -1357 1027 -1351 1061
rect -1397 989 -1351 1027
rect -1397 955 -1391 989
rect -1357 955 -1351 989
rect -1397 917 -1351 955
rect -1397 883 -1391 917
rect -1357 883 -1351 917
rect -1397 845 -1351 883
rect -1397 811 -1391 845
rect -1357 811 -1351 845
rect -1397 773 -1351 811
rect -1397 739 -1391 773
rect -1357 739 -1351 773
rect -1397 701 -1351 739
rect -1397 667 -1391 701
rect -1357 667 -1351 701
rect -1397 629 -1351 667
rect -1397 595 -1391 629
rect -1357 595 -1351 629
rect -1397 557 -1351 595
rect -1397 523 -1391 557
rect -1357 523 -1351 557
rect -1397 485 -1351 523
rect -1397 451 -1391 485
rect -1357 451 -1351 485
rect -1397 413 -1351 451
rect -1397 379 -1391 413
rect -1357 379 -1351 413
rect -1397 341 -1351 379
rect -1397 307 -1391 341
rect -1357 307 -1351 341
rect -1397 269 -1351 307
rect -1397 235 -1391 269
rect -1357 235 -1351 269
rect -1397 197 -1351 235
rect -1397 163 -1391 197
rect -1357 163 -1351 197
rect -1397 125 -1351 163
rect -1397 91 -1391 125
rect -1357 91 -1351 125
rect -1397 53 -1351 91
rect -1397 19 -1391 53
rect -1357 19 -1351 53
rect -1397 -19 -1351 19
rect -1397 -53 -1391 -19
rect -1357 -53 -1351 -19
rect -1397 -91 -1351 -53
rect -1397 -125 -1391 -91
rect -1357 -125 -1351 -91
rect -1397 -163 -1351 -125
rect -1397 -197 -1391 -163
rect -1357 -197 -1351 -163
rect -1397 -235 -1351 -197
rect -1397 -269 -1391 -235
rect -1357 -269 -1351 -235
rect -1397 -307 -1351 -269
rect -1397 -341 -1391 -307
rect -1357 -341 -1351 -307
rect -1397 -379 -1351 -341
rect -1397 -413 -1391 -379
rect -1357 -413 -1351 -379
rect -1397 -451 -1351 -413
rect -1397 -485 -1391 -451
rect -1357 -485 -1351 -451
rect -1397 -523 -1351 -485
rect -1397 -557 -1391 -523
rect -1357 -557 -1351 -523
rect -1397 -595 -1351 -557
rect -1397 -629 -1391 -595
rect -1357 -629 -1351 -595
rect -1397 -667 -1351 -629
rect -1397 -701 -1391 -667
rect -1357 -701 -1351 -667
rect -1397 -739 -1351 -701
rect -1397 -773 -1391 -739
rect -1357 -773 -1351 -739
rect -1397 -811 -1351 -773
rect -1397 -845 -1391 -811
rect -1357 -845 -1351 -811
rect -1397 -883 -1351 -845
rect -1397 -917 -1391 -883
rect -1357 -917 -1351 -883
rect -1397 -955 -1351 -917
rect -1397 -989 -1391 -955
rect -1357 -989 -1351 -955
rect -1397 -1027 -1351 -989
rect -1397 -1061 -1391 -1027
rect -1357 -1061 -1351 -1027
rect -1397 -1099 -1351 -1061
rect -1397 -1133 -1391 -1099
rect -1357 -1133 -1351 -1099
rect -1397 -1171 -1351 -1133
rect -1397 -1205 -1391 -1171
rect -1357 -1205 -1351 -1171
rect -1397 -1243 -1351 -1205
rect -1397 -1277 -1391 -1243
rect -1357 -1277 -1351 -1243
rect -1397 -1320 -1351 -1277
rect -939 1277 -893 1320
rect -939 1243 -933 1277
rect -899 1243 -893 1277
rect -939 1205 -893 1243
rect -939 1171 -933 1205
rect -899 1171 -893 1205
rect -939 1133 -893 1171
rect -939 1099 -933 1133
rect -899 1099 -893 1133
rect -939 1061 -893 1099
rect -939 1027 -933 1061
rect -899 1027 -893 1061
rect -939 989 -893 1027
rect -939 955 -933 989
rect -899 955 -893 989
rect -939 917 -893 955
rect -939 883 -933 917
rect -899 883 -893 917
rect -939 845 -893 883
rect -939 811 -933 845
rect -899 811 -893 845
rect -939 773 -893 811
rect -939 739 -933 773
rect -899 739 -893 773
rect -939 701 -893 739
rect -939 667 -933 701
rect -899 667 -893 701
rect -939 629 -893 667
rect -939 595 -933 629
rect -899 595 -893 629
rect -939 557 -893 595
rect -939 523 -933 557
rect -899 523 -893 557
rect -939 485 -893 523
rect -939 451 -933 485
rect -899 451 -893 485
rect -939 413 -893 451
rect -939 379 -933 413
rect -899 379 -893 413
rect -939 341 -893 379
rect -939 307 -933 341
rect -899 307 -893 341
rect -939 269 -893 307
rect -939 235 -933 269
rect -899 235 -893 269
rect -939 197 -893 235
rect -939 163 -933 197
rect -899 163 -893 197
rect -939 125 -893 163
rect -939 91 -933 125
rect -899 91 -893 125
rect -939 53 -893 91
rect -939 19 -933 53
rect -899 19 -893 53
rect -939 -19 -893 19
rect -939 -53 -933 -19
rect -899 -53 -893 -19
rect -939 -91 -893 -53
rect -939 -125 -933 -91
rect -899 -125 -893 -91
rect -939 -163 -893 -125
rect -939 -197 -933 -163
rect -899 -197 -893 -163
rect -939 -235 -893 -197
rect -939 -269 -933 -235
rect -899 -269 -893 -235
rect -939 -307 -893 -269
rect -939 -341 -933 -307
rect -899 -341 -893 -307
rect -939 -379 -893 -341
rect -939 -413 -933 -379
rect -899 -413 -893 -379
rect -939 -451 -893 -413
rect -939 -485 -933 -451
rect -899 -485 -893 -451
rect -939 -523 -893 -485
rect -939 -557 -933 -523
rect -899 -557 -893 -523
rect -939 -595 -893 -557
rect -939 -629 -933 -595
rect -899 -629 -893 -595
rect -939 -667 -893 -629
rect -939 -701 -933 -667
rect -899 -701 -893 -667
rect -939 -739 -893 -701
rect -939 -773 -933 -739
rect -899 -773 -893 -739
rect -939 -811 -893 -773
rect -939 -845 -933 -811
rect -899 -845 -893 -811
rect -939 -883 -893 -845
rect -939 -917 -933 -883
rect -899 -917 -893 -883
rect -939 -955 -893 -917
rect -939 -989 -933 -955
rect -899 -989 -893 -955
rect -939 -1027 -893 -989
rect -939 -1061 -933 -1027
rect -899 -1061 -893 -1027
rect -939 -1099 -893 -1061
rect -939 -1133 -933 -1099
rect -899 -1133 -893 -1099
rect -939 -1171 -893 -1133
rect -939 -1205 -933 -1171
rect -899 -1205 -893 -1171
rect -939 -1243 -893 -1205
rect -939 -1277 -933 -1243
rect -899 -1277 -893 -1243
rect -939 -1320 -893 -1277
rect -481 1277 -435 1320
rect -481 1243 -475 1277
rect -441 1243 -435 1277
rect -481 1205 -435 1243
rect -481 1171 -475 1205
rect -441 1171 -435 1205
rect -481 1133 -435 1171
rect -481 1099 -475 1133
rect -441 1099 -435 1133
rect -481 1061 -435 1099
rect -481 1027 -475 1061
rect -441 1027 -435 1061
rect -481 989 -435 1027
rect -481 955 -475 989
rect -441 955 -435 989
rect -481 917 -435 955
rect -481 883 -475 917
rect -441 883 -435 917
rect -481 845 -435 883
rect -481 811 -475 845
rect -441 811 -435 845
rect -481 773 -435 811
rect -481 739 -475 773
rect -441 739 -435 773
rect -481 701 -435 739
rect -481 667 -475 701
rect -441 667 -435 701
rect -481 629 -435 667
rect -481 595 -475 629
rect -441 595 -435 629
rect -481 557 -435 595
rect -481 523 -475 557
rect -441 523 -435 557
rect -481 485 -435 523
rect -481 451 -475 485
rect -441 451 -435 485
rect -481 413 -435 451
rect -481 379 -475 413
rect -441 379 -435 413
rect -481 341 -435 379
rect -481 307 -475 341
rect -441 307 -435 341
rect -481 269 -435 307
rect -481 235 -475 269
rect -441 235 -435 269
rect -481 197 -435 235
rect -481 163 -475 197
rect -441 163 -435 197
rect -481 125 -435 163
rect -481 91 -475 125
rect -441 91 -435 125
rect -481 53 -435 91
rect -481 19 -475 53
rect -441 19 -435 53
rect -481 -19 -435 19
rect -481 -53 -475 -19
rect -441 -53 -435 -19
rect -481 -91 -435 -53
rect -481 -125 -475 -91
rect -441 -125 -435 -91
rect -481 -163 -435 -125
rect -481 -197 -475 -163
rect -441 -197 -435 -163
rect -481 -235 -435 -197
rect -481 -269 -475 -235
rect -441 -269 -435 -235
rect -481 -307 -435 -269
rect -481 -341 -475 -307
rect -441 -341 -435 -307
rect -481 -379 -435 -341
rect -481 -413 -475 -379
rect -441 -413 -435 -379
rect -481 -451 -435 -413
rect -481 -485 -475 -451
rect -441 -485 -435 -451
rect -481 -523 -435 -485
rect -481 -557 -475 -523
rect -441 -557 -435 -523
rect -481 -595 -435 -557
rect -481 -629 -475 -595
rect -441 -629 -435 -595
rect -481 -667 -435 -629
rect -481 -701 -475 -667
rect -441 -701 -435 -667
rect -481 -739 -435 -701
rect -481 -773 -475 -739
rect -441 -773 -435 -739
rect -481 -811 -435 -773
rect -481 -845 -475 -811
rect -441 -845 -435 -811
rect -481 -883 -435 -845
rect -481 -917 -475 -883
rect -441 -917 -435 -883
rect -481 -955 -435 -917
rect -481 -989 -475 -955
rect -441 -989 -435 -955
rect -481 -1027 -435 -989
rect -481 -1061 -475 -1027
rect -441 -1061 -435 -1027
rect -481 -1099 -435 -1061
rect -481 -1133 -475 -1099
rect -441 -1133 -435 -1099
rect -481 -1171 -435 -1133
rect -481 -1205 -475 -1171
rect -441 -1205 -435 -1171
rect -481 -1243 -435 -1205
rect -481 -1277 -475 -1243
rect -441 -1277 -435 -1243
rect -481 -1320 -435 -1277
rect -23 1277 23 1320
rect -23 1243 -17 1277
rect 17 1243 23 1277
rect -23 1205 23 1243
rect -23 1171 -17 1205
rect 17 1171 23 1205
rect -23 1133 23 1171
rect -23 1099 -17 1133
rect 17 1099 23 1133
rect -23 1061 23 1099
rect -23 1027 -17 1061
rect 17 1027 23 1061
rect -23 989 23 1027
rect -23 955 -17 989
rect 17 955 23 989
rect -23 917 23 955
rect -23 883 -17 917
rect 17 883 23 917
rect -23 845 23 883
rect -23 811 -17 845
rect 17 811 23 845
rect -23 773 23 811
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -811 23 -773
rect -23 -845 -17 -811
rect 17 -845 23 -811
rect -23 -883 23 -845
rect -23 -917 -17 -883
rect 17 -917 23 -883
rect -23 -955 23 -917
rect -23 -989 -17 -955
rect 17 -989 23 -955
rect -23 -1027 23 -989
rect -23 -1061 -17 -1027
rect 17 -1061 23 -1027
rect -23 -1099 23 -1061
rect -23 -1133 -17 -1099
rect 17 -1133 23 -1099
rect -23 -1171 23 -1133
rect -23 -1205 -17 -1171
rect 17 -1205 23 -1171
rect -23 -1243 23 -1205
rect -23 -1277 -17 -1243
rect 17 -1277 23 -1243
rect -23 -1320 23 -1277
rect 435 1277 481 1320
rect 435 1243 441 1277
rect 475 1243 481 1277
rect 435 1205 481 1243
rect 435 1171 441 1205
rect 475 1171 481 1205
rect 435 1133 481 1171
rect 435 1099 441 1133
rect 475 1099 481 1133
rect 435 1061 481 1099
rect 435 1027 441 1061
rect 475 1027 481 1061
rect 435 989 481 1027
rect 435 955 441 989
rect 475 955 481 989
rect 435 917 481 955
rect 435 883 441 917
rect 475 883 481 917
rect 435 845 481 883
rect 435 811 441 845
rect 475 811 481 845
rect 435 773 481 811
rect 435 739 441 773
rect 475 739 481 773
rect 435 701 481 739
rect 435 667 441 701
rect 475 667 481 701
rect 435 629 481 667
rect 435 595 441 629
rect 475 595 481 629
rect 435 557 481 595
rect 435 523 441 557
rect 475 523 481 557
rect 435 485 481 523
rect 435 451 441 485
rect 475 451 481 485
rect 435 413 481 451
rect 435 379 441 413
rect 475 379 481 413
rect 435 341 481 379
rect 435 307 441 341
rect 475 307 481 341
rect 435 269 481 307
rect 435 235 441 269
rect 475 235 481 269
rect 435 197 481 235
rect 435 163 441 197
rect 475 163 481 197
rect 435 125 481 163
rect 435 91 441 125
rect 475 91 481 125
rect 435 53 481 91
rect 435 19 441 53
rect 475 19 481 53
rect 435 -19 481 19
rect 435 -53 441 -19
rect 475 -53 481 -19
rect 435 -91 481 -53
rect 435 -125 441 -91
rect 475 -125 481 -91
rect 435 -163 481 -125
rect 435 -197 441 -163
rect 475 -197 481 -163
rect 435 -235 481 -197
rect 435 -269 441 -235
rect 475 -269 481 -235
rect 435 -307 481 -269
rect 435 -341 441 -307
rect 475 -341 481 -307
rect 435 -379 481 -341
rect 435 -413 441 -379
rect 475 -413 481 -379
rect 435 -451 481 -413
rect 435 -485 441 -451
rect 475 -485 481 -451
rect 435 -523 481 -485
rect 435 -557 441 -523
rect 475 -557 481 -523
rect 435 -595 481 -557
rect 435 -629 441 -595
rect 475 -629 481 -595
rect 435 -667 481 -629
rect 435 -701 441 -667
rect 475 -701 481 -667
rect 435 -739 481 -701
rect 435 -773 441 -739
rect 475 -773 481 -739
rect 435 -811 481 -773
rect 435 -845 441 -811
rect 475 -845 481 -811
rect 435 -883 481 -845
rect 435 -917 441 -883
rect 475 -917 481 -883
rect 435 -955 481 -917
rect 435 -989 441 -955
rect 475 -989 481 -955
rect 435 -1027 481 -989
rect 435 -1061 441 -1027
rect 475 -1061 481 -1027
rect 435 -1099 481 -1061
rect 435 -1133 441 -1099
rect 475 -1133 481 -1099
rect 435 -1171 481 -1133
rect 435 -1205 441 -1171
rect 475 -1205 481 -1171
rect 435 -1243 481 -1205
rect 435 -1277 441 -1243
rect 475 -1277 481 -1243
rect 435 -1320 481 -1277
rect 893 1277 939 1320
rect 893 1243 899 1277
rect 933 1243 939 1277
rect 893 1205 939 1243
rect 893 1171 899 1205
rect 933 1171 939 1205
rect 893 1133 939 1171
rect 893 1099 899 1133
rect 933 1099 939 1133
rect 893 1061 939 1099
rect 893 1027 899 1061
rect 933 1027 939 1061
rect 893 989 939 1027
rect 893 955 899 989
rect 933 955 939 989
rect 893 917 939 955
rect 893 883 899 917
rect 933 883 939 917
rect 893 845 939 883
rect 893 811 899 845
rect 933 811 939 845
rect 893 773 939 811
rect 893 739 899 773
rect 933 739 939 773
rect 893 701 939 739
rect 893 667 899 701
rect 933 667 939 701
rect 893 629 939 667
rect 893 595 899 629
rect 933 595 939 629
rect 893 557 939 595
rect 893 523 899 557
rect 933 523 939 557
rect 893 485 939 523
rect 893 451 899 485
rect 933 451 939 485
rect 893 413 939 451
rect 893 379 899 413
rect 933 379 939 413
rect 893 341 939 379
rect 893 307 899 341
rect 933 307 939 341
rect 893 269 939 307
rect 893 235 899 269
rect 933 235 939 269
rect 893 197 939 235
rect 893 163 899 197
rect 933 163 939 197
rect 893 125 939 163
rect 893 91 899 125
rect 933 91 939 125
rect 893 53 939 91
rect 893 19 899 53
rect 933 19 939 53
rect 893 -19 939 19
rect 893 -53 899 -19
rect 933 -53 939 -19
rect 893 -91 939 -53
rect 893 -125 899 -91
rect 933 -125 939 -91
rect 893 -163 939 -125
rect 893 -197 899 -163
rect 933 -197 939 -163
rect 893 -235 939 -197
rect 893 -269 899 -235
rect 933 -269 939 -235
rect 893 -307 939 -269
rect 893 -341 899 -307
rect 933 -341 939 -307
rect 893 -379 939 -341
rect 893 -413 899 -379
rect 933 -413 939 -379
rect 893 -451 939 -413
rect 893 -485 899 -451
rect 933 -485 939 -451
rect 893 -523 939 -485
rect 893 -557 899 -523
rect 933 -557 939 -523
rect 893 -595 939 -557
rect 893 -629 899 -595
rect 933 -629 939 -595
rect 893 -667 939 -629
rect 893 -701 899 -667
rect 933 -701 939 -667
rect 893 -739 939 -701
rect 893 -773 899 -739
rect 933 -773 939 -739
rect 893 -811 939 -773
rect 893 -845 899 -811
rect 933 -845 939 -811
rect 893 -883 939 -845
rect 893 -917 899 -883
rect 933 -917 939 -883
rect 893 -955 939 -917
rect 893 -989 899 -955
rect 933 -989 939 -955
rect 893 -1027 939 -989
rect 893 -1061 899 -1027
rect 933 -1061 939 -1027
rect 893 -1099 939 -1061
rect 893 -1133 899 -1099
rect 933 -1133 939 -1099
rect 893 -1171 939 -1133
rect 893 -1205 899 -1171
rect 933 -1205 939 -1171
rect 893 -1243 939 -1205
rect 893 -1277 899 -1243
rect 933 -1277 939 -1243
rect 893 -1320 939 -1277
rect 1351 1277 1397 1320
rect 1351 1243 1357 1277
rect 1391 1243 1397 1277
rect 1351 1205 1397 1243
rect 1351 1171 1357 1205
rect 1391 1171 1397 1205
rect 1351 1133 1397 1171
rect 1351 1099 1357 1133
rect 1391 1099 1397 1133
rect 1351 1061 1397 1099
rect 1351 1027 1357 1061
rect 1391 1027 1397 1061
rect 1351 989 1397 1027
rect 1351 955 1357 989
rect 1391 955 1397 989
rect 1351 917 1397 955
rect 1351 883 1357 917
rect 1391 883 1397 917
rect 1351 845 1397 883
rect 1351 811 1357 845
rect 1391 811 1397 845
rect 1351 773 1397 811
rect 1351 739 1357 773
rect 1391 739 1397 773
rect 1351 701 1397 739
rect 1351 667 1357 701
rect 1391 667 1397 701
rect 1351 629 1397 667
rect 1351 595 1357 629
rect 1391 595 1397 629
rect 1351 557 1397 595
rect 1351 523 1357 557
rect 1391 523 1397 557
rect 1351 485 1397 523
rect 1351 451 1357 485
rect 1391 451 1397 485
rect 1351 413 1397 451
rect 1351 379 1357 413
rect 1391 379 1397 413
rect 1351 341 1397 379
rect 1351 307 1357 341
rect 1391 307 1397 341
rect 1351 269 1397 307
rect 1351 235 1357 269
rect 1391 235 1397 269
rect 1351 197 1397 235
rect 1351 163 1357 197
rect 1391 163 1397 197
rect 1351 125 1397 163
rect 1351 91 1357 125
rect 1391 91 1397 125
rect 1351 53 1397 91
rect 1351 19 1357 53
rect 1391 19 1397 53
rect 1351 -19 1397 19
rect 1351 -53 1357 -19
rect 1391 -53 1397 -19
rect 1351 -91 1397 -53
rect 1351 -125 1357 -91
rect 1391 -125 1397 -91
rect 1351 -163 1397 -125
rect 1351 -197 1357 -163
rect 1391 -197 1397 -163
rect 1351 -235 1397 -197
rect 1351 -269 1357 -235
rect 1391 -269 1397 -235
rect 1351 -307 1397 -269
rect 1351 -341 1357 -307
rect 1391 -341 1397 -307
rect 1351 -379 1397 -341
rect 1351 -413 1357 -379
rect 1391 -413 1397 -379
rect 1351 -451 1397 -413
rect 1351 -485 1357 -451
rect 1391 -485 1397 -451
rect 1351 -523 1397 -485
rect 1351 -557 1357 -523
rect 1391 -557 1397 -523
rect 1351 -595 1397 -557
rect 1351 -629 1357 -595
rect 1391 -629 1397 -595
rect 1351 -667 1397 -629
rect 1351 -701 1357 -667
rect 1391 -701 1397 -667
rect 1351 -739 1397 -701
rect 1351 -773 1357 -739
rect 1391 -773 1397 -739
rect 1351 -811 1397 -773
rect 1351 -845 1357 -811
rect 1391 -845 1397 -811
rect 1351 -883 1397 -845
rect 1351 -917 1357 -883
rect 1391 -917 1397 -883
rect 1351 -955 1397 -917
rect 1351 -989 1357 -955
rect 1391 -989 1397 -955
rect 1351 -1027 1397 -989
rect 1351 -1061 1357 -1027
rect 1391 -1061 1397 -1027
rect 1351 -1099 1397 -1061
rect 1351 -1133 1357 -1099
rect 1391 -1133 1397 -1099
rect 1351 -1171 1397 -1133
rect 1351 -1205 1357 -1171
rect 1391 -1205 1397 -1171
rect 1351 -1243 1397 -1205
rect 1351 -1277 1357 -1243
rect 1391 -1277 1397 -1243
rect 1351 -1320 1397 -1277
rect 1809 1277 1855 1320
rect 1809 1243 1815 1277
rect 1849 1243 1855 1277
rect 1809 1205 1855 1243
rect 1809 1171 1815 1205
rect 1849 1171 1855 1205
rect 1809 1133 1855 1171
rect 1809 1099 1815 1133
rect 1849 1099 1855 1133
rect 1809 1061 1855 1099
rect 1809 1027 1815 1061
rect 1849 1027 1855 1061
rect 1809 989 1855 1027
rect 1809 955 1815 989
rect 1849 955 1855 989
rect 1809 917 1855 955
rect 1809 883 1815 917
rect 1849 883 1855 917
rect 1809 845 1855 883
rect 1809 811 1815 845
rect 1849 811 1855 845
rect 1809 773 1855 811
rect 1809 739 1815 773
rect 1849 739 1855 773
rect 1809 701 1855 739
rect 1809 667 1815 701
rect 1849 667 1855 701
rect 1809 629 1855 667
rect 1809 595 1815 629
rect 1849 595 1855 629
rect 1809 557 1855 595
rect 1809 523 1815 557
rect 1849 523 1855 557
rect 1809 485 1855 523
rect 1809 451 1815 485
rect 1849 451 1855 485
rect 1809 413 1855 451
rect 1809 379 1815 413
rect 1849 379 1855 413
rect 1809 341 1855 379
rect 1809 307 1815 341
rect 1849 307 1855 341
rect 1809 269 1855 307
rect 1809 235 1815 269
rect 1849 235 1855 269
rect 1809 197 1855 235
rect 1809 163 1815 197
rect 1849 163 1855 197
rect 1809 125 1855 163
rect 1809 91 1815 125
rect 1849 91 1855 125
rect 1809 53 1855 91
rect 1809 19 1815 53
rect 1849 19 1855 53
rect 1809 -19 1855 19
rect 1809 -53 1815 -19
rect 1849 -53 1855 -19
rect 1809 -91 1855 -53
rect 1809 -125 1815 -91
rect 1849 -125 1855 -91
rect 1809 -163 1855 -125
rect 1809 -197 1815 -163
rect 1849 -197 1855 -163
rect 1809 -235 1855 -197
rect 1809 -269 1815 -235
rect 1849 -269 1855 -235
rect 1809 -307 1855 -269
rect 1809 -341 1815 -307
rect 1849 -341 1855 -307
rect 1809 -379 1855 -341
rect 1809 -413 1815 -379
rect 1849 -413 1855 -379
rect 1809 -451 1855 -413
rect 1809 -485 1815 -451
rect 1849 -485 1855 -451
rect 1809 -523 1855 -485
rect 1809 -557 1815 -523
rect 1849 -557 1855 -523
rect 1809 -595 1855 -557
rect 1809 -629 1815 -595
rect 1849 -629 1855 -595
rect 1809 -667 1855 -629
rect 1809 -701 1815 -667
rect 1849 -701 1855 -667
rect 1809 -739 1855 -701
rect 1809 -773 1815 -739
rect 1849 -773 1855 -739
rect 1809 -811 1855 -773
rect 1809 -845 1815 -811
rect 1849 -845 1855 -811
rect 1809 -883 1855 -845
rect 1809 -917 1815 -883
rect 1849 -917 1855 -883
rect 1809 -955 1855 -917
rect 1809 -989 1815 -955
rect 1849 -989 1855 -955
rect 1809 -1027 1855 -989
rect 1809 -1061 1815 -1027
rect 1849 -1061 1855 -1027
rect 1809 -1099 1855 -1061
rect 1809 -1133 1815 -1099
rect 1849 -1133 1855 -1099
rect 1809 -1171 1855 -1133
rect 1809 -1205 1815 -1171
rect 1849 -1205 1855 -1171
rect 1809 -1243 1855 -1205
rect 1809 -1277 1815 -1243
rect 1849 -1277 1855 -1243
rect 1809 -1320 1855 -1277
rect 2267 1277 2313 1320
rect 2267 1243 2273 1277
rect 2307 1243 2313 1277
rect 2267 1205 2313 1243
rect 2267 1171 2273 1205
rect 2307 1171 2313 1205
rect 2267 1133 2313 1171
rect 2267 1099 2273 1133
rect 2307 1099 2313 1133
rect 2267 1061 2313 1099
rect 2267 1027 2273 1061
rect 2307 1027 2313 1061
rect 2267 989 2313 1027
rect 2267 955 2273 989
rect 2307 955 2313 989
rect 2267 917 2313 955
rect 2267 883 2273 917
rect 2307 883 2313 917
rect 2267 845 2313 883
rect 2267 811 2273 845
rect 2307 811 2313 845
rect 2267 773 2313 811
rect 2267 739 2273 773
rect 2307 739 2313 773
rect 2267 701 2313 739
rect 2267 667 2273 701
rect 2307 667 2313 701
rect 2267 629 2313 667
rect 2267 595 2273 629
rect 2307 595 2313 629
rect 2267 557 2313 595
rect 2267 523 2273 557
rect 2307 523 2313 557
rect 2267 485 2313 523
rect 2267 451 2273 485
rect 2307 451 2313 485
rect 2267 413 2313 451
rect 2267 379 2273 413
rect 2307 379 2313 413
rect 2267 341 2313 379
rect 2267 307 2273 341
rect 2307 307 2313 341
rect 2267 269 2313 307
rect 2267 235 2273 269
rect 2307 235 2313 269
rect 2267 197 2313 235
rect 2267 163 2273 197
rect 2307 163 2313 197
rect 2267 125 2313 163
rect 2267 91 2273 125
rect 2307 91 2313 125
rect 2267 53 2313 91
rect 2267 19 2273 53
rect 2307 19 2313 53
rect 2267 -19 2313 19
rect 2267 -53 2273 -19
rect 2307 -53 2313 -19
rect 2267 -91 2313 -53
rect 2267 -125 2273 -91
rect 2307 -125 2313 -91
rect 2267 -163 2313 -125
rect 2267 -197 2273 -163
rect 2307 -197 2313 -163
rect 2267 -235 2313 -197
rect 2267 -269 2273 -235
rect 2307 -269 2313 -235
rect 2267 -307 2313 -269
rect 2267 -341 2273 -307
rect 2307 -341 2313 -307
rect 2267 -379 2313 -341
rect 2267 -413 2273 -379
rect 2307 -413 2313 -379
rect 2267 -451 2313 -413
rect 2267 -485 2273 -451
rect 2307 -485 2313 -451
rect 2267 -523 2313 -485
rect 2267 -557 2273 -523
rect 2307 -557 2313 -523
rect 2267 -595 2313 -557
rect 2267 -629 2273 -595
rect 2307 -629 2313 -595
rect 2267 -667 2313 -629
rect 2267 -701 2273 -667
rect 2307 -701 2313 -667
rect 2267 -739 2313 -701
rect 2267 -773 2273 -739
rect 2307 -773 2313 -739
rect 2267 -811 2313 -773
rect 2267 -845 2273 -811
rect 2307 -845 2313 -811
rect 2267 -883 2313 -845
rect 2267 -917 2273 -883
rect 2307 -917 2313 -883
rect 2267 -955 2313 -917
rect 2267 -989 2273 -955
rect 2307 -989 2313 -955
rect 2267 -1027 2313 -989
rect 2267 -1061 2273 -1027
rect 2307 -1061 2313 -1027
rect 2267 -1099 2313 -1061
rect 2267 -1133 2273 -1099
rect 2307 -1133 2313 -1099
rect 2267 -1171 2313 -1133
rect 2267 -1205 2273 -1171
rect 2307 -1205 2313 -1171
rect 2267 -1243 2313 -1205
rect 2267 -1277 2273 -1243
rect 2307 -1277 2313 -1243
rect 2267 -1320 2313 -1277
rect -2399 -1460 2399 -1454
rect -2399 -1494 -2357 -1460
rect -2323 -1494 -2285 -1460
rect -2251 -1494 -2213 -1460
rect -2179 -1494 -2141 -1460
rect -2107 -1494 -2069 -1460
rect -2035 -1494 -1997 -1460
rect -1963 -1494 -1925 -1460
rect -1891 -1494 -1853 -1460
rect -1819 -1494 -1781 -1460
rect -1747 -1494 -1709 -1460
rect -1675 -1494 -1637 -1460
rect -1603 -1494 -1565 -1460
rect -1531 -1494 -1493 -1460
rect -1459 -1494 -1421 -1460
rect -1387 -1494 -1349 -1460
rect -1315 -1494 -1277 -1460
rect -1243 -1494 -1205 -1460
rect -1171 -1494 -1133 -1460
rect -1099 -1494 -1061 -1460
rect -1027 -1494 -989 -1460
rect -955 -1494 -917 -1460
rect -883 -1494 -845 -1460
rect -811 -1494 -773 -1460
rect -739 -1494 -701 -1460
rect -667 -1494 -629 -1460
rect -595 -1494 -557 -1460
rect -523 -1494 -485 -1460
rect -451 -1494 -413 -1460
rect -379 -1494 -341 -1460
rect -307 -1494 -269 -1460
rect -235 -1494 -197 -1460
rect -163 -1494 -125 -1460
rect -91 -1494 -53 -1460
rect -19 -1494 19 -1460
rect 53 -1494 91 -1460
rect 125 -1494 163 -1460
rect 197 -1494 235 -1460
rect 269 -1494 307 -1460
rect 341 -1494 379 -1460
rect 413 -1494 451 -1460
rect 485 -1494 523 -1460
rect 557 -1494 595 -1460
rect 629 -1494 667 -1460
rect 701 -1494 739 -1460
rect 773 -1494 811 -1460
rect 845 -1494 883 -1460
rect 917 -1494 955 -1460
rect 989 -1494 1027 -1460
rect 1061 -1494 1099 -1460
rect 1133 -1494 1171 -1460
rect 1205 -1494 1243 -1460
rect 1277 -1494 1315 -1460
rect 1349 -1494 1387 -1460
rect 1421 -1494 1459 -1460
rect 1493 -1494 1531 -1460
rect 1565 -1494 1603 -1460
rect 1637 -1494 1675 -1460
rect 1709 -1494 1747 -1460
rect 1781 -1494 1819 -1460
rect 1853 -1494 1891 -1460
rect 1925 -1494 1963 -1460
rect 1997 -1494 2035 -1460
rect 2069 -1494 2107 -1460
rect 2141 -1494 2179 -1460
rect 2213 -1494 2251 -1460
rect 2285 -1494 2323 -1460
rect 2357 -1494 2399 -1460
rect -2399 -1500 2399 -1494
<< properties >>
string FIXED_BBOX -2404 -1477 2404 1477
<< end >>
