magic
tech sky130A
magscale 1 2
timestamp 1608050792
<< nwell >>
rect -854 -1549 854 1549
<< pmos >>
rect -658 -1330 -258 1330
rect -200 -1330 200 1330
rect 258 -1330 658 1330
<< pdiff >>
rect -716 1318 -658 1330
rect -716 -1318 -704 1318
rect -670 -1318 -658 1318
rect -716 -1330 -658 -1318
rect -258 1318 -200 1330
rect -258 -1318 -246 1318
rect -212 -1318 -200 1318
rect -258 -1330 -200 -1318
rect 200 1318 258 1330
rect 200 -1318 212 1318
rect 246 -1318 258 1318
rect 200 -1330 258 -1318
rect 658 1318 716 1330
rect 658 -1318 670 1318
rect 704 -1318 716 1318
rect 658 -1330 716 -1318
<< pdiffc >>
rect -704 -1318 -670 1318
rect -246 -1318 -212 1318
rect 212 -1318 246 1318
rect 670 -1318 704 1318
<< nsubdiff >>
rect -818 1479 -722 1513
rect 722 1479 818 1513
rect -818 1417 -784 1479
rect 784 1417 818 1479
rect -818 -1479 -784 -1417
rect 784 -1479 818 -1417
rect -818 -1513 -722 -1479
rect 722 -1513 818 -1479
<< nsubdiffcont >>
rect -722 1479 722 1513
rect -818 -1417 -784 1417
rect 784 -1417 818 1417
rect -722 -1513 722 -1479
<< poly >>
rect -511 1411 -405 1427
rect -511 1394 -495 1411
rect -658 1377 -495 1394
rect -421 1394 -405 1411
rect -53 1411 53 1427
rect -53 1394 -37 1411
rect -421 1377 -258 1394
rect -658 1330 -258 1377
rect -200 1377 -37 1394
rect 37 1394 53 1411
rect 405 1411 511 1427
rect 405 1394 421 1411
rect 37 1377 200 1394
rect -200 1330 200 1377
rect 258 1377 421 1394
rect 495 1394 511 1411
rect 495 1377 658 1394
rect 258 1330 658 1377
rect -658 -1377 -258 -1330
rect -658 -1394 -495 -1377
rect -511 -1411 -495 -1394
rect -421 -1394 -258 -1377
rect -200 -1377 200 -1330
rect -200 -1394 -37 -1377
rect -421 -1411 -405 -1394
rect -511 -1427 -405 -1411
rect -53 -1411 -37 -1394
rect 37 -1394 200 -1377
rect 258 -1377 658 -1330
rect 258 -1394 421 -1377
rect 37 -1411 53 -1394
rect -53 -1427 53 -1411
rect 405 -1411 421 -1394
rect 495 -1394 658 -1377
rect 495 -1411 511 -1394
rect 405 -1427 511 -1411
<< polycont >>
rect -495 1377 -421 1411
rect -37 1377 37 1411
rect 421 1377 495 1411
rect -495 -1411 -421 -1377
rect -37 -1411 37 -1377
rect 421 -1411 495 -1377
<< locali >>
rect -818 1417 -784 1513
rect 784 1417 818 1513
rect -511 1377 -495 1411
rect -421 1377 -405 1411
rect -53 1377 -37 1411
rect 37 1377 53 1411
rect 405 1377 421 1411
rect 495 1377 511 1411
rect -704 1318 -670 1334
rect -704 -1334 -670 -1318
rect -246 1318 -212 1334
rect -246 -1334 -212 -1318
rect 212 1318 246 1334
rect 212 -1334 246 -1318
rect 670 1318 704 1334
rect 670 -1334 704 -1318
rect -511 -1411 -495 -1377
rect -421 -1411 -405 -1377
rect -53 -1411 -37 -1377
rect 37 -1411 53 -1377
rect 405 -1411 421 -1377
rect 495 -1411 511 -1377
rect -818 -1479 -784 -1417
rect 784 -1479 818 -1417
rect -818 -1513 -722 -1479
rect 722 -1513 818 -1479
<< viali >>
rect -784 1479 -722 1513
rect -722 1479 722 1513
rect 722 1479 784 1513
rect -704 -1318 -670 1318
rect -246 -1318 -212 1318
rect 212 -1318 246 1318
rect 670 -1318 704 1318
<< metal1 >>
rect -796 1513 796 1519
rect -796 1479 -784 1513
rect 784 1479 796 1513
rect -796 1473 796 1479
rect -710 1318 -664 1330
rect -710 -1318 -704 1318
rect -670 -1318 -664 1318
rect -710 -1330 -664 -1318
rect -252 1318 -206 1330
rect -252 -1318 -246 1318
rect -212 -1318 -206 1318
rect -252 -1330 -206 -1318
rect 206 1318 252 1330
rect 206 -1318 212 1318
rect 246 -1318 252 1318
rect 206 -1330 252 -1318
rect 664 1318 710 1330
rect 664 -1318 670 1318
rect 704 -1318 710 1318
rect 664 -1330 710 -1318
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -801 -1496 801 1496
string parameters w 13.3 l 2 m 1 nf 3 diffcov 100 polycov 20 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 100 viagb 0 viagate 0 viadrn 100 viasrc 100
string library sky130
<< end >>
