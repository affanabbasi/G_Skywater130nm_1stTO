magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -98 1838 1124 1872
rect -98 1458 -64 1838
rect 1090 1458 1124 1838
rect -98 1424 1124 1458
rect 1196 1838 2418 1872
rect 1196 1458 1230 1838
rect 2384 1458 2418 1838
rect 1196 1424 2418 1458
rect 1192 806 2414 840
rect 1192 426 1226 806
rect 2380 426 2414 806
rect 1192 392 2414 426
<< nmoslvt >>
rect 66 1598 96 1698
rect 162 1598 192 1698
rect 258 1598 288 1698
rect 354 1598 384 1698
rect 450 1598 480 1698
rect 546 1598 576 1698
rect 642 1598 672 1698
rect 738 1598 768 1698
rect 834 1598 864 1698
rect 930 1598 960 1698
rect 1360 1598 1390 1698
rect 1456 1598 1486 1698
rect 1552 1598 1582 1698
rect 1648 1598 1678 1698
rect 1744 1598 1774 1698
rect 1840 1598 1870 1698
rect 1936 1598 1966 1698
rect 2032 1598 2062 1698
rect 2128 1598 2158 1698
rect 2224 1598 2254 1698
rect 1356 566 1386 666
rect 1452 566 1482 666
rect 1548 566 1578 666
rect 1644 566 1674 666
rect 1740 566 1770 666
rect 1836 566 1866 666
rect 1932 566 1962 666
rect 2028 566 2058 666
rect 2124 566 2154 666
rect 2220 566 2250 666
<< ndiff >>
rect 4 1665 66 1698
rect 4 1631 16 1665
rect 50 1631 66 1665
rect 4 1598 66 1631
rect 96 1665 162 1698
rect 96 1631 112 1665
rect 146 1631 162 1665
rect 96 1598 162 1631
rect 192 1665 258 1698
rect 192 1631 208 1665
rect 242 1631 258 1665
rect 192 1598 258 1631
rect 288 1665 354 1698
rect 288 1631 304 1665
rect 338 1631 354 1665
rect 288 1598 354 1631
rect 384 1665 450 1698
rect 384 1631 400 1665
rect 434 1631 450 1665
rect 384 1598 450 1631
rect 480 1665 546 1698
rect 480 1631 496 1665
rect 530 1631 546 1665
rect 480 1598 546 1631
rect 576 1665 642 1698
rect 576 1631 592 1665
rect 626 1631 642 1665
rect 576 1598 642 1631
rect 672 1665 738 1698
rect 672 1631 688 1665
rect 722 1631 738 1665
rect 672 1598 738 1631
rect 768 1665 834 1698
rect 768 1631 784 1665
rect 818 1631 834 1665
rect 768 1598 834 1631
rect 864 1665 930 1698
rect 864 1631 880 1665
rect 914 1631 930 1665
rect 864 1598 930 1631
rect 960 1665 1022 1698
rect 960 1631 976 1665
rect 1010 1631 1022 1665
rect 960 1598 1022 1631
rect 1298 1665 1360 1698
rect 1298 1631 1310 1665
rect 1344 1631 1360 1665
rect 1298 1598 1360 1631
rect 1390 1665 1456 1698
rect 1390 1631 1406 1665
rect 1440 1631 1456 1665
rect 1390 1598 1456 1631
rect 1486 1665 1552 1698
rect 1486 1631 1502 1665
rect 1536 1631 1552 1665
rect 1486 1598 1552 1631
rect 1582 1665 1648 1698
rect 1582 1631 1598 1665
rect 1632 1631 1648 1665
rect 1582 1598 1648 1631
rect 1678 1665 1744 1698
rect 1678 1631 1694 1665
rect 1728 1631 1744 1665
rect 1678 1598 1744 1631
rect 1774 1665 1840 1698
rect 1774 1631 1790 1665
rect 1824 1631 1840 1665
rect 1774 1598 1840 1631
rect 1870 1665 1936 1698
rect 1870 1631 1886 1665
rect 1920 1631 1936 1665
rect 1870 1598 1936 1631
rect 1966 1665 2032 1698
rect 1966 1631 1982 1665
rect 2016 1631 2032 1665
rect 1966 1598 2032 1631
rect 2062 1665 2128 1698
rect 2062 1631 2078 1665
rect 2112 1631 2128 1665
rect 2062 1598 2128 1631
rect 2158 1665 2224 1698
rect 2158 1631 2174 1665
rect 2208 1631 2224 1665
rect 2158 1598 2224 1631
rect 2254 1665 2316 1698
rect 2254 1631 2270 1665
rect 2304 1631 2316 1665
rect 2254 1598 2316 1631
rect 1294 633 1356 666
rect 1294 599 1306 633
rect 1340 599 1356 633
rect 1294 566 1356 599
rect 1386 633 1452 666
rect 1386 599 1402 633
rect 1436 599 1452 633
rect 1386 566 1452 599
rect 1482 633 1548 666
rect 1482 599 1498 633
rect 1532 599 1548 633
rect 1482 566 1548 599
rect 1578 633 1644 666
rect 1578 599 1594 633
rect 1628 599 1644 633
rect 1578 566 1644 599
rect 1674 633 1740 666
rect 1674 599 1690 633
rect 1724 599 1740 633
rect 1674 566 1740 599
rect 1770 633 1836 666
rect 1770 599 1786 633
rect 1820 599 1836 633
rect 1770 566 1836 599
rect 1866 633 1932 666
rect 1866 599 1882 633
rect 1916 599 1932 633
rect 1866 566 1932 599
rect 1962 633 2028 666
rect 1962 599 1978 633
rect 2012 599 2028 633
rect 1962 566 2028 599
rect 2058 633 2124 666
rect 2058 599 2074 633
rect 2108 599 2124 633
rect 2058 566 2124 599
rect 2154 633 2220 666
rect 2154 599 2170 633
rect 2204 599 2220 633
rect 2154 566 2220 599
rect 2250 633 2312 666
rect 2250 599 2266 633
rect 2300 599 2312 633
rect 2250 566 2312 599
<< pdiff >>
rect -1196 6356 -1138 6391
rect -1196 6322 -1184 6356
rect -1150 6322 -1138 6356
rect -1196 6288 -1138 6322
rect -1196 6254 -1184 6288
rect -1150 6254 -1138 6288
rect -1196 6220 -1138 6254
rect -1196 6186 -1184 6220
rect -1150 6186 -1138 6220
rect -1196 6152 -1138 6186
rect -1196 6118 -1184 6152
rect -1150 6118 -1138 6152
rect -1196 6084 -1138 6118
rect -1196 6050 -1184 6084
rect -1150 6050 -1138 6084
rect -1196 6016 -1138 6050
rect -1196 5982 -1184 6016
rect -1150 5982 -1138 6016
rect -1196 5948 -1138 5982
rect -1196 5914 -1184 5948
rect -1150 5914 -1138 5948
rect -1196 5880 -1138 5914
rect -1196 5846 -1184 5880
rect -1150 5846 -1138 5880
rect -1196 5812 -1138 5846
rect -1196 5778 -1184 5812
rect -1150 5778 -1138 5812
rect -1196 5744 -1138 5778
rect -1196 5710 -1184 5744
rect -1150 5710 -1138 5744
rect -1196 5676 -1138 5710
rect -1196 5642 -1184 5676
rect -1150 5642 -1138 5676
rect -1196 5608 -1138 5642
rect -1196 5574 -1184 5608
rect -1150 5574 -1138 5608
rect -1196 5540 -1138 5574
rect -1196 5506 -1184 5540
rect -1150 5506 -1138 5540
rect -1196 5472 -1138 5506
rect -1196 5438 -1184 5472
rect -1150 5438 -1138 5472
rect -1196 5404 -1138 5438
rect -1196 5370 -1184 5404
rect -1150 5370 -1138 5404
rect -1196 5336 -1138 5370
rect -1196 5302 -1184 5336
rect -1150 5302 -1138 5336
rect -1196 5268 -1138 5302
rect -1196 5234 -1184 5268
rect -1150 5234 -1138 5268
rect -1196 5200 -1138 5234
rect -1196 5166 -1184 5200
rect -1150 5166 -1138 5200
rect -1196 5132 -1138 5166
rect -1196 5098 -1184 5132
rect -1150 5098 -1138 5132
rect -1196 5064 -1138 5098
rect -1196 5030 -1184 5064
rect -1150 5030 -1138 5064
rect -1196 4996 -1138 5030
rect -1196 4962 -1184 4996
rect -1150 4962 -1138 4996
rect -1196 4928 -1138 4962
rect -1196 4894 -1184 4928
rect -1150 4894 -1138 4928
rect -1196 4860 -1138 4894
rect -1196 4826 -1184 4860
rect -1150 4826 -1138 4860
rect -1196 4791 -1138 4826
rect -738 6356 -680 6391
rect -738 6322 -726 6356
rect -692 6322 -680 6356
rect -738 6288 -680 6322
rect -738 6254 -726 6288
rect -692 6254 -680 6288
rect -738 6220 -680 6254
rect -738 6186 -726 6220
rect -692 6186 -680 6220
rect -738 6152 -680 6186
rect -738 6118 -726 6152
rect -692 6118 -680 6152
rect -738 6084 -680 6118
rect -738 6050 -726 6084
rect -692 6050 -680 6084
rect -738 6016 -680 6050
rect -738 5982 -726 6016
rect -692 5982 -680 6016
rect -738 5948 -680 5982
rect -738 5914 -726 5948
rect -692 5914 -680 5948
rect -738 5880 -680 5914
rect -738 5846 -726 5880
rect -692 5846 -680 5880
rect -738 5812 -680 5846
rect -738 5778 -726 5812
rect -692 5778 -680 5812
rect -738 5744 -680 5778
rect -738 5710 -726 5744
rect -692 5710 -680 5744
rect -738 5676 -680 5710
rect -738 5642 -726 5676
rect -692 5642 -680 5676
rect -738 5608 -680 5642
rect -738 5574 -726 5608
rect -692 5574 -680 5608
rect -738 5540 -680 5574
rect -738 5506 -726 5540
rect -692 5506 -680 5540
rect -738 5472 -680 5506
rect -738 5438 -726 5472
rect -692 5438 -680 5472
rect -738 5404 -680 5438
rect -738 5370 -726 5404
rect -692 5370 -680 5404
rect -738 5336 -680 5370
rect -738 5302 -726 5336
rect -692 5302 -680 5336
rect -738 5268 -680 5302
rect -738 5234 -726 5268
rect -692 5234 -680 5268
rect -738 5200 -680 5234
rect -738 5166 -726 5200
rect -692 5166 -680 5200
rect -738 5132 -680 5166
rect -738 5098 -726 5132
rect -692 5098 -680 5132
rect -738 5064 -680 5098
rect -738 5030 -726 5064
rect -692 5030 -680 5064
rect -738 4996 -680 5030
rect -738 4962 -726 4996
rect -692 4962 -680 4996
rect -738 4928 -680 4962
rect -738 4894 -726 4928
rect -692 4894 -680 4928
rect -738 4860 -680 4894
rect -738 4826 -726 4860
rect -692 4826 -680 4860
rect -738 4791 -680 4826
rect -280 6356 -222 6391
rect -280 6322 -268 6356
rect -234 6322 -222 6356
rect -280 6288 -222 6322
rect -280 6254 -268 6288
rect -234 6254 -222 6288
rect -280 6220 -222 6254
rect -280 6186 -268 6220
rect -234 6186 -222 6220
rect -280 6152 -222 6186
rect -280 6118 -268 6152
rect -234 6118 -222 6152
rect -280 6084 -222 6118
rect -280 6050 -268 6084
rect -234 6050 -222 6084
rect -280 6016 -222 6050
rect -280 5982 -268 6016
rect -234 5982 -222 6016
rect -280 5948 -222 5982
rect -280 5914 -268 5948
rect -234 5914 -222 5948
rect -280 5880 -222 5914
rect -280 5846 -268 5880
rect -234 5846 -222 5880
rect -280 5812 -222 5846
rect -280 5778 -268 5812
rect -234 5778 -222 5812
rect -280 5744 -222 5778
rect -280 5710 -268 5744
rect -234 5710 -222 5744
rect -280 5676 -222 5710
rect -280 5642 -268 5676
rect -234 5642 -222 5676
rect -280 5608 -222 5642
rect -280 5574 -268 5608
rect -234 5574 -222 5608
rect -280 5540 -222 5574
rect -280 5506 -268 5540
rect -234 5506 -222 5540
rect -280 5472 -222 5506
rect -280 5438 -268 5472
rect -234 5438 -222 5472
rect -280 5404 -222 5438
rect -280 5370 -268 5404
rect -234 5370 -222 5404
rect -280 5336 -222 5370
rect -280 5302 -268 5336
rect -234 5302 -222 5336
rect -280 5268 -222 5302
rect -280 5234 -268 5268
rect -234 5234 -222 5268
rect -280 5200 -222 5234
rect -280 5166 -268 5200
rect -234 5166 -222 5200
rect -280 5132 -222 5166
rect -280 5098 -268 5132
rect -234 5098 -222 5132
rect -280 5064 -222 5098
rect -280 5030 -268 5064
rect -234 5030 -222 5064
rect -280 4996 -222 5030
rect -280 4962 -268 4996
rect -234 4962 -222 4996
rect -280 4928 -222 4962
rect -280 4894 -268 4928
rect -234 4894 -222 4928
rect -280 4860 -222 4894
rect -280 4826 -268 4860
rect -234 4826 -222 4860
rect -280 4791 -222 4826
rect 178 6356 236 6391
rect 178 6322 190 6356
rect 224 6322 236 6356
rect 178 6288 236 6322
rect 178 6254 190 6288
rect 224 6254 236 6288
rect 178 6220 236 6254
rect 178 6186 190 6220
rect 224 6186 236 6220
rect 178 6152 236 6186
rect 178 6118 190 6152
rect 224 6118 236 6152
rect 178 6084 236 6118
rect 178 6050 190 6084
rect 224 6050 236 6084
rect 178 6016 236 6050
rect 178 5982 190 6016
rect 224 5982 236 6016
rect 178 5948 236 5982
rect 178 5914 190 5948
rect 224 5914 236 5948
rect 178 5880 236 5914
rect 178 5846 190 5880
rect 224 5846 236 5880
rect 178 5812 236 5846
rect 178 5778 190 5812
rect 224 5778 236 5812
rect 178 5744 236 5778
rect 178 5710 190 5744
rect 224 5710 236 5744
rect 178 5676 236 5710
rect 178 5642 190 5676
rect 224 5642 236 5676
rect 178 5608 236 5642
rect 178 5574 190 5608
rect 224 5574 236 5608
rect 178 5540 236 5574
rect 178 5506 190 5540
rect 224 5506 236 5540
rect 178 5472 236 5506
rect 178 5438 190 5472
rect 224 5438 236 5472
rect 178 5404 236 5438
rect 178 5370 190 5404
rect 224 5370 236 5404
rect 178 5336 236 5370
rect 178 5302 190 5336
rect 224 5302 236 5336
rect 178 5268 236 5302
rect 178 5234 190 5268
rect 224 5234 236 5268
rect 178 5200 236 5234
rect 178 5166 190 5200
rect 224 5166 236 5200
rect 178 5132 236 5166
rect 178 5098 190 5132
rect 224 5098 236 5132
rect 178 5064 236 5098
rect 178 5030 190 5064
rect 224 5030 236 5064
rect 178 4996 236 5030
rect 178 4962 190 4996
rect 224 4962 236 4996
rect 178 4928 236 4962
rect 178 4894 190 4928
rect 224 4894 236 4928
rect 178 4860 236 4894
rect 178 4826 190 4860
rect 224 4826 236 4860
rect 178 4791 236 4826
rect 636 6356 694 6391
rect 636 6322 648 6356
rect 682 6322 694 6356
rect 636 6288 694 6322
rect 636 6254 648 6288
rect 682 6254 694 6288
rect 636 6220 694 6254
rect 636 6186 648 6220
rect 682 6186 694 6220
rect 636 6152 694 6186
rect 636 6118 648 6152
rect 682 6118 694 6152
rect 636 6084 694 6118
rect 636 6050 648 6084
rect 682 6050 694 6084
rect 636 6016 694 6050
rect 636 5982 648 6016
rect 682 5982 694 6016
rect 636 5948 694 5982
rect 636 5914 648 5948
rect 682 5914 694 5948
rect 636 5880 694 5914
rect 636 5846 648 5880
rect 682 5846 694 5880
rect 636 5812 694 5846
rect 636 5778 648 5812
rect 682 5778 694 5812
rect 636 5744 694 5778
rect 636 5710 648 5744
rect 682 5710 694 5744
rect 636 5676 694 5710
rect 636 5642 648 5676
rect 682 5642 694 5676
rect 636 5608 694 5642
rect 636 5574 648 5608
rect 682 5574 694 5608
rect 636 5540 694 5574
rect 636 5506 648 5540
rect 682 5506 694 5540
rect 636 5472 694 5506
rect 636 5438 648 5472
rect 682 5438 694 5472
rect 636 5404 694 5438
rect 636 5370 648 5404
rect 682 5370 694 5404
rect 636 5336 694 5370
rect 636 5302 648 5336
rect 682 5302 694 5336
rect 636 5268 694 5302
rect 636 5234 648 5268
rect 682 5234 694 5268
rect 636 5200 694 5234
rect 636 5166 648 5200
rect 682 5166 694 5200
rect 636 5132 694 5166
rect 636 5098 648 5132
rect 682 5098 694 5132
rect 636 5064 694 5098
rect 636 5030 648 5064
rect 682 5030 694 5064
rect 636 4996 694 5030
rect 636 4962 648 4996
rect 682 4962 694 4996
rect 636 4928 694 4962
rect 636 4894 648 4928
rect 682 4894 694 4928
rect 636 4860 694 4894
rect 636 4826 648 4860
rect 682 4826 694 4860
rect 636 4791 694 4826
rect 1094 6356 1152 6391
rect 1094 6322 1106 6356
rect 1140 6322 1152 6356
rect 1094 6288 1152 6322
rect 1094 6254 1106 6288
rect 1140 6254 1152 6288
rect 1094 6220 1152 6254
rect 1094 6186 1106 6220
rect 1140 6186 1152 6220
rect 1094 6152 1152 6186
rect 1094 6118 1106 6152
rect 1140 6118 1152 6152
rect 1094 6084 1152 6118
rect 1094 6050 1106 6084
rect 1140 6050 1152 6084
rect 1094 6016 1152 6050
rect 1094 5982 1106 6016
rect 1140 5982 1152 6016
rect 1094 5948 1152 5982
rect 1094 5914 1106 5948
rect 1140 5914 1152 5948
rect 1094 5880 1152 5914
rect 1094 5846 1106 5880
rect 1140 5846 1152 5880
rect 1094 5812 1152 5846
rect 1094 5778 1106 5812
rect 1140 5778 1152 5812
rect 1094 5744 1152 5778
rect 1094 5710 1106 5744
rect 1140 5710 1152 5744
rect 1094 5676 1152 5710
rect 1094 5642 1106 5676
rect 1140 5642 1152 5676
rect 1094 5608 1152 5642
rect 1094 5574 1106 5608
rect 1140 5574 1152 5608
rect 1094 5540 1152 5574
rect 1094 5506 1106 5540
rect 1140 5506 1152 5540
rect 1094 5472 1152 5506
rect 1094 5438 1106 5472
rect 1140 5438 1152 5472
rect 1094 5404 1152 5438
rect 1094 5370 1106 5404
rect 1140 5370 1152 5404
rect 1094 5336 1152 5370
rect 1094 5302 1106 5336
rect 1140 5302 1152 5336
rect 1094 5268 1152 5302
rect 1094 5234 1106 5268
rect 1140 5234 1152 5268
rect 1094 5200 1152 5234
rect 1094 5166 1106 5200
rect 1140 5166 1152 5200
rect 1094 5132 1152 5166
rect 1094 5098 1106 5132
rect 1140 5098 1152 5132
rect 1094 5064 1152 5098
rect 1094 5030 1106 5064
rect 1140 5030 1152 5064
rect 1094 4996 1152 5030
rect 1094 4962 1106 4996
rect 1140 4962 1152 4996
rect 1094 4928 1152 4962
rect 1094 4894 1106 4928
rect 1140 4894 1152 4928
rect 1094 4860 1152 4894
rect 1094 4826 1106 4860
rect 1140 4826 1152 4860
rect 1094 4791 1152 4826
rect -1196 4318 -1138 4353
rect -1196 4284 -1184 4318
rect -1150 4284 -1138 4318
rect -1196 4250 -1138 4284
rect -1196 4216 -1184 4250
rect -1150 4216 -1138 4250
rect -1196 4182 -1138 4216
rect -1196 4148 -1184 4182
rect -1150 4148 -1138 4182
rect -1196 4114 -1138 4148
rect -1196 4080 -1184 4114
rect -1150 4080 -1138 4114
rect -1196 4046 -1138 4080
rect -1196 4012 -1184 4046
rect -1150 4012 -1138 4046
rect -1196 3978 -1138 4012
rect -1196 3944 -1184 3978
rect -1150 3944 -1138 3978
rect -1196 3910 -1138 3944
rect -1196 3876 -1184 3910
rect -1150 3876 -1138 3910
rect -1196 3842 -1138 3876
rect -1196 3808 -1184 3842
rect -1150 3808 -1138 3842
rect -1196 3774 -1138 3808
rect -1196 3740 -1184 3774
rect -1150 3740 -1138 3774
rect -1196 3706 -1138 3740
rect -1196 3672 -1184 3706
rect -1150 3672 -1138 3706
rect -1196 3638 -1138 3672
rect -1196 3604 -1184 3638
rect -1150 3604 -1138 3638
rect -1196 3570 -1138 3604
rect -1196 3536 -1184 3570
rect -1150 3536 -1138 3570
rect -1196 3502 -1138 3536
rect -1196 3468 -1184 3502
rect -1150 3468 -1138 3502
rect -1196 3434 -1138 3468
rect -1196 3400 -1184 3434
rect -1150 3400 -1138 3434
rect -1196 3366 -1138 3400
rect -1196 3332 -1184 3366
rect -1150 3332 -1138 3366
rect -1196 3298 -1138 3332
rect -1196 3264 -1184 3298
rect -1150 3264 -1138 3298
rect -1196 3230 -1138 3264
rect -1196 3196 -1184 3230
rect -1150 3196 -1138 3230
rect -1196 3162 -1138 3196
rect -1196 3128 -1184 3162
rect -1150 3128 -1138 3162
rect -1196 3094 -1138 3128
rect -1196 3060 -1184 3094
rect -1150 3060 -1138 3094
rect -1196 3026 -1138 3060
rect -1196 2992 -1184 3026
rect -1150 2992 -1138 3026
rect -1196 2958 -1138 2992
rect -1196 2924 -1184 2958
rect -1150 2924 -1138 2958
rect -1196 2890 -1138 2924
rect -1196 2856 -1184 2890
rect -1150 2856 -1138 2890
rect -1196 2822 -1138 2856
rect -1196 2788 -1184 2822
rect -1150 2788 -1138 2822
rect -1196 2753 -1138 2788
rect -738 4318 -680 4353
rect -738 4284 -726 4318
rect -692 4284 -680 4318
rect -738 4250 -680 4284
rect -738 4216 -726 4250
rect -692 4216 -680 4250
rect -738 4182 -680 4216
rect -738 4148 -726 4182
rect -692 4148 -680 4182
rect -738 4114 -680 4148
rect -738 4080 -726 4114
rect -692 4080 -680 4114
rect -738 4046 -680 4080
rect -738 4012 -726 4046
rect -692 4012 -680 4046
rect -738 3978 -680 4012
rect -738 3944 -726 3978
rect -692 3944 -680 3978
rect -738 3910 -680 3944
rect -738 3876 -726 3910
rect -692 3876 -680 3910
rect -738 3842 -680 3876
rect -738 3808 -726 3842
rect -692 3808 -680 3842
rect -738 3774 -680 3808
rect -738 3740 -726 3774
rect -692 3740 -680 3774
rect -738 3706 -680 3740
rect -738 3672 -726 3706
rect -692 3672 -680 3706
rect -738 3638 -680 3672
rect -738 3604 -726 3638
rect -692 3604 -680 3638
rect -738 3570 -680 3604
rect -738 3536 -726 3570
rect -692 3536 -680 3570
rect -738 3502 -680 3536
rect -738 3468 -726 3502
rect -692 3468 -680 3502
rect -738 3434 -680 3468
rect -738 3400 -726 3434
rect -692 3400 -680 3434
rect -738 3366 -680 3400
rect -738 3332 -726 3366
rect -692 3332 -680 3366
rect -738 3298 -680 3332
rect -738 3264 -726 3298
rect -692 3264 -680 3298
rect -738 3230 -680 3264
rect -738 3196 -726 3230
rect -692 3196 -680 3230
rect -738 3162 -680 3196
rect -738 3128 -726 3162
rect -692 3128 -680 3162
rect -738 3094 -680 3128
rect -738 3060 -726 3094
rect -692 3060 -680 3094
rect -738 3026 -680 3060
rect -738 2992 -726 3026
rect -692 2992 -680 3026
rect -738 2958 -680 2992
rect -738 2924 -726 2958
rect -692 2924 -680 2958
rect -738 2890 -680 2924
rect -738 2856 -726 2890
rect -692 2856 -680 2890
rect -738 2822 -680 2856
rect -738 2788 -726 2822
rect -692 2788 -680 2822
rect -738 2753 -680 2788
rect -280 4318 -222 4353
rect -280 4284 -268 4318
rect -234 4284 -222 4318
rect -280 4250 -222 4284
rect -280 4216 -268 4250
rect -234 4216 -222 4250
rect -280 4182 -222 4216
rect -280 4148 -268 4182
rect -234 4148 -222 4182
rect -280 4114 -222 4148
rect -280 4080 -268 4114
rect -234 4080 -222 4114
rect -280 4046 -222 4080
rect -280 4012 -268 4046
rect -234 4012 -222 4046
rect -280 3978 -222 4012
rect -280 3944 -268 3978
rect -234 3944 -222 3978
rect -280 3910 -222 3944
rect -280 3876 -268 3910
rect -234 3876 -222 3910
rect -280 3842 -222 3876
rect -280 3808 -268 3842
rect -234 3808 -222 3842
rect -280 3774 -222 3808
rect -280 3740 -268 3774
rect -234 3740 -222 3774
rect -280 3706 -222 3740
rect -280 3672 -268 3706
rect -234 3672 -222 3706
rect -280 3638 -222 3672
rect -280 3604 -268 3638
rect -234 3604 -222 3638
rect -280 3570 -222 3604
rect -280 3536 -268 3570
rect -234 3536 -222 3570
rect -280 3502 -222 3536
rect -280 3468 -268 3502
rect -234 3468 -222 3502
rect -280 3434 -222 3468
rect -280 3400 -268 3434
rect -234 3400 -222 3434
rect -280 3366 -222 3400
rect -280 3332 -268 3366
rect -234 3332 -222 3366
rect -280 3298 -222 3332
rect -280 3264 -268 3298
rect -234 3264 -222 3298
rect -280 3230 -222 3264
rect -280 3196 -268 3230
rect -234 3196 -222 3230
rect -280 3162 -222 3196
rect -280 3128 -268 3162
rect -234 3128 -222 3162
rect -280 3094 -222 3128
rect -280 3060 -268 3094
rect -234 3060 -222 3094
rect -280 3026 -222 3060
rect -280 2992 -268 3026
rect -234 2992 -222 3026
rect -280 2958 -222 2992
rect -280 2924 -268 2958
rect -234 2924 -222 2958
rect -280 2890 -222 2924
rect -280 2856 -268 2890
rect -234 2856 -222 2890
rect -280 2822 -222 2856
rect -280 2788 -268 2822
rect -234 2788 -222 2822
rect -280 2753 -222 2788
rect 178 4318 236 4353
rect 178 4284 190 4318
rect 224 4284 236 4318
rect 178 4250 236 4284
rect 178 4216 190 4250
rect 224 4216 236 4250
rect 178 4182 236 4216
rect 178 4148 190 4182
rect 224 4148 236 4182
rect 178 4114 236 4148
rect 178 4080 190 4114
rect 224 4080 236 4114
rect 178 4046 236 4080
rect 178 4012 190 4046
rect 224 4012 236 4046
rect 178 3978 236 4012
rect 178 3944 190 3978
rect 224 3944 236 3978
rect 178 3910 236 3944
rect 178 3876 190 3910
rect 224 3876 236 3910
rect 178 3842 236 3876
rect 178 3808 190 3842
rect 224 3808 236 3842
rect 178 3774 236 3808
rect 178 3740 190 3774
rect 224 3740 236 3774
rect 178 3706 236 3740
rect 178 3672 190 3706
rect 224 3672 236 3706
rect 178 3638 236 3672
rect 178 3604 190 3638
rect 224 3604 236 3638
rect 178 3570 236 3604
rect 178 3536 190 3570
rect 224 3536 236 3570
rect 178 3502 236 3536
rect 178 3468 190 3502
rect 224 3468 236 3502
rect 178 3434 236 3468
rect 178 3400 190 3434
rect 224 3400 236 3434
rect 178 3366 236 3400
rect 178 3332 190 3366
rect 224 3332 236 3366
rect 178 3298 236 3332
rect 178 3264 190 3298
rect 224 3264 236 3298
rect 178 3230 236 3264
rect 178 3196 190 3230
rect 224 3196 236 3230
rect 178 3162 236 3196
rect 178 3128 190 3162
rect 224 3128 236 3162
rect 178 3094 236 3128
rect 178 3060 190 3094
rect 224 3060 236 3094
rect 178 3026 236 3060
rect 178 2992 190 3026
rect 224 2992 236 3026
rect 178 2958 236 2992
rect 178 2924 190 2958
rect 224 2924 236 2958
rect 178 2890 236 2924
rect 178 2856 190 2890
rect 224 2856 236 2890
rect 178 2822 236 2856
rect 178 2788 190 2822
rect 224 2788 236 2822
rect 178 2753 236 2788
rect 636 4318 694 4353
rect 636 4284 648 4318
rect 682 4284 694 4318
rect 636 4250 694 4284
rect 636 4216 648 4250
rect 682 4216 694 4250
rect 636 4182 694 4216
rect 636 4148 648 4182
rect 682 4148 694 4182
rect 636 4114 694 4148
rect 636 4080 648 4114
rect 682 4080 694 4114
rect 636 4046 694 4080
rect 636 4012 648 4046
rect 682 4012 694 4046
rect 636 3978 694 4012
rect 636 3944 648 3978
rect 682 3944 694 3978
rect 636 3910 694 3944
rect 636 3876 648 3910
rect 682 3876 694 3910
rect 636 3842 694 3876
rect 636 3808 648 3842
rect 682 3808 694 3842
rect 636 3774 694 3808
rect 636 3740 648 3774
rect 682 3740 694 3774
rect 636 3706 694 3740
rect 636 3672 648 3706
rect 682 3672 694 3706
rect 636 3638 694 3672
rect 636 3604 648 3638
rect 682 3604 694 3638
rect 636 3570 694 3604
rect 636 3536 648 3570
rect 682 3536 694 3570
rect 636 3502 694 3536
rect 636 3468 648 3502
rect 682 3468 694 3502
rect 636 3434 694 3468
rect 636 3400 648 3434
rect 682 3400 694 3434
rect 636 3366 694 3400
rect 636 3332 648 3366
rect 682 3332 694 3366
rect 636 3298 694 3332
rect 636 3264 648 3298
rect 682 3264 694 3298
rect 636 3230 694 3264
rect 636 3196 648 3230
rect 682 3196 694 3230
rect 636 3162 694 3196
rect 636 3128 648 3162
rect 682 3128 694 3162
rect 636 3094 694 3128
rect 636 3060 648 3094
rect 682 3060 694 3094
rect 636 3026 694 3060
rect 636 2992 648 3026
rect 682 2992 694 3026
rect 636 2958 694 2992
rect 636 2924 648 2958
rect 682 2924 694 2958
rect 636 2890 694 2924
rect 636 2856 648 2890
rect 682 2856 694 2890
rect 636 2822 694 2856
rect 636 2788 648 2822
rect 682 2788 694 2822
rect 636 2753 694 2788
rect 1094 4318 1152 4353
rect 1094 4284 1106 4318
rect 1140 4284 1152 4318
rect 1094 4250 1152 4284
rect 1094 4216 1106 4250
rect 1140 4216 1152 4250
rect 1094 4182 1152 4216
rect 1094 4148 1106 4182
rect 1140 4148 1152 4182
rect 1094 4114 1152 4148
rect 1094 4080 1106 4114
rect 1140 4080 1152 4114
rect 1094 4046 1152 4080
rect 1094 4012 1106 4046
rect 1140 4012 1152 4046
rect 1094 3978 1152 4012
rect 1094 3944 1106 3978
rect 1140 3944 1152 3978
rect 1094 3910 1152 3944
rect 1094 3876 1106 3910
rect 1140 3876 1152 3910
rect 1094 3842 1152 3876
rect 1094 3808 1106 3842
rect 1140 3808 1152 3842
rect 1094 3774 1152 3808
rect 1094 3740 1106 3774
rect 1140 3740 1152 3774
rect 1094 3706 1152 3740
rect 1094 3672 1106 3706
rect 1140 3672 1152 3706
rect 1094 3638 1152 3672
rect 1094 3604 1106 3638
rect 1140 3604 1152 3638
rect 1094 3570 1152 3604
rect 1094 3536 1106 3570
rect 1140 3536 1152 3570
rect 1094 3502 1152 3536
rect 1094 3468 1106 3502
rect 1140 3468 1152 3502
rect 1094 3434 1152 3468
rect 1094 3400 1106 3434
rect 1140 3400 1152 3434
rect 1094 3366 1152 3400
rect 1094 3332 1106 3366
rect 1140 3332 1152 3366
rect 1094 3298 1152 3332
rect 1094 3264 1106 3298
rect 1140 3264 1152 3298
rect 1094 3230 1152 3264
rect 1094 3196 1106 3230
rect 1140 3196 1152 3230
rect 1094 3162 1152 3196
rect 1094 3128 1106 3162
rect 1140 3128 1152 3162
rect 1094 3094 1152 3128
rect 1094 3060 1106 3094
rect 1140 3060 1152 3094
rect 1094 3026 1152 3060
rect 1094 2992 1106 3026
rect 1140 2992 1152 3026
rect 1094 2958 1152 2992
rect 1094 2924 1106 2958
rect 1140 2924 1152 2958
rect 1094 2890 1152 2924
rect 1094 2856 1106 2890
rect 1140 2856 1152 2890
rect 1094 2822 1152 2856
rect 1094 2788 1106 2822
rect 1140 2788 1152 2822
rect 1094 2753 1152 2788
<< ndiffc >>
rect 16 1631 50 1665
rect 112 1631 146 1665
rect 208 1631 242 1665
rect 304 1631 338 1665
rect 400 1631 434 1665
rect 496 1631 530 1665
rect 592 1631 626 1665
rect 688 1631 722 1665
rect 784 1631 818 1665
rect 880 1631 914 1665
rect 976 1631 1010 1665
rect 1310 1631 1344 1665
rect 1406 1631 1440 1665
rect 1502 1631 1536 1665
rect 1598 1631 1632 1665
rect 1694 1631 1728 1665
rect 1790 1631 1824 1665
rect 1886 1631 1920 1665
rect 1982 1631 2016 1665
rect 2078 1631 2112 1665
rect 2174 1631 2208 1665
rect 2270 1631 2304 1665
rect 1306 599 1340 633
rect 1402 599 1436 633
rect 1498 599 1532 633
rect 1594 599 1628 633
rect 1690 599 1724 633
rect 1786 599 1820 633
rect 1882 599 1916 633
rect 1978 599 2012 633
rect 2074 599 2108 633
rect 2170 599 2204 633
rect 2266 599 2300 633
<< pdiffc >>
rect -1184 6322 -1150 6356
rect -1184 6254 -1150 6288
rect -1184 6186 -1150 6220
rect -1184 6118 -1150 6152
rect -1184 6050 -1150 6084
rect -1184 5982 -1150 6016
rect -1184 5914 -1150 5948
rect -1184 5846 -1150 5880
rect -1184 5778 -1150 5812
rect -1184 5710 -1150 5744
rect -1184 5642 -1150 5676
rect -1184 5574 -1150 5608
rect -1184 5506 -1150 5540
rect -1184 5438 -1150 5472
rect -1184 5370 -1150 5404
rect -1184 5302 -1150 5336
rect -1184 5234 -1150 5268
rect -1184 5166 -1150 5200
rect -1184 5098 -1150 5132
rect -1184 5030 -1150 5064
rect -1184 4962 -1150 4996
rect -1184 4894 -1150 4928
rect -1184 4826 -1150 4860
rect -726 6322 -692 6356
rect -726 6254 -692 6288
rect -726 6186 -692 6220
rect -726 6118 -692 6152
rect -726 6050 -692 6084
rect -726 5982 -692 6016
rect -726 5914 -692 5948
rect -726 5846 -692 5880
rect -726 5778 -692 5812
rect -726 5710 -692 5744
rect -726 5642 -692 5676
rect -726 5574 -692 5608
rect -726 5506 -692 5540
rect -726 5438 -692 5472
rect -726 5370 -692 5404
rect -726 5302 -692 5336
rect -726 5234 -692 5268
rect -726 5166 -692 5200
rect -726 5098 -692 5132
rect -726 5030 -692 5064
rect -726 4962 -692 4996
rect -726 4894 -692 4928
rect -726 4826 -692 4860
rect -268 6322 -234 6356
rect -268 6254 -234 6288
rect -268 6186 -234 6220
rect -268 6118 -234 6152
rect -268 6050 -234 6084
rect -268 5982 -234 6016
rect -268 5914 -234 5948
rect -268 5846 -234 5880
rect -268 5778 -234 5812
rect -268 5710 -234 5744
rect -268 5642 -234 5676
rect -268 5574 -234 5608
rect -268 5506 -234 5540
rect -268 5438 -234 5472
rect -268 5370 -234 5404
rect -268 5302 -234 5336
rect -268 5234 -234 5268
rect -268 5166 -234 5200
rect -268 5098 -234 5132
rect -268 5030 -234 5064
rect -268 4962 -234 4996
rect -268 4894 -234 4928
rect -268 4826 -234 4860
rect 190 6322 224 6356
rect 190 6254 224 6288
rect 190 6186 224 6220
rect 190 6118 224 6152
rect 190 6050 224 6084
rect 190 5982 224 6016
rect 190 5914 224 5948
rect 190 5846 224 5880
rect 190 5778 224 5812
rect 190 5710 224 5744
rect 190 5642 224 5676
rect 190 5574 224 5608
rect 190 5506 224 5540
rect 190 5438 224 5472
rect 190 5370 224 5404
rect 190 5302 224 5336
rect 190 5234 224 5268
rect 190 5166 224 5200
rect 190 5098 224 5132
rect 190 5030 224 5064
rect 190 4962 224 4996
rect 190 4894 224 4928
rect 190 4826 224 4860
rect 648 6322 682 6356
rect 648 6254 682 6288
rect 648 6186 682 6220
rect 648 6118 682 6152
rect 648 6050 682 6084
rect 648 5982 682 6016
rect 648 5914 682 5948
rect 648 5846 682 5880
rect 648 5778 682 5812
rect 648 5710 682 5744
rect 648 5642 682 5676
rect 648 5574 682 5608
rect 648 5506 682 5540
rect 648 5438 682 5472
rect 648 5370 682 5404
rect 648 5302 682 5336
rect 648 5234 682 5268
rect 648 5166 682 5200
rect 648 5098 682 5132
rect 648 5030 682 5064
rect 648 4962 682 4996
rect 648 4894 682 4928
rect 648 4826 682 4860
rect 1106 6322 1140 6356
rect 1106 6254 1140 6288
rect 1106 6186 1140 6220
rect 1106 6118 1140 6152
rect 1106 6050 1140 6084
rect 1106 5982 1140 6016
rect 1106 5914 1140 5948
rect 1106 5846 1140 5880
rect 1106 5778 1140 5812
rect 1106 5710 1140 5744
rect 1106 5642 1140 5676
rect 1106 5574 1140 5608
rect 1106 5506 1140 5540
rect 1106 5438 1140 5472
rect 1106 5370 1140 5404
rect 1106 5302 1140 5336
rect 1106 5234 1140 5268
rect 1106 5166 1140 5200
rect 1106 5098 1140 5132
rect 1106 5030 1140 5064
rect 1106 4962 1140 4996
rect 1106 4894 1140 4928
rect 1106 4826 1140 4860
rect -1184 4284 -1150 4318
rect -1184 4216 -1150 4250
rect -1184 4148 -1150 4182
rect -1184 4080 -1150 4114
rect -1184 4012 -1150 4046
rect -1184 3944 -1150 3978
rect -1184 3876 -1150 3910
rect -1184 3808 -1150 3842
rect -1184 3740 -1150 3774
rect -1184 3672 -1150 3706
rect -1184 3604 -1150 3638
rect -1184 3536 -1150 3570
rect -1184 3468 -1150 3502
rect -1184 3400 -1150 3434
rect -1184 3332 -1150 3366
rect -1184 3264 -1150 3298
rect -1184 3196 -1150 3230
rect -1184 3128 -1150 3162
rect -1184 3060 -1150 3094
rect -1184 2992 -1150 3026
rect -1184 2924 -1150 2958
rect -1184 2856 -1150 2890
rect -1184 2788 -1150 2822
rect -726 4284 -692 4318
rect -726 4216 -692 4250
rect -726 4148 -692 4182
rect -726 4080 -692 4114
rect -726 4012 -692 4046
rect -726 3944 -692 3978
rect -726 3876 -692 3910
rect -726 3808 -692 3842
rect -726 3740 -692 3774
rect -726 3672 -692 3706
rect -726 3604 -692 3638
rect -726 3536 -692 3570
rect -726 3468 -692 3502
rect -726 3400 -692 3434
rect -726 3332 -692 3366
rect -726 3264 -692 3298
rect -726 3196 -692 3230
rect -726 3128 -692 3162
rect -726 3060 -692 3094
rect -726 2992 -692 3026
rect -726 2924 -692 2958
rect -726 2856 -692 2890
rect -726 2788 -692 2822
rect -268 4284 -234 4318
rect -268 4216 -234 4250
rect -268 4148 -234 4182
rect -268 4080 -234 4114
rect -268 4012 -234 4046
rect -268 3944 -234 3978
rect -268 3876 -234 3910
rect -268 3808 -234 3842
rect -268 3740 -234 3774
rect -268 3672 -234 3706
rect -268 3604 -234 3638
rect -268 3536 -234 3570
rect -268 3468 -234 3502
rect -268 3400 -234 3434
rect -268 3332 -234 3366
rect -268 3264 -234 3298
rect -268 3196 -234 3230
rect -268 3128 -234 3162
rect -268 3060 -234 3094
rect -268 2992 -234 3026
rect -268 2924 -234 2958
rect -268 2856 -234 2890
rect -268 2788 -234 2822
rect 190 4284 224 4318
rect 190 4216 224 4250
rect 190 4148 224 4182
rect 190 4080 224 4114
rect 190 4012 224 4046
rect 190 3944 224 3978
rect 190 3876 224 3910
rect 190 3808 224 3842
rect 190 3740 224 3774
rect 190 3672 224 3706
rect 190 3604 224 3638
rect 190 3536 224 3570
rect 190 3468 224 3502
rect 190 3400 224 3434
rect 190 3332 224 3366
rect 190 3264 224 3298
rect 190 3196 224 3230
rect 190 3128 224 3162
rect 190 3060 224 3094
rect 190 2992 224 3026
rect 190 2924 224 2958
rect 190 2856 224 2890
rect 190 2788 224 2822
rect 648 4284 682 4318
rect 648 4216 682 4250
rect 648 4148 682 4182
rect 648 4080 682 4114
rect 648 4012 682 4046
rect 648 3944 682 3978
rect 648 3876 682 3910
rect 648 3808 682 3842
rect 648 3740 682 3774
rect 648 3672 682 3706
rect 648 3604 682 3638
rect 648 3536 682 3570
rect 648 3468 682 3502
rect 648 3400 682 3434
rect 648 3332 682 3366
rect 648 3264 682 3298
rect 648 3196 682 3230
rect 648 3128 682 3162
rect 648 3060 682 3094
rect 648 2992 682 3026
rect 648 2924 682 2958
rect 648 2856 682 2890
rect 648 2788 682 2822
rect 1106 4284 1140 4318
rect 1106 4216 1140 4250
rect 1106 4148 1140 4182
rect 1106 4080 1140 4114
rect 1106 4012 1140 4046
rect 1106 3944 1140 3978
rect 1106 3876 1140 3910
rect 1106 3808 1140 3842
rect 1106 3740 1140 3774
rect 1106 3672 1140 3706
rect 1106 3604 1140 3638
rect 1106 3536 1140 3570
rect 1106 3468 1140 3502
rect 1106 3400 1140 3434
rect 1106 3332 1140 3366
rect 1106 3264 1140 3298
rect 1106 3196 1140 3230
rect 1106 3128 1140 3162
rect 1106 3060 1140 3094
rect 1106 2992 1140 3026
rect 1106 2924 1140 2958
rect 1106 2856 1140 2890
rect 1106 2788 1140 2822
<< psubdiff >>
rect -98 1838 20 1872
rect 54 1838 88 1872
rect 122 1838 156 1872
rect 190 1838 224 1872
rect 258 1838 292 1872
rect 326 1838 360 1872
rect 394 1838 428 1872
rect 462 1838 496 1872
rect 530 1838 564 1872
rect 598 1838 632 1872
rect 666 1838 700 1872
rect 734 1838 768 1872
rect 802 1838 836 1872
rect 870 1838 904 1872
rect 938 1838 972 1872
rect 1006 1838 1124 1872
rect -98 1767 -64 1838
rect -98 1699 -64 1733
rect 1090 1767 1124 1838
rect 1090 1699 1124 1733
rect -98 1631 -64 1665
rect 1090 1631 1124 1665
rect -98 1563 -64 1597
rect -98 1458 -64 1529
rect 1090 1563 1124 1597
rect 1090 1458 1124 1529
rect -98 1424 20 1458
rect 54 1424 88 1458
rect 122 1424 156 1458
rect 190 1424 224 1458
rect 258 1424 292 1458
rect 326 1424 360 1458
rect 394 1424 428 1458
rect 462 1424 496 1458
rect 530 1424 564 1458
rect 598 1424 632 1458
rect 666 1424 700 1458
rect 734 1424 768 1458
rect 802 1424 836 1458
rect 870 1424 904 1458
rect 938 1424 972 1458
rect 1006 1424 1124 1458
rect 1196 1838 1314 1872
rect 1348 1838 1382 1872
rect 1416 1838 1450 1872
rect 1484 1838 1518 1872
rect 1552 1838 1586 1872
rect 1620 1838 1654 1872
rect 1688 1838 1722 1872
rect 1756 1838 1790 1872
rect 1824 1838 1858 1872
rect 1892 1838 1926 1872
rect 1960 1838 1994 1872
rect 2028 1838 2062 1872
rect 2096 1838 2130 1872
rect 2164 1838 2198 1872
rect 2232 1838 2266 1872
rect 2300 1838 2418 1872
rect 1196 1767 1230 1838
rect 1196 1699 1230 1733
rect 2384 1767 2418 1838
rect 2384 1699 2418 1733
rect 1196 1631 1230 1665
rect 2384 1631 2418 1665
rect 1196 1563 1230 1597
rect 1196 1458 1230 1529
rect 2384 1563 2418 1597
rect 2384 1458 2418 1529
rect 1196 1424 1314 1458
rect 1348 1424 1382 1458
rect 1416 1424 1450 1458
rect 1484 1424 1518 1458
rect 1552 1424 1586 1458
rect 1620 1424 1654 1458
rect 1688 1424 1722 1458
rect 1756 1424 1790 1458
rect 1824 1424 1858 1458
rect 1892 1424 1926 1458
rect 1960 1424 1994 1458
rect 2028 1424 2062 1458
rect 2096 1424 2130 1458
rect 2164 1424 2198 1458
rect 2232 1424 2266 1458
rect 2300 1424 2418 1458
rect 1192 806 1310 840
rect 1344 806 1378 840
rect 1412 806 1446 840
rect 1480 806 1514 840
rect 1548 806 1582 840
rect 1616 806 1650 840
rect 1684 806 1718 840
rect 1752 806 1786 840
rect 1820 806 1854 840
rect 1888 806 1922 840
rect 1956 806 1990 840
rect 2024 806 2058 840
rect 2092 806 2126 840
rect 2160 806 2194 840
rect 2228 806 2262 840
rect 2296 806 2414 840
rect 1192 735 1226 806
rect 1192 667 1226 701
rect 2380 735 2414 806
rect 2380 667 2414 701
rect 1192 599 1226 633
rect 2380 599 2414 633
rect 1192 531 1226 565
rect 1192 426 1226 497
rect 2380 531 2414 565
rect 2380 426 2414 497
rect 1192 392 1310 426
rect 1344 392 1378 426
rect 1412 392 1446 426
rect 1480 392 1514 426
rect 1548 392 1582 426
rect 1616 392 1650 426
rect 1684 392 1718 426
rect 1752 392 1786 426
rect 1820 392 1854 426
rect 1888 392 1922 426
rect 1956 392 1990 426
rect 2024 392 2058 426
rect 2092 392 2126 426
rect 2160 392 2194 426
rect 2228 392 2262 426
rect 2296 392 2414 426
<< nsubdiff >>
rect -1298 6540 -1195 6574
rect -1161 6540 -1127 6574
rect -1093 6540 -1059 6574
rect -1025 6540 -991 6574
rect -957 6540 -923 6574
rect -889 6540 -855 6574
rect -821 6540 -787 6574
rect -753 6540 -719 6574
rect -685 6540 -651 6574
rect -617 6540 -583 6574
rect -549 6540 -515 6574
rect -481 6540 -447 6574
rect -413 6540 -379 6574
rect -345 6540 -311 6574
rect -277 6540 -243 6574
rect -209 6540 -175 6574
rect -141 6540 -107 6574
rect -73 6540 -39 6574
rect -5 6540 29 6574
rect 63 6540 97 6574
rect 131 6540 165 6574
rect 199 6540 233 6574
rect 267 6540 301 6574
rect 335 6540 369 6574
rect 403 6540 437 6574
rect 471 6540 505 6574
rect 539 6540 573 6574
rect 607 6540 641 6574
rect 675 6540 709 6574
rect 743 6540 777 6574
rect 811 6540 845 6574
rect 879 6540 913 6574
rect 947 6540 981 6574
rect 1015 6540 1049 6574
rect 1083 6540 1117 6574
rect 1151 6540 1254 6574
rect -1298 6458 -1264 6540
rect -1298 6390 -1264 6424
rect 1220 6458 1254 6540
rect -1298 6322 -1264 6356
rect -1298 6254 -1264 6288
rect -1298 6186 -1264 6220
rect -1298 6118 -1264 6152
rect -1298 6050 -1264 6084
rect -1298 5982 -1264 6016
rect -1298 5914 -1264 5948
rect -1298 5846 -1264 5880
rect -1298 5778 -1264 5812
rect -1298 5710 -1264 5744
rect -1298 5642 -1264 5676
rect -1298 5574 -1264 5608
rect -1298 5506 -1264 5540
rect -1298 5438 -1264 5472
rect -1298 5370 -1264 5404
rect -1298 5302 -1264 5336
rect -1298 5234 -1264 5268
rect -1298 5166 -1264 5200
rect -1298 5098 -1264 5132
rect -1298 5030 -1264 5064
rect -1298 4962 -1264 4996
rect -1298 4894 -1264 4928
rect -1298 4826 -1264 4860
rect -1298 4758 -1264 4792
rect 1220 6390 1254 6424
rect 1220 6322 1254 6356
rect 1220 6254 1254 6288
rect 1220 6186 1254 6220
rect 1220 6118 1254 6152
rect 1220 6050 1254 6084
rect 1220 5982 1254 6016
rect 1220 5914 1254 5948
rect 1220 5846 1254 5880
rect 1220 5778 1254 5812
rect 1220 5710 1254 5744
rect 1220 5642 1254 5676
rect 1220 5574 1254 5608
rect 1220 5506 1254 5540
rect 1220 5438 1254 5472
rect 1220 5370 1254 5404
rect 1220 5302 1254 5336
rect 1220 5234 1254 5268
rect 1220 5166 1254 5200
rect 1220 5098 1254 5132
rect 1220 5030 1254 5064
rect 1220 4962 1254 4996
rect 1220 4894 1254 4928
rect 1220 4826 1254 4860
rect -1298 4642 -1264 4724
rect 1220 4758 1254 4792
rect 1220 4642 1254 4724
rect -1298 4608 -1195 4642
rect -1161 4608 -1127 4642
rect -1093 4608 -1059 4642
rect -1025 4608 -991 4642
rect -957 4608 -923 4642
rect -889 4608 -855 4642
rect -821 4608 -787 4642
rect -753 4608 -719 4642
rect -685 4608 -651 4642
rect -617 4608 -583 4642
rect -549 4608 -515 4642
rect -481 4608 -447 4642
rect -413 4608 -379 4642
rect -345 4608 -311 4642
rect -277 4608 -243 4642
rect -209 4608 -175 4642
rect -141 4608 -107 4642
rect -73 4608 -39 4642
rect -5 4608 29 4642
rect 63 4608 97 4642
rect 131 4608 165 4642
rect 199 4608 233 4642
rect 267 4608 301 4642
rect 335 4608 369 4642
rect 403 4608 437 4642
rect 471 4608 505 4642
rect 539 4608 573 4642
rect 607 4608 641 4642
rect 675 4608 709 4642
rect 743 4608 777 4642
rect 811 4608 845 4642
rect 879 4608 913 4642
rect 947 4608 981 4642
rect 1015 4608 1049 4642
rect 1083 4608 1117 4642
rect 1151 4608 1254 4642
rect -1298 4502 -1195 4536
rect -1161 4502 -1127 4536
rect -1093 4502 -1059 4536
rect -1025 4502 -991 4536
rect -957 4502 -923 4536
rect -889 4502 -855 4536
rect -821 4502 -787 4536
rect -753 4502 -719 4536
rect -685 4502 -651 4536
rect -617 4502 -583 4536
rect -549 4502 -515 4536
rect -481 4502 -447 4536
rect -413 4502 -379 4536
rect -345 4502 -311 4536
rect -277 4502 -243 4536
rect -209 4502 -175 4536
rect -141 4502 -107 4536
rect -73 4502 -39 4536
rect -5 4502 29 4536
rect 63 4502 97 4536
rect 131 4502 165 4536
rect 199 4502 233 4536
rect 267 4502 301 4536
rect 335 4502 369 4536
rect 403 4502 437 4536
rect 471 4502 505 4536
rect 539 4502 573 4536
rect 607 4502 641 4536
rect 675 4502 709 4536
rect 743 4502 777 4536
rect 811 4502 845 4536
rect 879 4502 913 4536
rect 947 4502 981 4536
rect 1015 4502 1049 4536
rect 1083 4502 1117 4536
rect 1151 4502 1254 4536
rect -1298 4420 -1264 4502
rect -1298 4352 -1264 4386
rect 1220 4420 1254 4502
rect -1298 4284 -1264 4318
rect -1298 4216 -1264 4250
rect -1298 4148 -1264 4182
rect -1298 4080 -1264 4114
rect -1298 4012 -1264 4046
rect -1298 3944 -1264 3978
rect -1298 3876 -1264 3910
rect -1298 3808 -1264 3842
rect -1298 3740 -1264 3774
rect -1298 3672 -1264 3706
rect -1298 3604 -1264 3638
rect -1298 3536 -1264 3570
rect -1298 3468 -1264 3502
rect -1298 3400 -1264 3434
rect -1298 3332 -1264 3366
rect -1298 3264 -1264 3298
rect -1298 3196 -1264 3230
rect -1298 3128 -1264 3162
rect -1298 3060 -1264 3094
rect -1298 2992 -1264 3026
rect -1298 2924 -1264 2958
rect -1298 2856 -1264 2890
rect -1298 2788 -1264 2822
rect -1298 2720 -1264 2754
rect 1220 4352 1254 4386
rect 1220 4284 1254 4318
rect 1220 4216 1254 4250
rect 1220 4148 1254 4182
rect 1220 4080 1254 4114
rect 1220 4012 1254 4046
rect 1220 3944 1254 3978
rect 1220 3876 1254 3910
rect 1220 3808 1254 3842
rect 1220 3740 1254 3774
rect 1220 3672 1254 3706
rect 1220 3604 1254 3638
rect 1220 3536 1254 3570
rect 1220 3468 1254 3502
rect 1220 3400 1254 3434
rect 1220 3332 1254 3366
rect 1220 3264 1254 3298
rect 1220 3196 1254 3230
rect 1220 3128 1254 3162
rect 1220 3060 1254 3094
rect 1220 2992 1254 3026
rect 1220 2924 1254 2958
rect 1220 2856 1254 2890
rect 1220 2788 1254 2822
rect -1298 2604 -1264 2686
rect 1220 2720 1254 2754
rect 1220 2604 1254 2686
rect -1298 2570 -1195 2604
rect -1161 2570 -1127 2604
rect -1093 2570 -1059 2604
rect -1025 2570 -991 2604
rect -957 2570 -923 2604
rect -889 2570 -855 2604
rect -821 2570 -787 2604
rect -753 2570 -719 2604
rect -685 2570 -651 2604
rect -617 2570 -583 2604
rect -549 2570 -515 2604
rect -481 2570 -447 2604
rect -413 2570 -379 2604
rect -345 2570 -311 2604
rect -277 2570 -243 2604
rect -209 2570 -175 2604
rect -141 2570 -107 2604
rect -73 2570 -39 2604
rect -5 2570 29 2604
rect 63 2570 97 2604
rect 131 2570 165 2604
rect 199 2570 233 2604
rect 267 2570 301 2604
rect 335 2570 369 2604
rect 403 2570 437 2604
rect 471 2570 505 2604
rect 539 2570 573 2604
rect 607 2570 641 2604
rect 675 2570 709 2604
rect 743 2570 777 2604
rect 811 2570 845 2604
rect 879 2570 913 2604
rect 947 2570 981 2604
rect 1015 2570 1049 2604
rect 1083 2570 1117 2604
rect 1151 2570 1254 2604
<< psubdiffcont >>
rect 20 1838 54 1872
rect 88 1838 122 1872
rect 156 1838 190 1872
rect 224 1838 258 1872
rect 292 1838 326 1872
rect 360 1838 394 1872
rect 428 1838 462 1872
rect 496 1838 530 1872
rect 564 1838 598 1872
rect 632 1838 666 1872
rect 700 1838 734 1872
rect 768 1838 802 1872
rect 836 1838 870 1872
rect 904 1838 938 1872
rect 972 1838 1006 1872
rect -98 1733 -64 1767
rect -98 1665 -64 1699
rect 1090 1733 1124 1767
rect -98 1597 -64 1631
rect 1090 1665 1124 1699
rect -98 1529 -64 1563
rect 1090 1597 1124 1631
rect 1090 1529 1124 1563
rect 20 1424 54 1458
rect 88 1424 122 1458
rect 156 1424 190 1458
rect 224 1424 258 1458
rect 292 1424 326 1458
rect 360 1424 394 1458
rect 428 1424 462 1458
rect 496 1424 530 1458
rect 564 1424 598 1458
rect 632 1424 666 1458
rect 700 1424 734 1458
rect 768 1424 802 1458
rect 836 1424 870 1458
rect 904 1424 938 1458
rect 972 1424 1006 1458
rect 1314 1838 1348 1872
rect 1382 1838 1416 1872
rect 1450 1838 1484 1872
rect 1518 1838 1552 1872
rect 1586 1838 1620 1872
rect 1654 1838 1688 1872
rect 1722 1838 1756 1872
rect 1790 1838 1824 1872
rect 1858 1838 1892 1872
rect 1926 1838 1960 1872
rect 1994 1838 2028 1872
rect 2062 1838 2096 1872
rect 2130 1838 2164 1872
rect 2198 1838 2232 1872
rect 2266 1838 2300 1872
rect 1196 1733 1230 1767
rect 1196 1665 1230 1699
rect 2384 1733 2418 1767
rect 1196 1597 1230 1631
rect 2384 1665 2418 1699
rect 1196 1529 1230 1563
rect 2384 1597 2418 1631
rect 2384 1529 2418 1563
rect 1314 1424 1348 1458
rect 1382 1424 1416 1458
rect 1450 1424 1484 1458
rect 1518 1424 1552 1458
rect 1586 1424 1620 1458
rect 1654 1424 1688 1458
rect 1722 1424 1756 1458
rect 1790 1424 1824 1458
rect 1858 1424 1892 1458
rect 1926 1424 1960 1458
rect 1994 1424 2028 1458
rect 2062 1424 2096 1458
rect 2130 1424 2164 1458
rect 2198 1424 2232 1458
rect 2266 1424 2300 1458
rect 1310 806 1344 840
rect 1378 806 1412 840
rect 1446 806 1480 840
rect 1514 806 1548 840
rect 1582 806 1616 840
rect 1650 806 1684 840
rect 1718 806 1752 840
rect 1786 806 1820 840
rect 1854 806 1888 840
rect 1922 806 1956 840
rect 1990 806 2024 840
rect 2058 806 2092 840
rect 2126 806 2160 840
rect 2194 806 2228 840
rect 2262 806 2296 840
rect 1192 701 1226 735
rect 1192 633 1226 667
rect 2380 701 2414 735
rect 1192 565 1226 599
rect 2380 633 2414 667
rect 1192 497 1226 531
rect 2380 565 2414 599
rect 2380 497 2414 531
rect 1310 392 1344 426
rect 1378 392 1412 426
rect 1446 392 1480 426
rect 1514 392 1548 426
rect 1582 392 1616 426
rect 1650 392 1684 426
rect 1718 392 1752 426
rect 1786 392 1820 426
rect 1854 392 1888 426
rect 1922 392 1956 426
rect 1990 392 2024 426
rect 2058 392 2092 426
rect 2126 392 2160 426
rect 2194 392 2228 426
rect 2262 392 2296 426
<< nsubdiffcont >>
rect -1195 6540 -1161 6574
rect -1127 6540 -1093 6574
rect -1059 6540 -1025 6574
rect -991 6540 -957 6574
rect -923 6540 -889 6574
rect -855 6540 -821 6574
rect -787 6540 -753 6574
rect -719 6540 -685 6574
rect -651 6540 -617 6574
rect -583 6540 -549 6574
rect -515 6540 -481 6574
rect -447 6540 -413 6574
rect -379 6540 -345 6574
rect -311 6540 -277 6574
rect -243 6540 -209 6574
rect -175 6540 -141 6574
rect -107 6540 -73 6574
rect -39 6540 -5 6574
rect 29 6540 63 6574
rect 97 6540 131 6574
rect 165 6540 199 6574
rect 233 6540 267 6574
rect 301 6540 335 6574
rect 369 6540 403 6574
rect 437 6540 471 6574
rect 505 6540 539 6574
rect 573 6540 607 6574
rect 641 6540 675 6574
rect 709 6540 743 6574
rect 777 6540 811 6574
rect 845 6540 879 6574
rect 913 6540 947 6574
rect 981 6540 1015 6574
rect 1049 6540 1083 6574
rect 1117 6540 1151 6574
rect -1298 6424 -1264 6458
rect 1220 6424 1254 6458
rect -1298 6356 -1264 6390
rect -1298 6288 -1264 6322
rect -1298 6220 -1264 6254
rect -1298 6152 -1264 6186
rect -1298 6084 -1264 6118
rect -1298 6016 -1264 6050
rect -1298 5948 -1264 5982
rect -1298 5880 -1264 5914
rect -1298 5812 -1264 5846
rect -1298 5744 -1264 5778
rect -1298 5676 -1264 5710
rect -1298 5608 -1264 5642
rect -1298 5540 -1264 5574
rect -1298 5472 -1264 5506
rect -1298 5404 -1264 5438
rect -1298 5336 -1264 5370
rect -1298 5268 -1264 5302
rect -1298 5200 -1264 5234
rect -1298 5132 -1264 5166
rect -1298 5064 -1264 5098
rect -1298 4996 -1264 5030
rect -1298 4928 -1264 4962
rect -1298 4860 -1264 4894
rect -1298 4792 -1264 4826
rect 1220 6356 1254 6390
rect 1220 6288 1254 6322
rect 1220 6220 1254 6254
rect 1220 6152 1254 6186
rect 1220 6084 1254 6118
rect 1220 6016 1254 6050
rect 1220 5948 1254 5982
rect 1220 5880 1254 5914
rect 1220 5812 1254 5846
rect 1220 5744 1254 5778
rect 1220 5676 1254 5710
rect 1220 5608 1254 5642
rect 1220 5540 1254 5574
rect 1220 5472 1254 5506
rect 1220 5404 1254 5438
rect 1220 5336 1254 5370
rect 1220 5268 1254 5302
rect 1220 5200 1254 5234
rect 1220 5132 1254 5166
rect 1220 5064 1254 5098
rect 1220 4996 1254 5030
rect 1220 4928 1254 4962
rect 1220 4860 1254 4894
rect 1220 4792 1254 4826
rect -1298 4724 -1264 4758
rect 1220 4724 1254 4758
rect -1195 4608 -1161 4642
rect -1127 4608 -1093 4642
rect -1059 4608 -1025 4642
rect -991 4608 -957 4642
rect -923 4608 -889 4642
rect -855 4608 -821 4642
rect -787 4608 -753 4642
rect -719 4608 -685 4642
rect -651 4608 -617 4642
rect -583 4608 -549 4642
rect -515 4608 -481 4642
rect -447 4608 -413 4642
rect -379 4608 -345 4642
rect -311 4608 -277 4642
rect -243 4608 -209 4642
rect -175 4608 -141 4642
rect -107 4608 -73 4642
rect -39 4608 -5 4642
rect 29 4608 63 4642
rect 97 4608 131 4642
rect 165 4608 199 4642
rect 233 4608 267 4642
rect 301 4608 335 4642
rect 369 4608 403 4642
rect 437 4608 471 4642
rect 505 4608 539 4642
rect 573 4608 607 4642
rect 641 4608 675 4642
rect 709 4608 743 4642
rect 777 4608 811 4642
rect 845 4608 879 4642
rect 913 4608 947 4642
rect 981 4608 1015 4642
rect 1049 4608 1083 4642
rect 1117 4608 1151 4642
rect -1195 4502 -1161 4536
rect -1127 4502 -1093 4536
rect -1059 4502 -1025 4536
rect -991 4502 -957 4536
rect -923 4502 -889 4536
rect -855 4502 -821 4536
rect -787 4502 -753 4536
rect -719 4502 -685 4536
rect -651 4502 -617 4536
rect -583 4502 -549 4536
rect -515 4502 -481 4536
rect -447 4502 -413 4536
rect -379 4502 -345 4536
rect -311 4502 -277 4536
rect -243 4502 -209 4536
rect -175 4502 -141 4536
rect -107 4502 -73 4536
rect -39 4502 -5 4536
rect 29 4502 63 4536
rect 97 4502 131 4536
rect 165 4502 199 4536
rect 233 4502 267 4536
rect 301 4502 335 4536
rect 369 4502 403 4536
rect 437 4502 471 4536
rect 505 4502 539 4536
rect 573 4502 607 4536
rect 641 4502 675 4536
rect 709 4502 743 4536
rect 777 4502 811 4536
rect 845 4502 879 4536
rect 913 4502 947 4536
rect 981 4502 1015 4536
rect 1049 4502 1083 4536
rect 1117 4502 1151 4536
rect -1298 4386 -1264 4420
rect 1220 4386 1254 4420
rect -1298 4318 -1264 4352
rect -1298 4250 -1264 4284
rect -1298 4182 -1264 4216
rect -1298 4114 -1264 4148
rect -1298 4046 -1264 4080
rect -1298 3978 -1264 4012
rect -1298 3910 -1264 3944
rect -1298 3842 -1264 3876
rect -1298 3774 -1264 3808
rect -1298 3706 -1264 3740
rect -1298 3638 -1264 3672
rect -1298 3570 -1264 3604
rect -1298 3502 -1264 3536
rect -1298 3434 -1264 3468
rect -1298 3366 -1264 3400
rect -1298 3298 -1264 3332
rect -1298 3230 -1264 3264
rect -1298 3162 -1264 3196
rect -1298 3094 -1264 3128
rect -1298 3026 -1264 3060
rect -1298 2958 -1264 2992
rect -1298 2890 -1264 2924
rect -1298 2822 -1264 2856
rect -1298 2754 -1264 2788
rect 1220 4318 1254 4352
rect 1220 4250 1254 4284
rect 1220 4182 1254 4216
rect 1220 4114 1254 4148
rect 1220 4046 1254 4080
rect 1220 3978 1254 4012
rect 1220 3910 1254 3944
rect 1220 3842 1254 3876
rect 1220 3774 1254 3808
rect 1220 3706 1254 3740
rect 1220 3638 1254 3672
rect 1220 3570 1254 3604
rect 1220 3502 1254 3536
rect 1220 3434 1254 3468
rect 1220 3366 1254 3400
rect 1220 3298 1254 3332
rect 1220 3230 1254 3264
rect 1220 3162 1254 3196
rect 1220 3094 1254 3128
rect 1220 3026 1254 3060
rect 1220 2958 1254 2992
rect 1220 2890 1254 2924
rect 1220 2822 1254 2856
rect 1220 2754 1254 2788
rect -1298 2686 -1264 2720
rect 1220 2686 1254 2720
rect -1195 2570 -1161 2604
rect -1127 2570 -1093 2604
rect -1059 2570 -1025 2604
rect -991 2570 -957 2604
rect -923 2570 -889 2604
rect -855 2570 -821 2604
rect -787 2570 -753 2604
rect -719 2570 -685 2604
rect -651 2570 -617 2604
rect -583 2570 -549 2604
rect -515 2570 -481 2604
rect -447 2570 -413 2604
rect -379 2570 -345 2604
rect -311 2570 -277 2604
rect -243 2570 -209 2604
rect -175 2570 -141 2604
rect -107 2570 -73 2604
rect -39 2570 -5 2604
rect 29 2570 63 2604
rect 97 2570 131 2604
rect 165 2570 199 2604
rect 233 2570 267 2604
rect 301 2570 335 2604
rect 369 2570 403 2604
rect 437 2570 471 2604
rect 505 2570 539 2604
rect 573 2570 607 2604
rect 641 2570 675 2604
rect 709 2570 743 2604
rect 777 2570 811 2604
rect 845 2570 879 2604
rect 913 2570 947 2604
rect 981 2570 1015 2604
rect 1049 2570 1083 2604
rect 1117 2570 1151 2604
<< poly >>
rect 48 1770 114 1786
rect 48 1736 64 1770
rect 98 1736 114 1770
rect 48 1720 114 1736
rect 240 1770 306 1786
rect 240 1736 256 1770
rect 290 1736 306 1770
rect 66 1698 96 1720
rect 162 1698 192 1724
rect 240 1720 306 1736
rect 432 1770 498 1786
rect 432 1736 448 1770
rect 482 1736 498 1770
rect 258 1698 288 1720
rect 354 1698 384 1724
rect 432 1720 498 1736
rect 624 1770 690 1786
rect 624 1736 640 1770
rect 674 1736 690 1770
rect 450 1698 480 1720
rect 546 1698 576 1724
rect 624 1720 690 1736
rect 816 1770 960 1786
rect 816 1736 832 1770
rect 866 1736 960 1770
rect 642 1698 672 1720
rect 738 1698 768 1724
rect 816 1720 960 1736
rect 834 1698 864 1720
rect 930 1698 960 1720
rect 66 1576 96 1598
rect 162 1576 192 1598
rect 66 1560 210 1576
rect 258 1572 288 1598
rect 354 1576 384 1598
rect 66 1526 160 1560
rect 194 1526 210 1560
rect 66 1510 210 1526
rect 336 1560 402 1576
rect 450 1572 480 1598
rect 546 1576 576 1598
rect 336 1526 352 1560
rect 386 1526 402 1560
rect 336 1510 402 1526
rect 528 1560 594 1576
rect 642 1572 672 1598
rect 738 1576 768 1598
rect 528 1526 544 1560
rect 578 1526 594 1560
rect 528 1510 594 1526
rect 720 1560 786 1576
rect 834 1572 864 1598
rect 930 1576 960 1598
rect 720 1526 736 1560
rect 770 1526 786 1560
rect 720 1510 786 1526
rect 912 1560 978 1576
rect 912 1526 928 1560
rect 962 1526 978 1560
rect 912 1510 978 1526
rect 1342 1770 1408 1786
rect 1342 1736 1358 1770
rect 1392 1736 1408 1770
rect 1342 1720 1408 1736
rect 1534 1770 1600 1786
rect 1534 1736 1550 1770
rect 1584 1736 1600 1770
rect 1360 1698 1390 1720
rect 1456 1698 1486 1724
rect 1534 1720 1600 1736
rect 1726 1770 1792 1786
rect 1726 1736 1742 1770
rect 1776 1736 1792 1770
rect 1552 1698 1582 1720
rect 1648 1698 1678 1724
rect 1726 1720 1792 1736
rect 1918 1770 1984 1786
rect 1918 1736 1934 1770
rect 1968 1736 1984 1770
rect 1744 1698 1774 1720
rect 1840 1698 1870 1724
rect 1918 1720 1984 1736
rect 2110 1770 2254 1786
rect 2110 1736 2126 1770
rect 2160 1736 2254 1770
rect 1936 1698 1966 1720
rect 2032 1698 2062 1724
rect 2110 1720 2254 1736
rect 2128 1698 2158 1720
rect 2224 1698 2254 1720
rect 1360 1576 1390 1598
rect 1456 1576 1486 1598
rect 1360 1560 1504 1576
rect 1552 1572 1582 1598
rect 1648 1576 1678 1598
rect 1360 1526 1454 1560
rect 1488 1526 1504 1560
rect 1360 1510 1504 1526
rect 1630 1560 1696 1576
rect 1744 1572 1774 1598
rect 1840 1576 1870 1598
rect 1630 1526 1646 1560
rect 1680 1526 1696 1560
rect 1630 1510 1696 1526
rect 1822 1560 1888 1576
rect 1936 1572 1966 1598
rect 2032 1576 2062 1598
rect 1822 1526 1838 1560
rect 1872 1526 1888 1560
rect 1822 1510 1888 1526
rect 2014 1560 2080 1576
rect 2128 1572 2158 1598
rect 2224 1576 2254 1598
rect 2014 1526 2030 1560
rect 2064 1526 2080 1560
rect 2014 1510 2080 1526
rect 2206 1560 2272 1576
rect 2206 1526 2222 1560
rect 2256 1526 2272 1560
rect 2206 1510 2272 1526
rect 62 688 140 754
rect 1356 738 1500 754
rect 1356 704 1450 738
rect 1484 704 1500 738
rect 1356 688 1500 704
rect 1626 738 1692 754
rect 1626 704 1642 738
rect 1676 704 1692 738
rect 1356 666 1386 688
rect 1452 666 1482 688
rect 1548 666 1578 692
rect 1626 688 1692 704
rect 1818 738 1884 754
rect 1818 704 1834 738
rect 1868 704 1884 738
rect 1644 666 1674 688
rect 1740 666 1770 692
rect 1818 688 1884 704
rect 2010 738 2076 754
rect 2010 704 2026 738
rect 2060 704 2076 738
rect 1836 666 1866 688
rect 1932 666 1962 692
rect 2010 688 2076 704
rect 2202 738 2268 754
rect 2202 704 2218 738
rect 2252 704 2268 738
rect 2028 666 2058 688
rect 2124 666 2154 692
rect 2202 688 2268 704
rect 2220 666 2250 688
rect 878 478 956 544
rect 1356 544 1386 566
rect 1338 528 1404 544
rect 1452 540 1482 566
rect 1548 544 1578 566
rect 1338 494 1354 528
rect 1388 494 1404 528
rect 1338 478 1404 494
rect 1530 528 1596 544
rect 1644 540 1674 566
rect 1740 544 1770 566
rect 1530 494 1546 528
rect 1580 494 1596 528
rect 1530 478 1596 494
rect 1722 528 1788 544
rect 1836 540 1866 566
rect 1932 544 1962 566
rect 1722 494 1738 528
rect 1772 494 1788 528
rect 1722 478 1788 494
rect 1914 528 1980 544
rect 2028 540 2058 566
rect 2124 544 2154 566
rect 2220 544 2250 566
rect 1914 494 1930 528
rect 1964 494 1980 528
rect 1914 478 1980 494
rect 2106 528 2250 544
rect 2106 494 2122 528
rect 2156 494 2250 528
rect 2106 478 2250 494
<< polycont >>
rect 64 1736 98 1770
rect 256 1736 290 1770
rect 448 1736 482 1770
rect 640 1736 674 1770
rect 832 1736 866 1770
rect 160 1526 194 1560
rect 352 1526 386 1560
rect 544 1526 578 1560
rect 736 1526 770 1560
rect 928 1526 962 1560
rect 1358 1736 1392 1770
rect 1550 1736 1584 1770
rect 1742 1736 1776 1770
rect 1934 1736 1968 1770
rect 2126 1736 2160 1770
rect 1454 1526 1488 1560
rect 1646 1526 1680 1560
rect 1838 1526 1872 1560
rect 2030 1526 2064 1560
rect 2222 1526 2256 1560
rect 1450 704 1484 738
rect 1642 704 1676 738
rect 1834 704 1868 738
rect 2026 704 2060 738
rect 2218 704 2252 738
rect 1354 494 1388 528
rect 1546 494 1580 528
rect 1738 494 1772 528
rect 1930 494 1964 528
rect 2122 494 2156 528
<< locali >>
rect -1298 6540 -1195 6574
rect -1157 6540 -1127 6574
rect -1085 6540 -1059 6574
rect -1013 6540 -991 6574
rect -941 6540 -923 6574
rect -869 6540 -855 6574
rect -797 6540 -787 6574
rect -725 6540 -719 6574
rect -653 6540 -651 6574
rect -617 6540 -615 6574
rect -549 6540 -543 6574
rect -481 6540 -471 6574
rect -413 6540 -399 6574
rect -345 6540 -327 6574
rect -277 6540 -255 6574
rect -209 6540 -183 6574
rect -141 6540 -111 6574
rect -73 6540 -39 6574
rect -5 6540 29 6574
rect 67 6540 97 6574
rect 139 6540 165 6574
rect 211 6540 233 6574
rect 283 6540 301 6574
rect 355 6540 369 6574
rect 427 6540 437 6574
rect 499 6540 505 6574
rect 571 6540 573 6574
rect 607 6540 609 6574
rect 675 6540 681 6574
rect 743 6540 753 6574
rect 811 6540 825 6574
rect 879 6540 897 6574
rect 947 6540 969 6574
rect 1015 6540 1041 6574
rect 1083 6540 1113 6574
rect 1151 6540 1254 6574
rect 1422 6540 1433 6574
rect 1467 6540 1505 6574
rect 1539 6540 1577 6574
rect 1611 6540 1649 6574
rect 1683 6540 1721 6574
rect 1755 6540 1793 6574
rect 1827 6540 1865 6574
rect 1899 6540 1937 6574
rect 1971 6540 2009 6574
rect 2043 6540 2081 6574
rect 2115 6540 2153 6574
rect 2187 6540 2225 6574
rect 2259 6540 2297 6574
rect 2331 6540 2369 6574
rect 2403 6540 2441 6574
rect 2475 6540 2513 6574
rect 2547 6540 2585 6574
rect 2619 6540 2657 6574
rect 2691 6540 2729 6574
rect 2763 6540 2801 6574
rect 2835 6540 2873 6574
rect 2907 6540 2945 6574
rect 2979 6540 3017 6574
rect 3051 6540 3089 6574
rect 3123 6540 3161 6574
rect 3195 6540 3233 6574
rect 3267 6540 3305 6574
rect 3339 6540 3377 6574
rect 3411 6540 3449 6574
rect 3483 6540 3521 6574
rect 3555 6540 3593 6574
rect 3627 6540 3665 6574
rect 3699 6540 3737 6574
rect 3771 6540 3782 6574
rect -1298 6458 -1264 6540
rect 1220 6472 1254 6540
rect -982 6438 -726 6472
rect -692 6438 190 6472
rect 224 6438 916 6472
rect 946 6438 1106 6472
rect 1140 6438 1156 6472
rect -1298 6390 -1264 6424
rect 1220 6400 1254 6424
rect -1298 6322 -1264 6356
rect -1298 6254 -1264 6288
rect -1298 6186 -1264 6220
rect -1298 6118 -1264 6152
rect -1298 6050 -1264 6084
rect -1298 5982 -1264 6016
rect -1298 5914 -1264 5948
rect -1298 5846 -1264 5880
rect -1298 5778 -1264 5812
rect -1298 5710 -1264 5744
rect -1298 5642 -1264 5676
rect -1298 5574 -1264 5608
rect -1298 5506 -1264 5540
rect -1298 5438 -1264 5472
rect -1298 5370 -1264 5404
rect -1298 5302 -1264 5336
rect -1298 5234 -1264 5268
rect -1298 5166 -1264 5200
rect -1298 5098 -1264 5132
rect -1298 5030 -1264 5064
rect -1298 4962 -1264 4996
rect -1298 4894 -1264 4928
rect -1298 4826 -1264 4860
rect -1298 4758 -1264 4792
rect -1184 6364 -1150 6395
rect -1184 6292 -1150 6330
rect -1184 6220 -1150 6258
rect -1184 6148 -1150 6186
rect -1184 6076 -1150 6114
rect -1184 6004 -1150 6042
rect -1184 5932 -1150 5970
rect -1184 5860 -1150 5898
rect -1184 5788 -1150 5826
rect -1184 5716 -1150 5754
rect -1184 5644 -1150 5682
rect -1184 5572 -1150 5610
rect -1184 5500 -1150 5538
rect -1184 5428 -1150 5466
rect -1184 5356 -1150 5394
rect -1184 5284 -1150 5322
rect -1184 5212 -1150 5250
rect -1184 5140 -1150 5178
rect -1184 5068 -1150 5106
rect -1184 4996 -1150 5034
rect -1184 4924 -1150 4962
rect -1184 4852 -1150 4890
rect -1184 4787 -1150 4818
rect -726 6364 -692 6395
rect -726 6292 -692 6330
rect -726 6220 -692 6258
rect -726 6148 -692 6186
rect -726 6076 -692 6114
rect -726 6004 -692 6042
rect -726 5932 -692 5970
rect -726 5860 -692 5898
rect -726 5788 -692 5826
rect -726 5716 -692 5754
rect -726 5644 -692 5682
rect -726 5572 -692 5610
rect -726 5500 -692 5538
rect -726 5428 -692 5466
rect -726 5356 -692 5394
rect -726 5284 -692 5322
rect -726 5212 -692 5250
rect -726 5140 -692 5178
rect -726 5068 -692 5106
rect -726 4996 -692 5034
rect -726 4924 -692 4962
rect -726 4852 -692 4890
rect -726 4787 -692 4818
rect -268 6364 -234 6395
rect -268 6292 -234 6330
rect -268 6220 -234 6258
rect -268 6148 -234 6186
rect -268 6076 -234 6114
rect -268 6004 -234 6042
rect -268 5932 -234 5970
rect -268 5860 -234 5898
rect -268 5788 -234 5826
rect -268 5716 -234 5754
rect -268 5644 -234 5682
rect -268 5572 -234 5610
rect -268 5500 -234 5538
rect -268 5428 -234 5466
rect -268 5356 -234 5394
rect -268 5284 -234 5322
rect -268 5212 -234 5250
rect -268 5140 -234 5178
rect -268 5068 -234 5106
rect -268 4996 -234 5034
rect -268 4924 -234 4962
rect -268 4852 -234 4890
rect -268 4787 -234 4818
rect 190 6364 224 6395
rect 190 6292 224 6330
rect 190 6220 224 6258
rect 190 6148 224 6186
rect 190 6076 224 6114
rect 190 6004 224 6042
rect 190 5932 224 5970
rect 190 5860 224 5898
rect 190 5788 224 5826
rect 190 5716 224 5754
rect 190 5644 224 5682
rect 190 5572 224 5610
rect 190 5500 224 5538
rect 190 5428 224 5466
rect 190 5356 224 5394
rect 190 5284 224 5322
rect 190 5212 224 5250
rect 190 5140 224 5178
rect 190 5068 224 5106
rect 190 4996 224 5034
rect 190 4924 224 4962
rect 190 4852 224 4890
rect 190 4787 224 4818
rect 648 6364 682 6395
rect 648 6292 682 6330
rect 648 6220 682 6258
rect 648 6148 682 6186
rect 648 6076 682 6114
rect 648 6004 682 6042
rect 648 5932 682 5970
rect 648 5860 682 5898
rect 648 5788 682 5826
rect 648 5716 682 5754
rect 648 5644 682 5682
rect 648 5572 682 5610
rect 648 5500 682 5538
rect 648 5428 682 5466
rect 648 5356 682 5394
rect 648 5284 682 5322
rect 648 5212 682 5250
rect 648 5140 682 5178
rect 648 5068 682 5106
rect 648 4996 682 5034
rect 648 4924 682 4962
rect 648 4852 682 4890
rect 648 4787 682 4818
rect 1106 6364 1140 6395
rect 1106 6292 1140 6330
rect 1106 6220 1140 6258
rect 1106 6148 1140 6186
rect 1106 6076 1140 6114
rect 1106 6004 1140 6042
rect 1106 5932 1140 5970
rect 1106 5860 1140 5898
rect 1106 5788 1140 5826
rect 1106 5716 1140 5754
rect 1106 5644 1140 5682
rect 1106 5572 1140 5610
rect 1106 5500 1140 5538
rect 1106 5428 1140 5466
rect 1106 5356 1140 5394
rect 1106 5284 1140 5322
rect 1106 5212 1140 5250
rect 1106 5140 1140 5178
rect 1106 5068 1140 5106
rect 1106 4996 1140 5034
rect 1106 4924 1140 4962
rect 1106 4852 1140 4890
rect 1106 4787 1140 4818
rect 1220 6328 1254 6356
rect 1220 6256 1254 6288
rect 1220 6186 1254 6220
rect 1220 6118 1254 6150
rect 1220 6050 1254 6078
rect 1220 5982 1254 6006
rect 1220 5914 1254 5934
rect 1220 5846 1254 5862
rect 1220 5778 1254 5790
rect 1220 5710 1254 5718
rect 1220 5642 1254 5646
rect 1220 5536 1254 5540
rect 1220 5464 1254 5472
rect 1220 5392 1254 5404
rect 1220 5320 1254 5336
rect 1220 5248 1254 5268
rect 1220 5176 1254 5200
rect 1220 5104 1254 5132
rect 1220 5032 1254 5064
rect 1220 4962 1254 4996
rect 1220 4894 1254 4926
rect 1220 4826 1254 4854
rect 1220 4758 1254 4782
rect -1298 4642 -1264 4724
rect -980 4710 -726 4744
rect -692 4710 190 4744
rect 224 4710 918 4744
rect 946 4710 1106 4744
rect 1140 4710 1156 4744
rect 1220 4642 1254 4710
rect 1326 6472 1360 6478
rect 1424 6438 1440 6472
rect 1474 6438 1634 6472
rect 1640 6438 2356 6472
rect 2390 6438 3272 6472
rect 3306 6438 3544 6472
rect 1326 6400 1360 6438
rect 1326 6328 1360 6366
rect 1326 6256 1360 6294
rect 1326 6184 1360 6222
rect 1326 6112 1360 6150
rect 1326 6040 1360 6078
rect 1326 5968 1360 6006
rect 1326 5896 1360 5934
rect 1326 5824 1360 5862
rect 1326 5752 1360 5790
rect 1326 5680 1360 5718
rect 1326 5608 1360 5646
rect 1326 5536 1360 5574
rect 1326 5464 1360 5502
rect 1326 5392 1360 5430
rect 1326 5320 1360 5358
rect 1326 5248 1360 5286
rect 1326 5176 1360 5214
rect 1326 5104 1360 5142
rect 1326 5032 1360 5070
rect 1326 4960 1360 4998
rect 1326 4888 1360 4926
rect 1326 4816 1360 4854
rect 1326 4744 1360 4782
rect 1424 4710 1440 4744
rect 1474 4710 1634 4744
rect 1656 4710 2356 4744
rect 2390 4710 3272 4744
rect 3306 4710 3560 4744
rect 1326 4704 1360 4710
rect -1298 4608 -1263 4642
rect -1229 4608 -1195 4642
rect -1157 4608 -1127 4642
rect -1085 4608 -1059 4642
rect -1013 4608 -991 4642
rect -941 4608 -923 4642
rect -869 4608 -855 4642
rect -797 4608 -787 4642
rect -725 4608 -719 4642
rect -653 4608 -651 4642
rect -617 4608 -615 4642
rect -549 4608 -543 4642
rect -481 4608 -471 4642
rect -413 4608 -399 4642
rect -345 4608 -327 4642
rect -277 4608 -255 4642
rect -209 4608 -183 4642
rect -141 4608 -111 4642
rect -73 4608 -39 4642
rect -5 4608 29 4642
rect 67 4608 97 4642
rect 139 4608 165 4642
rect 211 4608 233 4642
rect 283 4608 301 4642
rect 355 4608 369 4642
rect 427 4608 437 4642
rect 499 4608 505 4642
rect 571 4608 573 4642
rect 607 4608 609 4642
rect 675 4608 681 4642
rect 743 4608 753 4642
rect 811 4608 825 4642
rect 879 4608 897 4642
rect 947 4608 969 4642
rect 1015 4608 1041 4642
rect 1083 4608 1113 4642
rect 1151 4608 1185 4642
rect 1219 4608 1254 4642
rect -1298 4502 -1263 4536
rect -1229 4502 -1195 4536
rect -1157 4502 -1127 4536
rect -1085 4502 -1059 4536
rect -1013 4502 -991 4536
rect -941 4502 -923 4536
rect -869 4502 -855 4536
rect -797 4502 -787 4536
rect -725 4502 -719 4536
rect -653 4502 -651 4536
rect -617 4502 -615 4536
rect -549 4502 -543 4536
rect -481 4502 -471 4536
rect -413 4502 -399 4536
rect -345 4502 -327 4536
rect -277 4502 -255 4536
rect -209 4502 -183 4536
rect -141 4502 -111 4536
rect -73 4502 -39 4536
rect -5 4502 29 4536
rect 67 4502 97 4536
rect 139 4502 165 4536
rect 211 4502 233 4536
rect 283 4502 301 4536
rect 355 4502 369 4536
rect 427 4502 437 4536
rect 499 4502 505 4536
rect 571 4502 573 4536
rect 607 4502 609 4536
rect 675 4502 681 4536
rect 743 4502 753 4536
rect 811 4502 825 4536
rect 879 4502 897 4536
rect 947 4502 969 4536
rect 1015 4502 1041 4536
rect 1083 4502 1113 4536
rect 1151 4502 1185 4536
rect 1219 4502 1254 4536
rect -1298 4420 -1264 4502
rect 1220 4434 1254 4502
rect -978 4400 920 4434
rect -1298 4352 -1264 4386
rect 1220 4362 1254 4386
rect -1298 4284 -1264 4318
rect -1298 4216 -1264 4250
rect -1298 4148 -1264 4182
rect -1298 4080 -1264 4114
rect -1298 4012 -1264 4046
rect -1298 3944 -1264 3978
rect -1298 3876 -1264 3910
rect -1298 3808 -1264 3842
rect -1298 3740 -1264 3774
rect -1298 3672 -1264 3706
rect -1298 3604 -1264 3638
rect -1298 3536 -1264 3570
rect -1298 3468 -1264 3502
rect -1298 3400 -1264 3434
rect -1298 3332 -1264 3366
rect -1298 3264 -1264 3298
rect -1298 3196 -1264 3230
rect -1298 3128 -1264 3162
rect -1298 3060 -1264 3094
rect -1298 2992 -1264 3026
rect -1298 2924 -1264 2958
rect -1298 2856 -1264 2890
rect -1298 2788 -1264 2822
rect -1298 2720 -1264 2754
rect -1184 4326 -1150 4357
rect -1184 4254 -1150 4292
rect -1184 4182 -1150 4220
rect -1184 4110 -1150 4148
rect -1184 4038 -1150 4076
rect -1184 3966 -1150 4004
rect -1184 3894 -1150 3932
rect -1184 3822 -1150 3860
rect -1184 3750 -1150 3788
rect -1184 3678 -1150 3716
rect -1184 3606 -1150 3644
rect -1184 3534 -1150 3572
rect -1184 3462 -1150 3500
rect -1184 3390 -1150 3428
rect -1184 3318 -1150 3356
rect -1184 3246 -1150 3284
rect -1184 3174 -1150 3212
rect -1184 3102 -1150 3140
rect -1184 3030 -1150 3068
rect -1184 2958 -1150 2996
rect -1184 2886 -1150 2924
rect -1184 2814 -1150 2852
rect -1184 2749 -1150 2780
rect -726 4326 -692 4357
rect -726 4254 -692 4292
rect -726 4182 -692 4220
rect -726 4110 -692 4148
rect -726 4038 -692 4076
rect -726 3966 -692 4004
rect -726 3894 -692 3932
rect -726 3822 -692 3860
rect -726 3750 -692 3788
rect -726 3678 -692 3716
rect -726 3606 -692 3644
rect -726 3534 -692 3572
rect -726 3462 -692 3500
rect -726 3390 -692 3428
rect -726 3318 -692 3356
rect -726 3246 -692 3284
rect -726 3174 -692 3212
rect -726 3102 -692 3140
rect -726 3030 -692 3068
rect -726 2958 -692 2996
rect -726 2886 -692 2924
rect -726 2814 -692 2852
rect -726 2749 -692 2780
rect -268 4326 -234 4357
rect -268 4254 -234 4292
rect -268 4182 -234 4220
rect -268 4110 -234 4148
rect -268 4038 -234 4076
rect -268 3966 -234 4004
rect -268 3894 -234 3932
rect -268 3822 -234 3860
rect -268 3750 -234 3788
rect -268 3678 -234 3716
rect -268 3606 -234 3644
rect -268 3534 -234 3572
rect -268 3462 -234 3500
rect -268 3390 -234 3428
rect -268 3318 -234 3356
rect -268 3246 -234 3284
rect -268 3174 -234 3212
rect -268 3102 -234 3140
rect -268 3030 -234 3068
rect -268 2958 -234 2996
rect -268 2886 -234 2924
rect -268 2814 -234 2852
rect -268 2749 -234 2780
rect 190 4326 224 4357
rect 190 4254 224 4292
rect 190 4182 224 4220
rect 190 4110 224 4148
rect 190 4038 224 4076
rect 190 3966 224 4004
rect 190 3894 224 3932
rect 190 3822 224 3860
rect 190 3750 224 3788
rect 190 3678 224 3716
rect 190 3606 224 3644
rect 190 3534 224 3572
rect 190 3462 224 3500
rect 190 3390 224 3428
rect 190 3318 224 3356
rect 190 3246 224 3284
rect 190 3174 224 3212
rect 190 3102 224 3140
rect 190 3030 224 3068
rect 190 2958 224 2996
rect 190 2886 224 2924
rect 190 2814 224 2852
rect 190 2749 224 2780
rect 648 4326 682 4357
rect 648 4254 682 4292
rect 648 4182 682 4220
rect 648 4110 682 4148
rect 648 4038 682 4076
rect 648 3966 682 4004
rect 648 3894 682 3932
rect 648 3822 682 3860
rect 648 3750 682 3788
rect 648 3678 682 3716
rect 648 3606 682 3644
rect 648 3534 682 3572
rect 648 3462 682 3500
rect 648 3390 682 3428
rect 648 3318 682 3356
rect 648 3246 682 3284
rect 648 3174 682 3212
rect 648 3102 682 3140
rect 648 3030 682 3068
rect 648 2958 682 2996
rect 648 2886 682 2924
rect 648 2814 682 2852
rect 648 2749 682 2780
rect 1106 4326 1140 4357
rect 1106 4254 1140 4292
rect 1106 4182 1140 4220
rect 1106 4110 1140 4148
rect 1106 4038 1140 4076
rect 1106 3966 1140 4004
rect 1106 3894 1140 3932
rect 1106 3822 1140 3860
rect 1106 3750 1140 3788
rect 1106 3678 1140 3716
rect 1106 3606 1140 3644
rect 1106 3534 1140 3572
rect 1106 3462 1140 3500
rect 1106 3390 1140 3428
rect 1106 3318 1140 3356
rect 1106 3246 1140 3284
rect 1106 3174 1140 3212
rect 1106 3102 1140 3140
rect 1106 3030 1140 3068
rect 1106 2958 1140 2996
rect 1106 2886 1140 2924
rect 1106 2814 1140 2852
rect 1106 2749 1140 2780
rect 1220 4290 1254 4318
rect 1220 4218 1254 4250
rect 1220 4148 1254 4182
rect 1220 4080 1254 4112
rect 1220 4012 1254 4040
rect 1220 3944 1254 3968
rect 1220 3876 1254 3896
rect 1220 3808 1254 3824
rect 1220 3740 1254 3752
rect 1220 3672 1254 3680
rect 1220 3604 1254 3608
rect 1220 3498 1254 3502
rect 1220 3426 1254 3434
rect 1220 3354 1254 3366
rect 1220 3282 1254 3298
rect 1220 3210 1254 3230
rect 1220 3138 1254 3162
rect 1220 3066 1254 3094
rect 1220 2994 1254 3026
rect 1220 2924 1254 2958
rect 1220 2856 1254 2888
rect 1220 2788 1254 2816
rect 1220 2720 1254 2744
rect -1298 2604 -1264 2686
rect -982 2672 860 2706
rect 894 2672 916 2706
rect 1220 2604 1254 2672
rect 1326 4434 1360 4440
rect 1680 4400 3560 4434
rect 1326 4362 1360 4400
rect 1326 4290 1360 4328
rect 1326 4218 1360 4256
rect 1326 4146 1360 4184
rect 1326 4074 1360 4112
rect 1326 4002 1360 4040
rect 1326 3930 1360 3968
rect 1326 3858 1360 3896
rect 1326 3786 1360 3824
rect 1326 3714 1360 3752
rect 1326 3642 1360 3680
rect 1326 3570 1360 3608
rect 1326 3498 1360 3536
rect 1326 3426 1360 3464
rect 1326 3354 1360 3392
rect 1326 3282 1360 3320
rect 1326 3210 1360 3248
rect 1326 3138 1360 3176
rect 1326 3066 1360 3104
rect 1326 2994 1360 3032
rect 1326 2922 1360 2960
rect 1326 2850 1360 2888
rect 1326 2778 1360 2816
rect 1326 2706 1360 2744
rect 1634 2672 1655 2706
rect 1689 2672 3514 2706
rect 1326 2666 1360 2672
rect -1298 2570 -1195 2604
rect -1161 2570 -1127 2604
rect -1093 2570 -1059 2604
rect -1025 2570 -991 2604
rect -957 2570 -923 2604
rect -889 2570 -855 2604
rect -821 2570 -787 2604
rect -753 2570 -719 2604
rect -685 2570 -651 2604
rect -617 2570 -583 2604
rect -549 2570 -515 2604
rect -481 2570 -447 2604
rect -413 2570 -379 2604
rect -345 2570 -311 2604
rect -277 2570 -243 2604
rect -209 2570 -175 2604
rect -141 2570 -107 2604
rect -73 2570 -39 2604
rect -5 2570 29 2604
rect 63 2570 97 2604
rect 131 2570 165 2604
rect 199 2570 233 2604
rect 267 2570 301 2604
rect 335 2570 369 2604
rect 403 2570 437 2604
rect 471 2570 505 2604
rect 539 2570 573 2604
rect 607 2570 641 2604
rect 675 2570 709 2604
rect 743 2570 777 2604
rect 811 2570 845 2604
rect 879 2570 913 2604
rect 947 2570 981 2604
rect 1015 2570 1049 2604
rect 1083 2570 1117 2604
rect 1151 2570 1254 2604
rect -98 1838 20 1872
rect 54 1838 88 1872
rect 122 1838 156 1872
rect 190 1838 224 1872
rect 258 1838 292 1872
rect 326 1838 360 1872
rect 394 1838 428 1872
rect 462 1838 496 1872
rect 530 1838 564 1872
rect 598 1838 632 1872
rect 666 1838 700 1872
rect 734 1838 768 1872
rect 802 1838 836 1872
rect 870 1838 904 1872
rect 938 1838 972 1872
rect 1006 1838 1124 1872
rect -98 1767 -64 1838
rect 48 1736 64 1770
rect 98 1736 256 1770
rect 290 1736 448 1770
rect 482 1736 640 1770
rect 674 1736 832 1770
rect 866 1736 882 1770
rect 1090 1767 1124 1838
rect -98 1699 -64 1733
rect -98 1631 -64 1665
rect -98 1563 -64 1597
rect 16 1665 50 1702
rect 16 1594 50 1631
rect 112 1665 146 1702
rect 112 1594 146 1631
rect 208 1665 242 1702
rect 208 1594 242 1631
rect 304 1665 338 1702
rect 304 1594 338 1631
rect 400 1665 434 1702
rect 400 1594 434 1631
rect 496 1665 530 1702
rect 496 1594 530 1631
rect 592 1665 626 1702
rect 592 1594 626 1631
rect 688 1665 722 1702
rect 688 1594 722 1631
rect 784 1665 818 1702
rect 784 1594 818 1631
rect 880 1665 914 1702
rect 880 1594 914 1631
rect 976 1665 1010 1702
rect 976 1594 1010 1631
rect 1090 1699 1124 1733
rect 1090 1631 1124 1665
rect 1090 1563 1124 1597
rect -98 1458 -64 1529
rect 66 1526 116 1560
rect 150 1526 160 1560
rect 194 1526 352 1560
rect 386 1526 544 1560
rect 578 1526 736 1560
rect 770 1526 928 1560
rect 962 1526 978 1560
rect 1090 1458 1124 1529
rect -98 1424 20 1458
rect 54 1424 88 1458
rect 122 1424 156 1458
rect 190 1424 224 1458
rect 258 1424 292 1458
rect 326 1424 360 1458
rect 394 1424 428 1458
rect 462 1424 496 1458
rect 530 1424 564 1458
rect 598 1424 632 1458
rect 666 1424 700 1458
rect 734 1424 768 1458
rect 802 1424 836 1458
rect 870 1424 904 1458
rect 938 1424 972 1458
rect 1006 1424 1124 1458
rect 1196 1838 1314 1872
rect 1348 1838 1382 1872
rect 1416 1838 1450 1872
rect 1484 1838 1518 1872
rect 1552 1838 1586 1872
rect 1620 1838 1654 1872
rect 1688 1838 1722 1872
rect 1756 1838 1790 1872
rect 1824 1838 1858 1872
rect 1892 1838 1926 1872
rect 1960 1838 1994 1872
rect 2028 1838 2062 1872
rect 2096 1838 2130 1872
rect 2164 1838 2198 1872
rect 2232 1838 2266 1872
rect 2300 1838 2418 1872
rect 1196 1767 1230 1838
rect 1342 1736 1358 1770
rect 1392 1736 1550 1770
rect 1584 1736 1742 1770
rect 1776 1736 1934 1770
rect 1968 1736 2126 1770
rect 2160 1736 2302 1770
rect 2336 1736 2340 1770
rect 2384 1767 2418 1838
rect 1196 1699 1230 1733
rect 1196 1631 1230 1665
rect 1196 1563 1230 1597
rect 1310 1665 1344 1702
rect 1310 1594 1344 1631
rect 1406 1665 1440 1702
rect 1406 1594 1440 1631
rect 1502 1665 1536 1702
rect 1502 1594 1536 1631
rect 1598 1665 1632 1702
rect 1598 1594 1632 1631
rect 1694 1665 1728 1702
rect 1694 1594 1728 1631
rect 1790 1665 1824 1702
rect 1790 1594 1824 1631
rect 1886 1665 1920 1702
rect 1886 1594 1920 1631
rect 1982 1665 2016 1702
rect 1982 1594 2016 1631
rect 2078 1665 2112 1702
rect 2078 1594 2112 1631
rect 2174 1665 2208 1702
rect 2174 1594 2208 1631
rect 2270 1665 2304 1702
rect 2270 1594 2304 1631
rect 2384 1699 2418 1733
rect 2384 1631 2418 1665
rect 2384 1563 2418 1597
rect 1196 1458 1230 1529
rect 1438 1526 1454 1560
rect 1488 1526 1646 1560
rect 1680 1526 1838 1560
rect 1872 1526 2030 1560
rect 2064 1526 2222 1560
rect 2256 1526 2272 1560
rect 2384 1458 2418 1529
rect 1196 1424 1314 1458
rect 1348 1424 1382 1458
rect 1416 1424 1450 1458
rect 1484 1424 1518 1458
rect 1552 1424 1586 1458
rect 1620 1424 1654 1458
rect 1688 1424 1722 1458
rect 1756 1424 1790 1458
rect 1824 1424 1858 1458
rect 1892 1424 1926 1458
rect 1960 1424 1994 1458
rect 2028 1424 2062 1458
rect 2096 1424 2130 1458
rect 2164 1424 2198 1458
rect 2232 1424 2266 1458
rect 2300 1424 2418 1458
rect -98 838 -64 1424
rect 2380 840 2414 1424
rect 1192 806 1310 840
rect 1344 806 1378 840
rect 1412 806 1446 840
rect 1480 806 1514 840
rect 1548 806 1582 840
rect 1616 806 1650 840
rect 1684 806 1718 840
rect 1752 806 1786 840
rect 1820 806 1854 840
rect 1888 806 1922 840
rect 1956 806 1990 840
rect 2024 806 2058 840
rect 2092 806 2126 840
rect 2160 806 2194 840
rect 2228 806 2262 840
rect 2296 806 2414 840
rect 62 704 114 738
rect 148 704 974 738
rect 1192 735 1226 806
rect 1434 704 1450 738
rect 1484 704 1642 738
rect 1676 704 1834 738
rect 1868 704 2026 738
rect 2060 704 2218 738
rect 2252 704 2268 738
rect 2380 735 2414 806
rect 1192 667 1226 701
rect 1192 599 1226 633
rect 1192 531 1226 565
rect 1306 633 1340 670
rect 1306 562 1340 599
rect 1402 633 1436 670
rect 1402 562 1436 599
rect 1498 633 1532 670
rect 1498 562 1532 599
rect 1594 633 1628 670
rect 1594 562 1628 599
rect 1690 633 1724 670
rect 1690 562 1724 599
rect 1786 633 1820 670
rect 1786 562 1820 599
rect 1882 633 1916 670
rect 1882 562 1916 599
rect 1978 633 2012 670
rect 1978 562 2012 599
rect 2074 633 2108 670
rect 2074 562 2108 599
rect 2170 633 2204 670
rect 2170 562 2204 599
rect 2266 633 2300 670
rect 2266 562 2300 599
rect 2380 667 2414 701
rect 2380 599 2414 633
rect 44 494 878 528
rect 2380 531 2414 565
rect 1192 426 1226 497
rect 1338 494 1354 528
rect 1388 494 1546 528
rect 1580 494 1738 528
rect 1772 494 1930 528
rect 1964 494 2122 528
rect 2156 494 2296 528
rect 2330 494 2336 528
rect 2380 426 2414 497
rect -102 -392 -50 412
rect 1192 392 1310 426
rect 1344 392 1378 426
rect 1412 392 1446 426
rect 1480 392 1514 426
rect 1548 392 1582 426
rect 1616 392 1650 426
rect 1684 392 1718 426
rect 1752 392 1786 426
rect 1820 392 1854 426
rect 1888 392 1922 426
rect 1956 392 1990 426
rect 2024 392 2058 426
rect 2092 392 2126 426
rect 2160 392 2194 426
rect 2228 392 2262 426
rect 2296 392 2414 426
rect 2360 -394 2412 392
rect -943 -510 3271 -476
rect -949 -3262 -915 -3228
rect -881 -3262 3275 -3228
<< viali >>
rect -1191 6540 -1161 6574
rect -1161 6540 -1157 6574
rect -1119 6540 -1093 6574
rect -1093 6540 -1085 6574
rect -1047 6540 -1025 6574
rect -1025 6540 -1013 6574
rect -975 6540 -957 6574
rect -957 6540 -941 6574
rect -903 6540 -889 6574
rect -889 6540 -869 6574
rect -831 6540 -821 6574
rect -821 6540 -797 6574
rect -759 6540 -753 6574
rect -753 6540 -725 6574
rect -687 6540 -685 6574
rect -685 6540 -653 6574
rect -615 6540 -583 6574
rect -583 6540 -581 6574
rect -543 6540 -515 6574
rect -515 6540 -509 6574
rect -471 6540 -447 6574
rect -447 6540 -437 6574
rect -399 6540 -379 6574
rect -379 6540 -365 6574
rect -327 6540 -311 6574
rect -311 6540 -293 6574
rect -255 6540 -243 6574
rect -243 6540 -221 6574
rect -183 6540 -175 6574
rect -175 6540 -149 6574
rect -111 6540 -107 6574
rect -107 6540 -77 6574
rect -39 6540 -5 6574
rect 33 6540 63 6574
rect 63 6540 67 6574
rect 105 6540 131 6574
rect 131 6540 139 6574
rect 177 6540 199 6574
rect 199 6540 211 6574
rect 249 6540 267 6574
rect 267 6540 283 6574
rect 321 6540 335 6574
rect 335 6540 355 6574
rect 393 6540 403 6574
rect 403 6540 427 6574
rect 465 6540 471 6574
rect 471 6540 499 6574
rect 537 6540 539 6574
rect 539 6540 571 6574
rect 609 6540 641 6574
rect 641 6540 643 6574
rect 681 6540 709 6574
rect 709 6540 715 6574
rect 753 6540 777 6574
rect 777 6540 787 6574
rect 825 6540 845 6574
rect 845 6540 859 6574
rect 897 6540 913 6574
rect 913 6540 931 6574
rect 969 6540 981 6574
rect 981 6540 1003 6574
rect 1041 6540 1049 6574
rect 1049 6540 1075 6574
rect 1113 6540 1117 6574
rect 1117 6540 1147 6574
rect 1433 6540 1467 6574
rect 1505 6540 1539 6574
rect 1577 6540 1611 6574
rect 1649 6540 1683 6574
rect 1721 6540 1755 6574
rect 1793 6540 1827 6574
rect 1865 6540 1899 6574
rect 1937 6540 1971 6574
rect 2009 6540 2043 6574
rect 2081 6540 2115 6574
rect 2153 6540 2187 6574
rect 2225 6540 2259 6574
rect 2297 6540 2331 6574
rect 2369 6540 2403 6574
rect 2441 6540 2475 6574
rect 2513 6540 2547 6574
rect 2585 6540 2619 6574
rect 2657 6540 2691 6574
rect 2729 6540 2763 6574
rect 2801 6540 2835 6574
rect 2873 6540 2907 6574
rect 2945 6540 2979 6574
rect 3017 6540 3051 6574
rect 3089 6540 3123 6574
rect 3161 6540 3195 6574
rect 3233 6540 3267 6574
rect 3305 6540 3339 6574
rect 3377 6540 3411 6574
rect 3449 6540 3483 6574
rect 3521 6540 3555 6574
rect 3593 6540 3627 6574
rect 3665 6540 3699 6574
rect 3737 6540 3771 6574
rect -726 6438 -692 6472
rect 190 6438 224 6472
rect 1106 6438 1140 6472
rect 1220 6458 1254 6472
rect 1220 6438 1254 6458
rect -1184 6330 -1150 6364
rect -1184 6258 -1150 6292
rect -1184 6186 -1150 6220
rect -1184 6114 -1150 6148
rect -1184 6042 -1150 6076
rect -1184 5970 -1150 6004
rect -1184 5898 -1150 5932
rect -1184 5826 -1150 5860
rect -1184 5754 -1150 5788
rect -1184 5682 -1150 5716
rect -1184 5610 -1150 5644
rect -1184 5538 -1150 5572
rect -1184 5466 -1150 5500
rect -1184 5394 -1150 5428
rect -1184 5322 -1150 5356
rect -1184 5250 -1150 5284
rect -1184 5178 -1150 5212
rect -1184 5106 -1150 5140
rect -1184 5034 -1150 5068
rect -1184 4962 -1150 4996
rect -1184 4890 -1150 4924
rect -1184 4818 -1150 4852
rect -726 6330 -692 6364
rect -726 6258 -692 6292
rect -726 6186 -692 6220
rect -726 6114 -692 6148
rect -726 6042 -692 6076
rect -726 5970 -692 6004
rect -726 5898 -692 5932
rect -726 5826 -692 5860
rect -726 5754 -692 5788
rect -726 5682 -692 5716
rect -726 5610 -692 5644
rect -726 5538 -692 5572
rect -726 5466 -692 5500
rect -726 5394 -692 5428
rect -726 5322 -692 5356
rect -726 5250 -692 5284
rect -726 5178 -692 5212
rect -726 5106 -692 5140
rect -726 5034 -692 5068
rect -726 4962 -692 4996
rect -726 4890 -692 4924
rect -726 4818 -692 4852
rect -268 6330 -234 6364
rect -268 6258 -234 6292
rect -268 6186 -234 6220
rect -268 6114 -234 6148
rect -268 6042 -234 6076
rect -268 5970 -234 6004
rect -268 5898 -234 5932
rect -268 5826 -234 5860
rect -268 5754 -234 5788
rect -268 5682 -234 5716
rect -268 5610 -234 5644
rect -268 5538 -234 5572
rect -268 5466 -234 5500
rect -268 5394 -234 5428
rect -268 5322 -234 5356
rect -268 5250 -234 5284
rect -268 5178 -234 5212
rect -268 5106 -234 5140
rect -268 5034 -234 5068
rect -268 4962 -234 4996
rect -268 4890 -234 4924
rect -268 4818 -234 4852
rect 190 6330 224 6364
rect 190 6258 224 6292
rect 190 6186 224 6220
rect 190 6114 224 6148
rect 190 6042 224 6076
rect 190 5970 224 6004
rect 190 5898 224 5932
rect 190 5826 224 5860
rect 190 5754 224 5788
rect 190 5682 224 5716
rect 190 5610 224 5644
rect 190 5538 224 5572
rect 190 5466 224 5500
rect 190 5394 224 5428
rect 190 5322 224 5356
rect 190 5250 224 5284
rect 190 5178 224 5212
rect 190 5106 224 5140
rect 190 5034 224 5068
rect 190 4962 224 4996
rect 190 4890 224 4924
rect 190 4818 224 4852
rect 648 6330 682 6364
rect 648 6258 682 6292
rect 648 6186 682 6220
rect 648 6114 682 6148
rect 648 6042 682 6076
rect 648 5970 682 6004
rect 648 5898 682 5932
rect 648 5826 682 5860
rect 648 5754 682 5788
rect 648 5682 682 5716
rect 648 5610 682 5644
rect 648 5538 682 5572
rect 648 5466 682 5500
rect 648 5394 682 5428
rect 648 5322 682 5356
rect 648 5250 682 5284
rect 648 5178 682 5212
rect 648 5106 682 5140
rect 648 5034 682 5068
rect 648 4962 682 4996
rect 648 4890 682 4924
rect 648 4818 682 4852
rect 1106 6330 1140 6364
rect 1106 6258 1140 6292
rect 1106 6186 1140 6220
rect 1106 6114 1140 6148
rect 1106 6042 1140 6076
rect 1106 5970 1140 6004
rect 1106 5898 1140 5932
rect 1106 5826 1140 5860
rect 1106 5754 1140 5788
rect 1106 5682 1140 5716
rect 1106 5610 1140 5644
rect 1106 5538 1140 5572
rect 1106 5466 1140 5500
rect 1106 5394 1140 5428
rect 1106 5322 1140 5356
rect 1106 5250 1140 5284
rect 1106 5178 1140 5212
rect 1106 5106 1140 5140
rect 1106 5034 1140 5068
rect 1106 4962 1140 4996
rect 1106 4890 1140 4924
rect 1106 4818 1140 4852
rect 1220 6390 1254 6400
rect 1220 6366 1254 6390
rect 1220 6322 1254 6328
rect 1220 6294 1254 6322
rect 1220 6254 1254 6256
rect 1220 6222 1254 6254
rect 1220 6152 1254 6184
rect 1220 6150 1254 6152
rect 1220 6084 1254 6112
rect 1220 6078 1254 6084
rect 1220 6016 1254 6040
rect 1220 6006 1254 6016
rect 1220 5948 1254 5968
rect 1220 5934 1254 5948
rect 1220 5880 1254 5896
rect 1220 5862 1254 5880
rect 1220 5812 1254 5824
rect 1220 5790 1254 5812
rect 1220 5744 1254 5752
rect 1220 5718 1254 5744
rect 1220 5676 1254 5680
rect 1220 5646 1254 5676
rect 1220 5574 1254 5608
rect 1220 5506 1254 5536
rect 1220 5502 1254 5506
rect 1220 5438 1254 5464
rect 1220 5430 1254 5438
rect 1220 5370 1254 5392
rect 1220 5358 1254 5370
rect 1220 5302 1254 5320
rect 1220 5286 1254 5302
rect 1220 5234 1254 5248
rect 1220 5214 1254 5234
rect 1220 5166 1254 5176
rect 1220 5142 1254 5166
rect 1220 5098 1254 5104
rect 1220 5070 1254 5098
rect 1220 5030 1254 5032
rect 1220 4998 1254 5030
rect 1220 4928 1254 4960
rect 1220 4926 1254 4928
rect 1220 4860 1254 4888
rect 1220 4854 1254 4860
rect 1220 4792 1254 4816
rect 1220 4782 1254 4792
rect -726 4710 -692 4744
rect 190 4710 224 4744
rect 1106 4710 1140 4744
rect 1220 4724 1254 4744
rect 1220 4710 1254 4724
rect 1326 6438 1360 6472
rect 1440 6438 1474 6472
rect 2356 6438 2390 6472
rect 3272 6438 3306 6472
rect 1326 6366 1360 6400
rect 1326 6294 1360 6328
rect 1326 6222 1360 6256
rect 1326 6150 1360 6184
rect 1326 6078 1360 6112
rect 1326 6006 1360 6040
rect 1326 5934 1360 5968
rect 1326 5862 1360 5896
rect 1326 5790 1360 5824
rect 1326 5718 1360 5752
rect 1326 5646 1360 5680
rect 1326 5574 1360 5608
rect 1326 5502 1360 5536
rect 1326 5430 1360 5464
rect 1326 5358 1360 5392
rect 1326 5286 1360 5320
rect 1326 5214 1360 5248
rect 1326 5142 1360 5176
rect 1326 5070 1360 5104
rect 1326 4998 1360 5032
rect 1326 4926 1360 4960
rect 1326 4854 1360 4888
rect 1326 4782 1360 4816
rect 1326 4710 1360 4744
rect 1440 4710 1474 4744
rect 2356 4710 2390 4744
rect 3272 4710 3306 4744
rect -1263 4608 -1229 4642
rect -1191 4608 -1161 4642
rect -1161 4608 -1157 4642
rect -1119 4608 -1093 4642
rect -1093 4608 -1085 4642
rect -1047 4608 -1025 4642
rect -1025 4608 -1013 4642
rect -975 4608 -957 4642
rect -957 4608 -941 4642
rect -903 4608 -889 4642
rect -889 4608 -869 4642
rect -831 4608 -821 4642
rect -821 4608 -797 4642
rect -759 4608 -753 4642
rect -753 4608 -725 4642
rect -687 4608 -685 4642
rect -685 4608 -653 4642
rect -615 4608 -583 4642
rect -583 4608 -581 4642
rect -543 4608 -515 4642
rect -515 4608 -509 4642
rect -471 4608 -447 4642
rect -447 4608 -437 4642
rect -399 4608 -379 4642
rect -379 4608 -365 4642
rect -327 4608 -311 4642
rect -311 4608 -293 4642
rect -255 4608 -243 4642
rect -243 4608 -221 4642
rect -183 4608 -175 4642
rect -175 4608 -149 4642
rect -111 4608 -107 4642
rect -107 4608 -77 4642
rect -39 4608 -5 4642
rect 33 4608 63 4642
rect 63 4608 67 4642
rect 105 4608 131 4642
rect 131 4608 139 4642
rect 177 4608 199 4642
rect 199 4608 211 4642
rect 249 4608 267 4642
rect 267 4608 283 4642
rect 321 4608 335 4642
rect 335 4608 355 4642
rect 393 4608 403 4642
rect 403 4608 427 4642
rect 465 4608 471 4642
rect 471 4608 499 4642
rect 537 4608 539 4642
rect 539 4608 571 4642
rect 609 4608 641 4642
rect 641 4608 643 4642
rect 681 4608 709 4642
rect 709 4608 715 4642
rect 753 4608 777 4642
rect 777 4608 787 4642
rect 825 4608 845 4642
rect 845 4608 859 4642
rect 897 4608 913 4642
rect 913 4608 931 4642
rect 969 4608 981 4642
rect 981 4608 1003 4642
rect 1041 4608 1049 4642
rect 1049 4608 1075 4642
rect 1113 4608 1117 4642
rect 1117 4608 1147 4642
rect 1185 4608 1219 4642
rect -1263 4502 -1229 4536
rect -1191 4502 -1161 4536
rect -1161 4502 -1157 4536
rect -1119 4502 -1093 4536
rect -1093 4502 -1085 4536
rect -1047 4502 -1025 4536
rect -1025 4502 -1013 4536
rect -975 4502 -957 4536
rect -957 4502 -941 4536
rect -903 4502 -889 4536
rect -889 4502 -869 4536
rect -831 4502 -821 4536
rect -821 4502 -797 4536
rect -759 4502 -753 4536
rect -753 4502 -725 4536
rect -687 4502 -685 4536
rect -685 4502 -653 4536
rect -615 4502 -583 4536
rect -583 4502 -581 4536
rect -543 4502 -515 4536
rect -515 4502 -509 4536
rect -471 4502 -447 4536
rect -447 4502 -437 4536
rect -399 4502 -379 4536
rect -379 4502 -365 4536
rect -327 4502 -311 4536
rect -311 4502 -293 4536
rect -255 4502 -243 4536
rect -243 4502 -221 4536
rect -183 4502 -175 4536
rect -175 4502 -149 4536
rect -111 4502 -107 4536
rect -107 4502 -77 4536
rect -39 4502 -5 4536
rect 33 4502 63 4536
rect 63 4502 67 4536
rect 105 4502 131 4536
rect 131 4502 139 4536
rect 177 4502 199 4536
rect 199 4502 211 4536
rect 249 4502 267 4536
rect 267 4502 283 4536
rect 321 4502 335 4536
rect 335 4502 355 4536
rect 393 4502 403 4536
rect 403 4502 427 4536
rect 465 4502 471 4536
rect 471 4502 499 4536
rect 537 4502 539 4536
rect 539 4502 571 4536
rect 609 4502 641 4536
rect 641 4502 643 4536
rect 681 4502 709 4536
rect 709 4502 715 4536
rect 753 4502 777 4536
rect 777 4502 787 4536
rect 825 4502 845 4536
rect 845 4502 859 4536
rect 897 4502 913 4536
rect 913 4502 931 4536
rect 969 4502 981 4536
rect 981 4502 1003 4536
rect 1041 4502 1049 4536
rect 1049 4502 1075 4536
rect 1113 4502 1117 4536
rect 1117 4502 1147 4536
rect 1185 4502 1219 4536
rect 1220 4420 1254 4434
rect 1220 4400 1254 4420
rect -1184 4292 -1150 4326
rect -1184 4220 -1150 4254
rect -1184 4148 -1150 4182
rect -1184 4076 -1150 4110
rect -1184 4004 -1150 4038
rect -1184 3932 -1150 3966
rect -1184 3860 -1150 3894
rect -1184 3788 -1150 3822
rect -1184 3716 -1150 3750
rect -1184 3644 -1150 3678
rect -1184 3572 -1150 3606
rect -1184 3500 -1150 3534
rect -1184 3428 -1150 3462
rect -1184 3356 -1150 3390
rect -1184 3284 -1150 3318
rect -1184 3212 -1150 3246
rect -1184 3140 -1150 3174
rect -1184 3068 -1150 3102
rect -1184 2996 -1150 3030
rect -1184 2924 -1150 2958
rect -1184 2852 -1150 2886
rect -1184 2780 -1150 2814
rect -726 4292 -692 4326
rect -726 4220 -692 4254
rect -726 4148 -692 4182
rect -726 4076 -692 4110
rect -726 4004 -692 4038
rect -726 3932 -692 3966
rect -726 3860 -692 3894
rect -726 3788 -692 3822
rect -726 3716 -692 3750
rect -726 3644 -692 3678
rect -726 3572 -692 3606
rect -726 3500 -692 3534
rect -726 3428 -692 3462
rect -726 3356 -692 3390
rect -726 3284 -692 3318
rect -726 3212 -692 3246
rect -726 3140 -692 3174
rect -726 3068 -692 3102
rect -726 2996 -692 3030
rect -726 2924 -692 2958
rect -726 2852 -692 2886
rect -726 2780 -692 2814
rect -268 4292 -234 4326
rect -268 4220 -234 4254
rect -268 4148 -234 4182
rect -268 4076 -234 4110
rect -268 4004 -234 4038
rect -268 3932 -234 3966
rect -268 3860 -234 3894
rect -268 3788 -234 3822
rect -268 3716 -234 3750
rect -268 3644 -234 3678
rect -268 3572 -234 3606
rect -268 3500 -234 3534
rect -268 3428 -234 3462
rect -268 3356 -234 3390
rect -268 3284 -234 3318
rect -268 3212 -234 3246
rect -268 3140 -234 3174
rect -268 3068 -234 3102
rect -268 2996 -234 3030
rect -268 2924 -234 2958
rect -268 2852 -234 2886
rect -268 2780 -234 2814
rect 190 4292 224 4326
rect 190 4220 224 4254
rect 190 4148 224 4182
rect 190 4076 224 4110
rect 190 4004 224 4038
rect 190 3932 224 3966
rect 190 3860 224 3894
rect 190 3788 224 3822
rect 190 3716 224 3750
rect 190 3644 224 3678
rect 190 3572 224 3606
rect 190 3500 224 3534
rect 190 3428 224 3462
rect 190 3356 224 3390
rect 190 3284 224 3318
rect 190 3212 224 3246
rect 190 3140 224 3174
rect 190 3068 224 3102
rect 190 2996 224 3030
rect 190 2924 224 2958
rect 190 2852 224 2886
rect 190 2780 224 2814
rect 648 4292 682 4326
rect 648 4220 682 4254
rect 648 4148 682 4182
rect 648 4076 682 4110
rect 648 4004 682 4038
rect 648 3932 682 3966
rect 648 3860 682 3894
rect 648 3788 682 3822
rect 648 3716 682 3750
rect 648 3644 682 3678
rect 648 3572 682 3606
rect 648 3500 682 3534
rect 648 3428 682 3462
rect 648 3356 682 3390
rect 648 3284 682 3318
rect 648 3212 682 3246
rect 648 3140 682 3174
rect 648 3068 682 3102
rect 648 2996 682 3030
rect 648 2924 682 2958
rect 648 2852 682 2886
rect 648 2780 682 2814
rect 1106 4292 1140 4326
rect 1106 4220 1140 4254
rect 1106 4148 1140 4182
rect 1106 4076 1140 4110
rect 1106 4004 1140 4038
rect 1106 3932 1140 3966
rect 1106 3860 1140 3894
rect 1106 3788 1140 3822
rect 1106 3716 1140 3750
rect 1106 3644 1140 3678
rect 1106 3572 1140 3606
rect 1106 3500 1140 3534
rect 1106 3428 1140 3462
rect 1106 3356 1140 3390
rect 1106 3284 1140 3318
rect 1106 3212 1140 3246
rect 1106 3140 1140 3174
rect 1106 3068 1140 3102
rect 1106 2996 1140 3030
rect 1106 2924 1140 2958
rect 1106 2852 1140 2886
rect 1106 2780 1140 2814
rect 1220 4352 1254 4362
rect 1220 4328 1254 4352
rect 1220 4284 1254 4290
rect 1220 4256 1254 4284
rect 1220 4216 1254 4218
rect 1220 4184 1254 4216
rect 1220 4114 1254 4146
rect 1220 4112 1254 4114
rect 1220 4046 1254 4074
rect 1220 4040 1254 4046
rect 1220 3978 1254 4002
rect 1220 3968 1254 3978
rect 1220 3910 1254 3930
rect 1220 3896 1254 3910
rect 1220 3842 1254 3858
rect 1220 3824 1254 3842
rect 1220 3774 1254 3786
rect 1220 3752 1254 3774
rect 1220 3706 1254 3714
rect 1220 3680 1254 3706
rect 1220 3638 1254 3642
rect 1220 3608 1254 3638
rect 1220 3536 1254 3570
rect 1220 3468 1254 3498
rect 1220 3464 1254 3468
rect 1220 3400 1254 3426
rect 1220 3392 1254 3400
rect 1220 3332 1254 3354
rect 1220 3320 1254 3332
rect 1220 3264 1254 3282
rect 1220 3248 1254 3264
rect 1220 3196 1254 3210
rect 1220 3176 1254 3196
rect 1220 3128 1254 3138
rect 1220 3104 1254 3128
rect 1220 3060 1254 3066
rect 1220 3032 1254 3060
rect 1220 2992 1254 2994
rect 1220 2960 1254 2992
rect 1220 2890 1254 2922
rect 1220 2888 1254 2890
rect 1220 2822 1254 2850
rect 1220 2816 1254 2822
rect 1220 2754 1254 2778
rect 1220 2744 1254 2754
rect 860 2672 894 2706
rect 1220 2686 1254 2706
rect 1220 2672 1254 2686
rect 1326 4400 1360 4434
rect 1326 4328 1360 4362
rect 1326 4256 1360 4290
rect 1326 4184 1360 4218
rect 1326 4112 1360 4146
rect 1326 4040 1360 4074
rect 1326 3968 1360 4002
rect 1326 3896 1360 3930
rect 1326 3824 1360 3858
rect 1326 3752 1360 3786
rect 1326 3680 1360 3714
rect 1326 3608 1360 3642
rect 1326 3536 1360 3570
rect 1326 3464 1360 3498
rect 1326 3392 1360 3426
rect 1326 3320 1360 3354
rect 1326 3248 1360 3282
rect 1326 3176 1360 3210
rect 1326 3104 1360 3138
rect 1326 3032 1360 3066
rect 1326 2960 1360 2994
rect 1326 2888 1360 2922
rect 1326 2816 1360 2850
rect 1326 2744 1360 2778
rect 1326 2672 1360 2706
rect 1655 2672 1689 2706
rect 16 1631 50 1665
rect 112 1631 146 1665
rect 208 1631 242 1665
rect 304 1631 338 1665
rect 400 1631 434 1665
rect 496 1631 530 1665
rect 592 1631 626 1665
rect 688 1631 722 1665
rect 784 1631 818 1665
rect 880 1631 914 1665
rect 976 1631 1010 1665
rect 116 1526 150 1560
rect 2302 1736 2336 1770
rect 1310 1631 1344 1665
rect 1406 1631 1440 1665
rect 1502 1631 1536 1665
rect 1598 1631 1632 1665
rect 1694 1631 1728 1665
rect 1790 1631 1824 1665
rect 1886 1631 1920 1665
rect 1982 1631 2016 1665
rect 2078 1631 2112 1665
rect 2174 1631 2208 1665
rect 2270 1631 2304 1665
rect 114 704 148 738
rect 1306 599 1340 633
rect 1402 599 1436 633
rect 1498 599 1532 633
rect 1594 599 1628 633
rect 1690 599 1724 633
rect 1786 599 1820 633
rect 1882 599 1916 633
rect 1978 599 2012 633
rect 2074 599 2108 633
rect 2170 599 2204 633
rect 2266 599 2300 633
rect 2296 494 2330 528
rect -915 -3262 -881 -3228
<< metal1 >>
rect -1212 6605 3792 6610
rect -1212 6580 -1200 6605
rect -1214 6553 -1200 6580
rect -1148 6553 -1136 6605
rect -1084 6553 -1072 6605
rect -1020 6574 -1008 6605
rect -956 6574 -944 6605
rect -892 6574 -880 6605
rect -828 6574 -816 6605
rect -764 6574 -752 6605
rect -1013 6553 -1008 6574
rect -764 6553 -759 6574
rect -700 6553 -688 6605
rect -636 6553 -624 6605
rect -572 6553 -560 6605
rect -508 6553 -496 6605
rect -444 6574 -432 6605
rect -380 6574 -368 6605
rect -316 6574 -304 6605
rect -252 6574 -240 6605
rect -188 6574 -176 6605
rect -437 6553 -432 6574
rect -188 6553 -183 6574
rect -124 6553 -112 6605
rect -60 6553 -48 6605
rect 4 6553 16 6605
rect 68 6553 80 6605
rect 132 6574 144 6605
rect 196 6574 208 6605
rect 260 6574 272 6605
rect 324 6574 336 6605
rect 388 6574 400 6605
rect 139 6553 144 6574
rect 388 6553 393 6574
rect 452 6553 464 6605
rect 516 6553 528 6605
rect 580 6553 592 6605
rect 644 6553 656 6605
rect 708 6574 720 6605
rect 772 6574 784 6605
rect 836 6574 848 6605
rect 900 6574 912 6605
rect 964 6574 976 6605
rect 715 6553 720 6574
rect 964 6553 969 6574
rect 1028 6553 1040 6605
rect 1092 6553 1104 6605
rect 1156 6553 1168 6605
rect 1220 6553 1232 6605
rect 1284 6553 1296 6605
rect 1348 6553 1360 6605
rect 1412 6553 1424 6605
rect 1476 6553 1488 6605
rect 1540 6553 1552 6605
rect 1604 6574 1616 6605
rect 1668 6574 1680 6605
rect 1732 6574 1744 6605
rect 1796 6574 1808 6605
rect 1860 6574 1872 6605
rect 1611 6553 1616 6574
rect 1860 6553 1865 6574
rect 1924 6553 1936 6605
rect 1988 6553 2000 6605
rect 2052 6553 2064 6605
rect 2116 6553 2128 6605
rect 2180 6574 2192 6605
rect 2244 6574 2256 6605
rect 2308 6574 2320 6605
rect 2372 6574 2384 6605
rect 2436 6574 2448 6605
rect 2187 6553 2192 6574
rect 2436 6553 2441 6574
rect 2500 6553 2512 6605
rect 2564 6553 2576 6605
rect 2628 6553 2640 6605
rect 2692 6553 2704 6605
rect 2756 6574 2768 6605
rect 2820 6574 2832 6605
rect 2884 6574 2896 6605
rect 2948 6574 2960 6605
rect 3012 6574 3024 6605
rect 2763 6553 2768 6574
rect 3012 6553 3017 6574
rect 3076 6553 3088 6605
rect 3140 6553 3152 6605
rect 3204 6553 3216 6605
rect 3268 6553 3280 6605
rect 3332 6574 3344 6605
rect 3396 6574 3408 6605
rect 3460 6574 3472 6605
rect 3524 6574 3536 6605
rect 3588 6574 3600 6605
rect 3339 6553 3344 6574
rect 3588 6553 3593 6574
rect 3652 6553 3664 6605
rect 3716 6553 3728 6605
rect 3780 6580 3792 6605
rect 3780 6553 3794 6580
rect -1214 6540 -1191 6553
rect -1157 6540 -1119 6553
rect -1085 6540 -1047 6553
rect -1013 6540 -975 6553
rect -941 6540 -903 6553
rect -869 6540 -831 6553
rect -797 6540 -759 6553
rect -725 6540 -687 6553
rect -653 6540 -615 6553
rect -581 6540 -543 6553
rect -509 6540 -471 6553
rect -437 6540 -399 6553
rect -365 6540 -327 6553
rect -293 6540 -255 6553
rect -221 6540 -183 6553
rect -149 6540 -111 6553
rect -77 6540 -39 6553
rect -5 6540 33 6553
rect 67 6540 105 6553
rect 139 6540 177 6553
rect 211 6540 249 6553
rect 283 6540 321 6553
rect 355 6540 393 6553
rect 427 6540 465 6553
rect 499 6540 537 6553
rect 571 6540 609 6553
rect 643 6540 681 6553
rect 715 6540 753 6553
rect 787 6540 825 6553
rect 859 6540 897 6553
rect 931 6540 969 6553
rect 1003 6540 1041 6553
rect 1075 6540 1113 6553
rect 1147 6548 1433 6553
rect 1147 6540 1170 6548
rect -1214 6534 1170 6540
rect 1410 6540 1433 6548
rect 1467 6540 1505 6553
rect 1539 6540 1577 6553
rect 1611 6540 1649 6553
rect 1683 6540 1721 6553
rect 1755 6540 1793 6553
rect 1827 6540 1865 6553
rect 1899 6540 1937 6553
rect 1971 6540 2009 6553
rect 2043 6540 2081 6553
rect 2115 6540 2153 6553
rect 2187 6540 2225 6553
rect 2259 6540 2297 6553
rect 2331 6540 2369 6553
rect 2403 6540 2441 6553
rect 2475 6540 2513 6553
rect 2547 6540 2585 6553
rect 2619 6540 2657 6553
rect 2691 6540 2729 6553
rect 2763 6540 2801 6553
rect 2835 6540 2873 6553
rect 2907 6540 2945 6553
rect 2979 6540 3017 6553
rect 3051 6540 3089 6553
rect 3123 6540 3161 6553
rect 3195 6540 3233 6553
rect 3267 6540 3305 6553
rect 3339 6540 3377 6553
rect 3411 6540 3449 6553
rect 3483 6540 3521 6553
rect 3555 6540 3593 6553
rect 3627 6540 3665 6553
rect 3699 6540 3737 6553
rect 3771 6540 3794 6553
rect 1410 6534 3794 6540
rect -742 6472 -676 6482
rect -742 6438 -726 6472
rect -692 6438 -676 6472
rect -1190 6364 -1144 6391
rect -1190 6330 -1184 6364
rect -1150 6330 -1144 6364
rect -1190 6292 -1144 6330
rect -1190 6258 -1184 6292
rect -1150 6258 -1144 6292
rect -1190 6220 -1144 6258
rect -1190 6186 -1184 6220
rect -1150 6186 -1144 6220
rect -1190 6148 -1144 6186
rect -1190 6114 -1184 6148
rect -1150 6114 -1144 6148
rect -1190 6076 -1144 6114
rect -1190 6042 -1184 6076
rect -1150 6042 -1144 6076
rect -1190 6004 -1144 6042
rect -1190 5970 -1184 6004
rect -1150 5970 -1144 6004
rect -1190 5932 -1144 5970
rect -1190 5898 -1184 5932
rect -1150 5898 -1144 5932
rect -1190 5860 -1144 5898
rect -1190 5826 -1184 5860
rect -1150 5826 -1144 5860
rect -1190 5788 -1144 5826
rect -1190 5754 -1184 5788
rect -1150 5754 -1144 5788
rect -1190 5716 -1144 5754
rect -1190 5682 -1184 5716
rect -1150 5682 -1144 5716
rect -1190 5644 -1144 5682
rect -1190 5610 -1184 5644
rect -1150 5610 -1144 5644
rect -1190 5572 -1144 5610
rect -1190 5538 -1184 5572
rect -1150 5538 -1144 5572
rect -1190 5500 -1144 5538
rect -1190 5466 -1184 5500
rect -1150 5466 -1144 5500
rect -1190 5428 -1144 5466
rect -1190 5394 -1184 5428
rect -1150 5394 -1144 5428
rect -1190 5356 -1144 5394
rect -1190 5322 -1184 5356
rect -1150 5322 -1144 5356
rect -1190 5284 -1144 5322
rect -1190 5250 -1184 5284
rect -1150 5250 -1144 5284
rect -1190 5212 -1144 5250
rect -1190 5178 -1184 5212
rect -1150 5178 -1144 5212
rect -1190 5140 -1144 5178
rect -1190 5106 -1184 5140
rect -1150 5106 -1144 5140
rect -1190 5068 -1144 5106
rect -1190 5034 -1184 5068
rect -1150 5034 -1144 5068
rect -1190 4996 -1144 5034
rect -1190 4962 -1184 4996
rect -1150 4962 -1144 4996
rect -1190 4924 -1144 4962
rect -1190 4890 -1184 4924
rect -1150 4890 -1144 4924
rect -1190 4852 -1144 4890
rect -1190 4818 -1184 4852
rect -1150 4818 -1144 4852
rect -1190 4648 -1144 4818
rect -742 6385 -676 6438
rect 174 6472 240 6482
rect 174 6438 190 6472
rect 224 6438 240 6472
rect -742 6333 -735 6385
rect -683 6333 -676 6385
rect -742 6330 -726 6333
rect -692 6330 -676 6333
rect -742 6321 -676 6330
rect -742 6269 -735 6321
rect -683 6269 -676 6321
rect -742 6258 -726 6269
rect -692 6258 -676 6269
rect -742 6257 -676 6258
rect -742 6205 -735 6257
rect -683 6205 -676 6257
rect -742 6193 -726 6205
rect -692 6193 -676 6205
rect -742 6141 -735 6193
rect -683 6141 -676 6193
rect -742 6129 -726 6141
rect -692 6129 -676 6141
rect -742 6077 -735 6129
rect -683 6077 -676 6129
rect -742 6076 -676 6077
rect -742 6065 -726 6076
rect -692 6065 -676 6076
rect -742 6013 -735 6065
rect -683 6013 -676 6065
rect -742 6004 -676 6013
rect -742 6001 -726 6004
rect -692 6001 -676 6004
rect -742 5949 -735 6001
rect -683 5949 -676 6001
rect -742 5937 -676 5949
rect -742 5885 -735 5937
rect -683 5885 -676 5937
rect -742 5873 -676 5885
rect -742 5821 -735 5873
rect -683 5821 -676 5873
rect -742 5809 -676 5821
rect -742 5757 -735 5809
rect -683 5757 -676 5809
rect -742 5754 -726 5757
rect -692 5754 -676 5757
rect -742 5745 -676 5754
rect -742 5693 -735 5745
rect -683 5693 -676 5745
rect -742 5682 -726 5693
rect -692 5682 -676 5693
rect -742 5681 -676 5682
rect -742 5629 -735 5681
rect -683 5629 -676 5681
rect -742 5617 -726 5629
rect -692 5617 -676 5629
rect -742 5565 -735 5617
rect -683 5565 -676 5617
rect -742 5553 -726 5565
rect -692 5553 -676 5565
rect -742 5501 -735 5553
rect -683 5501 -676 5553
rect -742 5500 -676 5501
rect -742 5489 -726 5500
rect -692 5489 -676 5500
rect -742 5437 -735 5489
rect -683 5437 -676 5489
rect -742 5428 -676 5437
rect -742 5425 -726 5428
rect -692 5425 -676 5428
rect -742 5373 -735 5425
rect -683 5373 -676 5425
rect -742 5361 -676 5373
rect -742 5309 -735 5361
rect -683 5309 -676 5361
rect -742 5297 -676 5309
rect -742 5245 -735 5297
rect -683 5245 -676 5297
rect -742 5233 -676 5245
rect -742 5181 -735 5233
rect -683 5181 -676 5233
rect -742 5178 -726 5181
rect -692 5178 -676 5181
rect -742 5169 -676 5178
rect -742 5117 -735 5169
rect -683 5117 -676 5169
rect -742 5106 -726 5117
rect -692 5106 -676 5117
rect -742 5105 -676 5106
rect -742 5053 -735 5105
rect -683 5053 -676 5105
rect -742 5041 -726 5053
rect -692 5041 -676 5053
rect -742 4989 -735 5041
rect -683 4989 -676 5041
rect -742 4977 -726 4989
rect -692 4977 -676 4989
rect -742 4925 -735 4977
rect -683 4925 -676 4977
rect -742 4924 -676 4925
rect -742 4913 -726 4924
rect -692 4913 -676 4924
rect -742 4861 -735 4913
rect -683 4861 -676 4913
rect -742 4852 -676 4861
rect -742 4849 -726 4852
rect -692 4849 -676 4852
rect -742 4797 -735 4849
rect -683 4797 -676 4849
rect -742 4744 -676 4797
rect -742 4710 -726 4744
rect -692 4710 -676 4744
rect -742 4694 -676 4710
rect -274 6364 -228 6391
rect -274 6330 -268 6364
rect -234 6330 -228 6364
rect -274 6292 -228 6330
rect -274 6258 -268 6292
rect -234 6258 -228 6292
rect -274 6220 -228 6258
rect -274 6186 -268 6220
rect -234 6186 -228 6220
rect -274 6148 -228 6186
rect -274 6114 -268 6148
rect -234 6114 -228 6148
rect -274 6076 -228 6114
rect -274 6042 -268 6076
rect -234 6042 -228 6076
rect -274 6004 -228 6042
rect -274 5970 -268 6004
rect -234 5970 -228 6004
rect -274 5932 -228 5970
rect -274 5898 -268 5932
rect -234 5898 -228 5932
rect -274 5860 -228 5898
rect -274 5826 -268 5860
rect -234 5826 -228 5860
rect -274 5788 -228 5826
rect -274 5754 -268 5788
rect -234 5754 -228 5788
rect -274 5716 -228 5754
rect -274 5682 -268 5716
rect -234 5682 -228 5716
rect -274 5644 -228 5682
rect -274 5610 -268 5644
rect -234 5610 -228 5644
rect -274 5572 -228 5610
rect -274 5538 -268 5572
rect -234 5538 -228 5572
rect -274 5500 -228 5538
rect -274 5466 -268 5500
rect -234 5466 -228 5500
rect -274 5428 -228 5466
rect -274 5394 -268 5428
rect -234 5394 -228 5428
rect -274 5356 -228 5394
rect -274 5322 -268 5356
rect -234 5322 -228 5356
rect -274 5284 -228 5322
rect -274 5250 -268 5284
rect -234 5250 -228 5284
rect -274 5212 -228 5250
rect -274 5178 -268 5212
rect -234 5178 -228 5212
rect -274 5140 -228 5178
rect -274 5106 -268 5140
rect -234 5106 -228 5140
rect -274 5068 -228 5106
rect -274 5034 -268 5068
rect -234 5034 -228 5068
rect -274 4996 -228 5034
rect -274 4962 -268 4996
rect -234 4962 -228 4996
rect -274 4924 -228 4962
rect -274 4890 -268 4924
rect -234 4890 -228 4924
rect -274 4852 -228 4890
rect -274 4818 -268 4852
rect -234 4818 -228 4852
rect -274 4648 -228 4818
rect 174 6385 240 6438
rect 1090 6472 1156 6482
rect 1090 6438 1106 6472
rect 1140 6438 1156 6472
rect 174 6333 181 6385
rect 233 6333 240 6385
rect 174 6330 190 6333
rect 224 6330 240 6333
rect 174 6321 240 6330
rect 174 6269 181 6321
rect 233 6269 240 6321
rect 174 6258 190 6269
rect 224 6258 240 6269
rect 174 6257 240 6258
rect 174 6205 181 6257
rect 233 6205 240 6257
rect 174 6193 190 6205
rect 224 6193 240 6205
rect 174 6141 181 6193
rect 233 6141 240 6193
rect 174 6129 190 6141
rect 224 6129 240 6141
rect 174 6077 181 6129
rect 233 6077 240 6129
rect 174 6076 240 6077
rect 174 6065 190 6076
rect 224 6065 240 6076
rect 174 6013 181 6065
rect 233 6013 240 6065
rect 174 6004 240 6013
rect 174 6001 190 6004
rect 224 6001 240 6004
rect 174 5949 181 6001
rect 233 5949 240 6001
rect 174 5937 240 5949
rect 174 5885 181 5937
rect 233 5885 240 5937
rect 174 5873 240 5885
rect 174 5821 181 5873
rect 233 5821 240 5873
rect 174 5809 240 5821
rect 174 5757 181 5809
rect 233 5757 240 5809
rect 174 5754 190 5757
rect 224 5754 240 5757
rect 174 5745 240 5754
rect 174 5693 181 5745
rect 233 5693 240 5745
rect 174 5682 190 5693
rect 224 5682 240 5693
rect 174 5681 240 5682
rect 174 5629 181 5681
rect 233 5629 240 5681
rect 174 5617 190 5629
rect 224 5617 240 5629
rect 174 5565 181 5617
rect 233 5565 240 5617
rect 174 5553 190 5565
rect 224 5553 240 5565
rect 174 5501 181 5553
rect 233 5501 240 5553
rect 174 5500 240 5501
rect 174 5489 190 5500
rect 224 5489 240 5500
rect 174 5437 181 5489
rect 233 5437 240 5489
rect 174 5428 240 5437
rect 174 5425 190 5428
rect 224 5425 240 5428
rect 174 5373 181 5425
rect 233 5373 240 5425
rect 174 5361 240 5373
rect 174 5309 181 5361
rect 233 5309 240 5361
rect 174 5297 240 5309
rect 174 5245 181 5297
rect 233 5245 240 5297
rect 174 5233 240 5245
rect 174 5181 181 5233
rect 233 5181 240 5233
rect 174 5178 190 5181
rect 224 5178 240 5181
rect 174 5169 240 5178
rect 174 5117 181 5169
rect 233 5117 240 5169
rect 174 5106 190 5117
rect 224 5106 240 5117
rect 174 5105 240 5106
rect 174 5053 181 5105
rect 233 5053 240 5105
rect 174 5041 190 5053
rect 224 5041 240 5053
rect 174 4989 181 5041
rect 233 4989 240 5041
rect 174 4977 190 4989
rect 224 4977 240 4989
rect 174 4925 181 4977
rect 233 4925 240 4977
rect 174 4924 240 4925
rect 174 4913 190 4924
rect 224 4913 240 4924
rect 174 4861 181 4913
rect 233 4861 240 4913
rect 174 4852 240 4861
rect 174 4849 190 4852
rect 224 4849 240 4852
rect 174 4797 181 4849
rect 233 4797 240 4849
rect 174 4744 240 4797
rect 174 4710 190 4744
rect 224 4710 240 4744
rect 174 4694 240 4710
rect 642 6364 688 6391
rect 642 6330 648 6364
rect 682 6330 688 6364
rect 642 6292 688 6330
rect 642 6258 648 6292
rect 682 6258 688 6292
rect 642 6220 688 6258
rect 642 6186 648 6220
rect 682 6186 688 6220
rect 642 6148 688 6186
rect 642 6114 648 6148
rect 682 6114 688 6148
rect 642 6076 688 6114
rect 642 6042 648 6076
rect 682 6042 688 6076
rect 642 6004 688 6042
rect 642 5970 648 6004
rect 682 5970 688 6004
rect 642 5932 688 5970
rect 642 5898 648 5932
rect 682 5898 688 5932
rect 642 5860 688 5898
rect 642 5826 648 5860
rect 682 5826 688 5860
rect 642 5788 688 5826
rect 642 5754 648 5788
rect 682 5754 688 5788
rect 642 5716 688 5754
rect 642 5682 648 5716
rect 682 5682 688 5716
rect 642 5644 688 5682
rect 642 5610 648 5644
rect 682 5610 688 5644
rect 642 5572 688 5610
rect 642 5538 648 5572
rect 682 5538 688 5572
rect 642 5500 688 5538
rect 642 5466 648 5500
rect 682 5466 688 5500
rect 642 5428 688 5466
rect 642 5394 648 5428
rect 682 5394 688 5428
rect 642 5356 688 5394
rect 642 5322 648 5356
rect 682 5322 688 5356
rect 642 5284 688 5322
rect 642 5250 648 5284
rect 682 5250 688 5284
rect 642 5212 688 5250
rect 642 5178 648 5212
rect 682 5178 688 5212
rect 642 5140 688 5178
rect 642 5106 648 5140
rect 682 5106 688 5140
rect 642 5068 688 5106
rect 642 5034 648 5068
rect 682 5034 688 5068
rect 642 4996 688 5034
rect 642 4962 648 4996
rect 682 4962 688 4996
rect 642 4924 688 4962
rect 642 4890 648 4924
rect 682 4890 688 4924
rect 642 4852 688 4890
rect 642 4818 648 4852
rect 682 4818 688 4852
rect 642 4648 688 4818
rect 1090 6385 1156 6438
rect 1090 6333 1097 6385
rect 1149 6333 1156 6385
rect 1090 6330 1106 6333
rect 1140 6330 1156 6333
rect 1090 6321 1156 6330
rect 1090 6269 1097 6321
rect 1149 6269 1156 6321
rect 1090 6258 1106 6269
rect 1140 6258 1156 6269
rect 1090 6257 1156 6258
rect 1090 6205 1097 6257
rect 1149 6205 1156 6257
rect 1090 6193 1106 6205
rect 1140 6193 1156 6205
rect 1090 6141 1097 6193
rect 1149 6141 1156 6193
rect 1090 6129 1106 6141
rect 1140 6129 1156 6141
rect 1090 6077 1097 6129
rect 1149 6077 1156 6129
rect 1090 6076 1156 6077
rect 1090 6065 1106 6076
rect 1140 6065 1156 6076
rect 1090 6013 1097 6065
rect 1149 6013 1156 6065
rect 1090 6004 1156 6013
rect 1090 6001 1106 6004
rect 1140 6001 1156 6004
rect 1090 5949 1097 6001
rect 1149 5949 1156 6001
rect 1090 5937 1156 5949
rect 1090 5885 1097 5937
rect 1149 5885 1156 5937
rect 1090 5873 1156 5885
rect 1090 5821 1097 5873
rect 1149 5821 1156 5873
rect 1090 5809 1156 5821
rect 1090 5757 1097 5809
rect 1149 5757 1156 5809
rect 1090 5754 1106 5757
rect 1140 5754 1156 5757
rect 1090 5745 1156 5754
rect 1090 5693 1097 5745
rect 1149 5693 1156 5745
rect 1090 5682 1106 5693
rect 1140 5682 1156 5693
rect 1090 5681 1156 5682
rect 1090 5629 1097 5681
rect 1149 5629 1156 5681
rect 1090 5617 1106 5629
rect 1140 5617 1156 5629
rect 1090 5565 1097 5617
rect 1149 5565 1156 5617
rect 1090 5553 1106 5565
rect 1140 5553 1156 5565
rect 1090 5501 1097 5553
rect 1149 5501 1156 5553
rect 1090 5500 1156 5501
rect 1090 5489 1106 5500
rect 1140 5489 1156 5500
rect 1090 5437 1097 5489
rect 1149 5437 1156 5489
rect 1090 5428 1156 5437
rect 1090 5425 1106 5428
rect 1140 5425 1156 5428
rect 1090 5373 1097 5425
rect 1149 5373 1156 5425
rect 1090 5361 1156 5373
rect 1090 5309 1097 5361
rect 1149 5309 1156 5361
rect 1090 5297 1156 5309
rect 1090 5245 1097 5297
rect 1149 5245 1156 5297
rect 1090 5233 1156 5245
rect 1090 5181 1097 5233
rect 1149 5181 1156 5233
rect 1090 5178 1106 5181
rect 1140 5178 1156 5181
rect 1090 5169 1156 5178
rect 1090 5117 1097 5169
rect 1149 5117 1156 5169
rect 1090 5106 1106 5117
rect 1140 5106 1156 5117
rect 1090 5105 1156 5106
rect 1090 5053 1097 5105
rect 1149 5053 1156 5105
rect 1090 5041 1106 5053
rect 1140 5041 1156 5053
rect 1090 4989 1097 5041
rect 1149 4989 1156 5041
rect 1090 4977 1106 4989
rect 1140 4977 1156 4989
rect 1090 4925 1097 4977
rect 1149 4925 1156 4977
rect 1090 4924 1156 4925
rect 1090 4913 1106 4924
rect 1140 4913 1156 4924
rect 1090 4861 1097 4913
rect 1149 4861 1156 4913
rect 1090 4852 1156 4861
rect 1090 4849 1106 4852
rect 1140 4849 1156 4852
rect 1090 4797 1097 4849
rect 1149 4797 1156 4849
rect 1090 4744 1156 4797
rect 1090 4710 1106 4744
rect 1140 4710 1156 4744
rect 1090 4694 1156 4710
rect 1206 6472 1372 6488
rect 1206 6438 1220 6472
rect 1254 6438 1326 6472
rect 1360 6438 1372 6472
rect 1206 6400 1372 6438
rect 1206 6366 1220 6400
rect 1254 6366 1326 6400
rect 1360 6366 1372 6400
rect 1206 6328 1372 6366
rect 1206 6294 1220 6328
rect 1254 6294 1326 6328
rect 1360 6294 1372 6328
rect 1206 6256 1372 6294
rect 1206 6222 1220 6256
rect 1254 6222 1326 6256
rect 1360 6222 1372 6256
rect 1206 6184 1372 6222
rect 1206 6150 1220 6184
rect 1254 6150 1326 6184
rect 1360 6150 1372 6184
rect 1206 6112 1372 6150
rect 1206 6078 1220 6112
rect 1254 6078 1326 6112
rect 1360 6078 1372 6112
rect 1206 6040 1372 6078
rect 1206 6006 1220 6040
rect 1254 6006 1326 6040
rect 1360 6006 1372 6040
rect 1206 5968 1372 6006
rect 1206 5934 1220 5968
rect 1254 5934 1326 5968
rect 1360 5934 1372 5968
rect 1206 5896 1372 5934
rect 1206 5862 1220 5896
rect 1254 5862 1326 5896
rect 1360 5862 1372 5896
rect 1206 5824 1372 5862
rect 1206 5790 1220 5824
rect 1254 5790 1326 5824
rect 1360 5790 1372 5824
rect 1206 5752 1372 5790
rect 1206 5718 1220 5752
rect 1254 5718 1326 5752
rect 1360 5718 1372 5752
rect 1206 5680 1372 5718
rect 1206 5646 1220 5680
rect 1254 5646 1326 5680
rect 1360 5646 1372 5680
rect 1206 5608 1372 5646
rect 1206 5574 1220 5608
rect 1254 5574 1326 5608
rect 1360 5574 1372 5608
rect 1206 5536 1372 5574
rect 1206 5502 1220 5536
rect 1254 5502 1326 5536
rect 1360 5502 1372 5536
rect 1206 5464 1372 5502
rect 1206 5430 1220 5464
rect 1254 5430 1326 5464
rect 1360 5430 1372 5464
rect 1206 5392 1372 5430
rect 1206 5358 1220 5392
rect 1254 5358 1326 5392
rect 1360 5358 1372 5392
rect 1206 5320 1372 5358
rect 1206 5286 1220 5320
rect 1254 5286 1326 5320
rect 1360 5286 1372 5320
rect 1206 5248 1372 5286
rect 1206 5214 1220 5248
rect 1254 5214 1326 5248
rect 1360 5214 1372 5248
rect 1206 5176 1372 5214
rect 1206 5142 1220 5176
rect 1254 5142 1326 5176
rect 1360 5142 1372 5176
rect 1206 5104 1372 5142
rect 1206 5070 1220 5104
rect 1254 5070 1326 5104
rect 1360 5070 1372 5104
rect 1206 5032 1372 5070
rect 1206 4998 1220 5032
rect 1254 4998 1326 5032
rect 1360 4998 1372 5032
rect 1206 4960 1372 4998
rect 1206 4926 1220 4960
rect 1254 4926 1326 4960
rect 1360 4926 1372 4960
rect 1206 4888 1372 4926
rect 1206 4854 1220 4888
rect 1254 4854 1326 4888
rect 1360 4854 1372 4888
rect 1206 4816 1372 4854
rect 1206 4782 1220 4816
rect 1254 4782 1326 4816
rect 1360 4782 1372 4816
rect 1206 4744 1372 4782
rect 1206 4710 1220 4744
rect 1254 4710 1326 4744
rect 1360 4710 1372 4744
rect 1206 4684 1372 4710
rect 1424 6472 1490 6488
rect 1424 6438 1440 6472
rect 1474 6438 1490 6472
rect 1424 6385 1490 6438
rect 1424 6333 1431 6385
rect 1483 6333 1490 6385
rect 1424 6321 1490 6333
rect 1424 6269 1431 6321
rect 1483 6269 1490 6321
rect 1424 6257 1490 6269
rect 1424 6205 1431 6257
rect 1483 6205 1490 6257
rect 1424 6193 1490 6205
rect 1424 6141 1431 6193
rect 1483 6141 1490 6193
rect 1424 6129 1490 6141
rect 1424 6077 1431 6129
rect 1483 6077 1490 6129
rect 1424 6065 1490 6077
rect 1424 6013 1431 6065
rect 1483 6013 1490 6065
rect 1424 6001 1490 6013
rect 1424 5949 1431 6001
rect 1483 5949 1490 6001
rect 1424 5937 1490 5949
rect 1424 5885 1431 5937
rect 1483 5885 1490 5937
rect 1424 5873 1490 5885
rect 1424 5821 1431 5873
rect 1483 5821 1490 5873
rect 1424 5809 1490 5821
rect 1424 5757 1431 5809
rect 1483 5757 1490 5809
rect 1424 5745 1490 5757
rect 1424 5693 1431 5745
rect 1483 5693 1490 5745
rect 1424 5681 1490 5693
rect 1424 5629 1431 5681
rect 1483 5629 1490 5681
rect 1424 5617 1490 5629
rect 1424 5565 1431 5617
rect 1483 5565 1490 5617
rect 1424 5553 1490 5565
rect 1424 5501 1431 5553
rect 1483 5501 1490 5553
rect 1424 5489 1490 5501
rect 1424 5437 1431 5489
rect 1483 5437 1490 5489
rect 1424 5425 1490 5437
rect 1424 5373 1431 5425
rect 1483 5373 1490 5425
rect 1424 5361 1490 5373
rect 1424 5309 1431 5361
rect 1483 5309 1490 5361
rect 1424 5297 1490 5309
rect 1424 5245 1431 5297
rect 1483 5245 1490 5297
rect 1424 5233 1490 5245
rect 1424 5181 1431 5233
rect 1483 5181 1490 5233
rect 1424 5169 1490 5181
rect 1424 5117 1431 5169
rect 1483 5117 1490 5169
rect 1424 5105 1490 5117
rect 1424 5053 1431 5105
rect 1483 5053 1490 5105
rect 1424 5041 1490 5053
rect 1424 4989 1431 5041
rect 1483 4989 1490 5041
rect 1424 4977 1490 4989
rect 1424 4925 1431 4977
rect 1483 4925 1490 4977
rect 1424 4913 1490 4925
rect 1424 4861 1431 4913
rect 1483 4861 1490 4913
rect 1424 4849 1490 4861
rect 1424 4797 1431 4849
rect 1483 4797 1490 4849
rect 2340 6472 2406 6488
rect 2340 6438 2356 6472
rect 2390 6438 2406 6472
rect 2340 6385 2406 6438
rect 2340 6333 2347 6385
rect 2399 6333 2406 6385
rect 2340 6321 2406 6333
rect 2340 6269 2347 6321
rect 2399 6269 2406 6321
rect 2340 6257 2406 6269
rect 2340 6205 2347 6257
rect 2399 6205 2406 6257
rect 2340 6193 2406 6205
rect 2340 6141 2347 6193
rect 2399 6141 2406 6193
rect 2340 6129 2406 6141
rect 2340 6077 2347 6129
rect 2399 6077 2406 6129
rect 2340 6065 2406 6077
rect 2340 6013 2347 6065
rect 2399 6013 2406 6065
rect 2340 6001 2406 6013
rect 2340 5949 2347 6001
rect 2399 5949 2406 6001
rect 2340 5937 2406 5949
rect 2340 5885 2347 5937
rect 2399 5885 2406 5937
rect 2340 5873 2406 5885
rect 2340 5821 2347 5873
rect 2399 5821 2406 5873
rect 2340 5809 2406 5821
rect 2340 5757 2347 5809
rect 2399 5757 2406 5809
rect 2340 5745 2406 5757
rect 2340 5693 2347 5745
rect 2399 5693 2406 5745
rect 2340 5681 2406 5693
rect 2340 5629 2347 5681
rect 2399 5629 2406 5681
rect 2340 5617 2406 5629
rect 2340 5565 2347 5617
rect 2399 5565 2406 5617
rect 2340 5553 2406 5565
rect 2340 5501 2347 5553
rect 2399 5501 2406 5553
rect 2340 5489 2406 5501
rect 2340 5437 2347 5489
rect 2399 5437 2406 5489
rect 2340 5425 2406 5437
rect 2340 5373 2347 5425
rect 2399 5373 2406 5425
rect 2340 5361 2406 5373
rect 2340 5309 2347 5361
rect 2399 5309 2406 5361
rect 2340 5297 2406 5309
rect 2340 5245 2347 5297
rect 2399 5245 2406 5297
rect 2340 5233 2406 5245
rect 2340 5181 2347 5233
rect 2399 5181 2406 5233
rect 2340 5169 2406 5181
rect 2340 5117 2347 5169
rect 2399 5117 2406 5169
rect 2340 5105 2406 5117
rect 2340 5053 2347 5105
rect 2399 5053 2406 5105
rect 2340 5041 2406 5053
rect 2340 4989 2347 5041
rect 2399 4989 2406 5041
rect 2340 4977 2406 4989
rect 2340 4925 2347 4977
rect 2399 4925 2406 4977
rect 2340 4913 2406 4925
rect 2340 4861 2347 4913
rect 2399 4861 2406 4913
rect 2340 4849 2406 4861
rect 1424 4744 1490 4797
rect 1424 4710 1440 4744
rect 1474 4710 1490 4744
rect 1424 4694 1490 4710
rect -1276 4642 1232 4648
rect 1892 4646 1938 4807
rect 2340 4797 2347 4849
rect 2399 4797 2406 4849
rect 3256 6472 3322 6488
rect 3256 6438 3272 6472
rect 3306 6438 3322 6472
rect 3256 6385 3322 6438
rect 3256 6333 3263 6385
rect 3315 6333 3322 6385
rect 3256 6321 3322 6333
rect 3256 6269 3263 6321
rect 3315 6269 3322 6321
rect 3256 6257 3322 6269
rect 3256 6205 3263 6257
rect 3315 6205 3322 6257
rect 3256 6193 3322 6205
rect 3256 6141 3263 6193
rect 3315 6141 3322 6193
rect 3256 6129 3322 6141
rect 3256 6077 3263 6129
rect 3315 6077 3322 6129
rect 3256 6065 3322 6077
rect 3256 6013 3263 6065
rect 3315 6013 3322 6065
rect 3256 6001 3322 6013
rect 3256 5949 3263 6001
rect 3315 5949 3322 6001
rect 3256 5937 3322 5949
rect 3256 5885 3263 5937
rect 3315 5885 3322 5937
rect 3256 5873 3322 5885
rect 3256 5821 3263 5873
rect 3315 5821 3322 5873
rect 3256 5809 3322 5821
rect 3256 5757 3263 5809
rect 3315 5757 3322 5809
rect 3256 5745 3322 5757
rect 3256 5693 3263 5745
rect 3315 5693 3322 5745
rect 3256 5681 3322 5693
rect 3256 5629 3263 5681
rect 3315 5629 3322 5681
rect 3256 5617 3322 5629
rect 3256 5565 3263 5617
rect 3315 5565 3322 5617
rect 3256 5553 3322 5565
rect 3256 5501 3263 5553
rect 3315 5501 3322 5553
rect 3256 5489 3322 5501
rect 3256 5437 3263 5489
rect 3315 5437 3322 5489
rect 3256 5425 3322 5437
rect 3256 5373 3263 5425
rect 3315 5373 3322 5425
rect 3256 5361 3322 5373
rect 3256 5309 3263 5361
rect 3315 5309 3322 5361
rect 3256 5297 3322 5309
rect 3256 5245 3263 5297
rect 3315 5245 3322 5297
rect 3256 5233 3322 5245
rect 3256 5181 3263 5233
rect 3315 5181 3322 5233
rect 3256 5169 3322 5181
rect 3256 5117 3263 5169
rect 3315 5117 3322 5169
rect 3256 5105 3322 5117
rect 3256 5053 3263 5105
rect 3315 5053 3322 5105
rect 3256 5041 3322 5053
rect 3256 4989 3263 5041
rect 3315 4989 3322 5041
rect 3256 4977 3322 4989
rect 3256 4925 3263 4977
rect 3315 4925 3322 4977
rect 3256 4913 3322 4925
rect 3256 4861 3263 4913
rect 3315 4861 3322 4913
rect 3256 4849 3322 4861
rect 2340 4744 2406 4797
rect 2340 4710 2356 4744
rect 2390 4710 2406 4744
rect 2340 4694 2406 4710
rect 2808 4646 2854 4807
rect 3256 4797 3263 4849
rect 3315 4797 3322 4849
rect 3256 4744 3322 4797
rect 3256 4710 3272 4744
rect 3306 4710 3322 4744
rect 3256 4694 3322 4710
rect 3724 4646 3770 4807
rect -1276 4608 -1263 4642
rect -1229 4608 -1191 4642
rect -1157 4608 -1119 4642
rect -1085 4608 -1047 4642
rect -1013 4608 -975 4642
rect -941 4608 -903 4642
rect -869 4608 -831 4642
rect -797 4608 -759 4642
rect -725 4608 -687 4642
rect -653 4608 -615 4642
rect -581 4608 -543 4642
rect -509 4608 -471 4642
rect -437 4608 -399 4642
rect -365 4608 -327 4642
rect -293 4608 -255 4642
rect -221 4608 -183 4642
rect -149 4608 -111 4642
rect -77 4608 -39 4642
rect -5 4608 33 4642
rect 67 4608 105 4642
rect 139 4608 177 4642
rect 211 4608 249 4642
rect 283 4608 321 4642
rect 355 4608 393 4642
rect 427 4608 465 4642
rect 499 4608 537 4642
rect 571 4608 609 4642
rect 643 4608 681 4642
rect 715 4608 753 4642
rect 787 4608 825 4642
rect 859 4608 897 4642
rect 931 4608 969 4642
rect 1003 4608 1041 4642
rect 1075 4608 1113 4642
rect 1147 4608 1185 4642
rect 1219 4608 1232 4642
rect -1276 4536 1232 4608
rect 1348 4540 3856 4604
rect -1276 4502 -1263 4536
rect -1229 4502 -1191 4536
rect -1157 4502 -1119 4536
rect -1085 4502 -1047 4536
rect -1013 4502 -975 4536
rect -941 4502 -903 4536
rect -869 4502 -831 4536
rect -797 4502 -759 4536
rect -725 4502 -687 4536
rect -653 4502 -615 4536
rect -581 4502 -543 4536
rect -509 4502 -471 4536
rect -437 4502 -399 4536
rect -365 4502 -327 4536
rect -293 4502 -255 4536
rect -221 4502 -183 4536
rect -149 4502 -111 4536
rect -77 4502 -39 4536
rect -5 4502 33 4536
rect 67 4502 105 4536
rect 139 4502 177 4536
rect 211 4502 249 4536
rect 283 4502 321 4536
rect 355 4502 393 4536
rect 427 4502 465 4536
rect 499 4502 537 4536
rect 571 4502 609 4536
rect 643 4502 681 4536
rect 715 4502 753 4536
rect 787 4502 825 4536
rect 859 4502 897 4536
rect 931 4502 969 4536
rect 1003 4502 1041 4536
rect 1075 4502 1113 4536
rect 1147 4502 1185 4536
rect 1219 4502 1232 4536
rect -1276 4496 1232 4502
rect -1190 4326 -1144 4496
rect -1190 4292 -1184 4326
rect -1150 4292 -1144 4326
rect -1190 4254 -1144 4292
rect -1190 4220 -1184 4254
rect -1150 4220 -1144 4254
rect -1190 4182 -1144 4220
rect -1190 4148 -1184 4182
rect -1150 4148 -1144 4182
rect -1190 4110 -1144 4148
rect -1190 4076 -1184 4110
rect -1150 4076 -1144 4110
rect -1190 4038 -1144 4076
rect -1190 4004 -1184 4038
rect -1150 4004 -1144 4038
rect -1190 3966 -1144 4004
rect -1190 3932 -1184 3966
rect -1150 3932 -1144 3966
rect -1190 3894 -1144 3932
rect -1190 3860 -1184 3894
rect -1150 3860 -1144 3894
rect -1190 3822 -1144 3860
rect -1190 3788 -1184 3822
rect -1150 3788 -1144 3822
rect -1190 3750 -1144 3788
rect -1190 3716 -1184 3750
rect -1150 3716 -1144 3750
rect -1190 3678 -1144 3716
rect -1190 3644 -1184 3678
rect -1150 3644 -1144 3678
rect -1190 3606 -1144 3644
rect -1190 3572 -1184 3606
rect -1150 3572 -1144 3606
rect -1190 3534 -1144 3572
rect -1190 3500 -1184 3534
rect -1150 3500 -1144 3534
rect -1190 3462 -1144 3500
rect -1190 3428 -1184 3462
rect -1150 3428 -1144 3462
rect -1190 3390 -1144 3428
rect -1190 3356 -1184 3390
rect -1150 3356 -1144 3390
rect -1190 3318 -1144 3356
rect -1190 3284 -1184 3318
rect -1150 3284 -1144 3318
rect -1190 3246 -1144 3284
rect -1190 3212 -1184 3246
rect -1150 3212 -1144 3246
rect -1190 3174 -1144 3212
rect -1190 3140 -1184 3174
rect -1150 3140 -1144 3174
rect -1190 3102 -1144 3140
rect -1190 3068 -1184 3102
rect -1150 3068 -1144 3102
rect -1190 3030 -1144 3068
rect -1190 2996 -1184 3030
rect -1150 2996 -1144 3030
rect -1190 2958 -1144 2996
rect -1190 2924 -1184 2958
rect -1150 2924 -1144 2958
rect -1190 2886 -1144 2924
rect -1190 2852 -1184 2886
rect -1150 2852 -1144 2886
rect -1190 2814 -1144 2852
rect -1190 2780 -1184 2814
rect -1150 2780 -1144 2814
rect -1190 2753 -1144 2780
rect -742 4347 -676 4360
rect -742 4295 -735 4347
rect -683 4295 -676 4347
rect -742 4292 -726 4295
rect -692 4292 -676 4295
rect -742 4283 -676 4292
rect -742 4231 -735 4283
rect -683 4231 -676 4283
rect -742 4220 -726 4231
rect -692 4220 -676 4231
rect -742 4219 -676 4220
rect -742 4167 -735 4219
rect -683 4167 -676 4219
rect -742 4155 -726 4167
rect -692 4155 -676 4167
rect -742 4103 -735 4155
rect -683 4103 -676 4155
rect -742 4091 -726 4103
rect -692 4091 -676 4103
rect -742 4039 -735 4091
rect -683 4039 -676 4091
rect -742 4038 -676 4039
rect -742 4027 -726 4038
rect -692 4027 -676 4038
rect -742 3975 -735 4027
rect -683 3975 -676 4027
rect -742 3966 -676 3975
rect -742 3963 -726 3966
rect -692 3963 -676 3966
rect -742 3911 -735 3963
rect -683 3911 -676 3963
rect -742 3899 -676 3911
rect -742 3847 -735 3899
rect -683 3847 -676 3899
rect -742 3835 -676 3847
rect -742 3783 -735 3835
rect -683 3783 -676 3835
rect -742 3771 -676 3783
rect -742 3719 -735 3771
rect -683 3719 -676 3771
rect -742 3716 -726 3719
rect -692 3716 -676 3719
rect -742 3707 -676 3716
rect -742 3655 -735 3707
rect -683 3655 -676 3707
rect -742 3644 -726 3655
rect -692 3644 -676 3655
rect -742 3643 -676 3644
rect -742 3591 -735 3643
rect -683 3591 -676 3643
rect -742 3579 -726 3591
rect -692 3579 -676 3591
rect -742 3527 -735 3579
rect -683 3527 -676 3579
rect -742 3515 -726 3527
rect -692 3515 -676 3527
rect -742 3463 -735 3515
rect -683 3463 -676 3515
rect -742 3462 -676 3463
rect -742 3451 -726 3462
rect -692 3451 -676 3462
rect -742 3399 -735 3451
rect -683 3399 -676 3451
rect -742 3390 -676 3399
rect -742 3387 -726 3390
rect -692 3387 -676 3390
rect -742 3335 -735 3387
rect -683 3335 -676 3387
rect -742 3323 -676 3335
rect -742 3271 -735 3323
rect -683 3271 -676 3323
rect -742 3259 -676 3271
rect -742 3207 -735 3259
rect -683 3207 -676 3259
rect -742 3195 -676 3207
rect -742 3143 -735 3195
rect -683 3143 -676 3195
rect -742 3140 -726 3143
rect -692 3140 -676 3143
rect -742 3131 -676 3140
rect -742 3079 -735 3131
rect -683 3079 -676 3131
rect -742 3068 -726 3079
rect -692 3068 -676 3079
rect -742 3067 -676 3068
rect -742 3015 -735 3067
rect -683 3015 -676 3067
rect -742 3003 -726 3015
rect -692 3003 -676 3015
rect -742 2951 -735 3003
rect -683 2951 -676 3003
rect -742 2939 -726 2951
rect -692 2939 -676 2951
rect -742 2887 -735 2939
rect -683 2887 -676 2939
rect -742 2886 -676 2887
rect -742 2875 -726 2886
rect -692 2875 -676 2886
rect -742 2823 -735 2875
rect -683 2823 -676 2875
rect -742 2814 -676 2823
rect -742 2811 -726 2814
rect -692 2811 -676 2814
rect -742 2759 -735 2811
rect -683 2759 -676 2811
rect -742 2746 -676 2759
rect -274 4326 -228 4496
rect -274 4292 -268 4326
rect -234 4292 -228 4326
rect -274 4254 -228 4292
rect -274 4220 -268 4254
rect -234 4220 -228 4254
rect -274 4182 -228 4220
rect -274 4148 -268 4182
rect -234 4148 -228 4182
rect -274 4110 -228 4148
rect -274 4076 -268 4110
rect -234 4076 -228 4110
rect -274 4038 -228 4076
rect -274 4004 -268 4038
rect -234 4004 -228 4038
rect -274 3966 -228 4004
rect -274 3932 -268 3966
rect -234 3932 -228 3966
rect -274 3894 -228 3932
rect -274 3860 -268 3894
rect -234 3860 -228 3894
rect -274 3822 -228 3860
rect -274 3788 -268 3822
rect -234 3788 -228 3822
rect -274 3750 -228 3788
rect -274 3716 -268 3750
rect -234 3716 -228 3750
rect -274 3678 -228 3716
rect -274 3644 -268 3678
rect -234 3644 -228 3678
rect -274 3606 -228 3644
rect -274 3572 -268 3606
rect -234 3572 -228 3606
rect -274 3534 -228 3572
rect -274 3500 -268 3534
rect -234 3500 -228 3534
rect -274 3462 -228 3500
rect -274 3428 -268 3462
rect -234 3428 -228 3462
rect -274 3390 -228 3428
rect -274 3356 -268 3390
rect -234 3356 -228 3390
rect -274 3318 -228 3356
rect -274 3284 -268 3318
rect -234 3284 -228 3318
rect -274 3246 -228 3284
rect -274 3212 -268 3246
rect -234 3212 -228 3246
rect -274 3174 -228 3212
rect -274 3140 -268 3174
rect -234 3140 -228 3174
rect -274 3102 -228 3140
rect -274 3068 -268 3102
rect -234 3068 -228 3102
rect -274 3030 -228 3068
rect -274 2996 -268 3030
rect -234 2996 -228 3030
rect -274 2958 -228 2996
rect -274 2924 -268 2958
rect -234 2924 -228 2958
rect -274 2886 -228 2924
rect -274 2852 -268 2886
rect -234 2852 -228 2886
rect -274 2814 -228 2852
rect -274 2780 -268 2814
rect -234 2780 -228 2814
rect -274 2753 -228 2780
rect 174 4347 240 4360
rect 174 4295 181 4347
rect 233 4295 240 4347
rect 174 4292 190 4295
rect 224 4292 240 4295
rect 174 4283 240 4292
rect 174 4231 181 4283
rect 233 4231 240 4283
rect 174 4220 190 4231
rect 224 4220 240 4231
rect 174 4219 240 4220
rect 174 4167 181 4219
rect 233 4167 240 4219
rect 174 4155 190 4167
rect 224 4155 240 4167
rect 174 4103 181 4155
rect 233 4103 240 4155
rect 174 4091 190 4103
rect 224 4091 240 4103
rect 174 4039 181 4091
rect 233 4039 240 4091
rect 174 4038 240 4039
rect 174 4027 190 4038
rect 224 4027 240 4038
rect 174 3975 181 4027
rect 233 3975 240 4027
rect 174 3966 240 3975
rect 174 3963 190 3966
rect 224 3963 240 3966
rect 174 3911 181 3963
rect 233 3911 240 3963
rect 174 3899 240 3911
rect 174 3847 181 3899
rect 233 3847 240 3899
rect 174 3835 240 3847
rect 174 3783 181 3835
rect 233 3783 240 3835
rect 174 3771 240 3783
rect 174 3719 181 3771
rect 233 3719 240 3771
rect 174 3716 190 3719
rect 224 3716 240 3719
rect 174 3707 240 3716
rect 174 3655 181 3707
rect 233 3655 240 3707
rect 174 3644 190 3655
rect 224 3644 240 3655
rect 174 3643 240 3644
rect 174 3591 181 3643
rect 233 3591 240 3643
rect 174 3579 190 3591
rect 224 3579 240 3591
rect 174 3527 181 3579
rect 233 3527 240 3579
rect 174 3515 190 3527
rect 224 3515 240 3527
rect 174 3463 181 3515
rect 233 3463 240 3515
rect 174 3462 240 3463
rect 174 3451 190 3462
rect 224 3451 240 3462
rect 174 3399 181 3451
rect 233 3399 240 3451
rect 174 3390 240 3399
rect 174 3387 190 3390
rect 224 3387 240 3390
rect 174 3335 181 3387
rect 233 3335 240 3387
rect 174 3323 240 3335
rect 174 3271 181 3323
rect 233 3271 240 3323
rect 174 3259 240 3271
rect 174 3207 181 3259
rect 233 3207 240 3259
rect 174 3195 240 3207
rect 174 3143 181 3195
rect 233 3143 240 3195
rect 174 3140 190 3143
rect 224 3140 240 3143
rect 174 3131 240 3140
rect 174 3079 181 3131
rect 233 3079 240 3131
rect 174 3068 190 3079
rect 224 3068 240 3079
rect 174 3067 240 3068
rect 174 3015 181 3067
rect 233 3015 240 3067
rect 174 3003 190 3015
rect 224 3003 240 3015
rect 174 2951 181 3003
rect 233 2951 240 3003
rect 174 2939 190 2951
rect 224 2939 240 2951
rect 174 2887 181 2939
rect 233 2887 240 2939
rect 174 2886 240 2887
rect 174 2875 190 2886
rect 224 2875 240 2886
rect 174 2823 181 2875
rect 233 2823 240 2875
rect 174 2814 240 2823
rect 174 2811 190 2814
rect 224 2811 240 2814
rect 174 2759 181 2811
rect 233 2759 240 2811
rect 174 2746 240 2759
rect 642 4326 688 4496
rect 1208 4434 1374 4456
rect 1208 4400 1220 4434
rect 1254 4400 1326 4434
rect 1360 4400 1374 4434
rect 1208 4362 1374 4400
rect 642 4292 648 4326
rect 682 4292 688 4326
rect 642 4254 688 4292
rect 642 4220 648 4254
rect 682 4220 688 4254
rect 642 4182 688 4220
rect 642 4148 648 4182
rect 682 4148 688 4182
rect 642 4110 688 4148
rect 642 4076 648 4110
rect 682 4076 688 4110
rect 642 4038 688 4076
rect 642 4004 648 4038
rect 682 4004 688 4038
rect 642 3966 688 4004
rect 642 3932 648 3966
rect 682 3932 688 3966
rect 642 3894 688 3932
rect 642 3860 648 3894
rect 682 3860 688 3894
rect 642 3822 688 3860
rect 642 3788 648 3822
rect 682 3788 688 3822
rect 642 3750 688 3788
rect 642 3716 648 3750
rect 682 3716 688 3750
rect 642 3678 688 3716
rect 642 3644 648 3678
rect 682 3644 688 3678
rect 642 3606 688 3644
rect 642 3572 648 3606
rect 682 3572 688 3606
rect 642 3534 688 3572
rect 642 3500 648 3534
rect 682 3500 688 3534
rect 642 3462 688 3500
rect 642 3428 648 3462
rect 682 3428 688 3462
rect 642 3390 688 3428
rect 642 3356 648 3390
rect 682 3356 688 3390
rect 642 3318 688 3356
rect 642 3284 648 3318
rect 682 3284 688 3318
rect 642 3246 688 3284
rect 642 3212 648 3246
rect 682 3212 688 3246
rect 642 3174 688 3212
rect 642 3140 648 3174
rect 682 3140 688 3174
rect 642 3102 688 3140
rect 642 3068 648 3102
rect 682 3068 688 3102
rect 642 3030 688 3068
rect 642 2996 648 3030
rect 682 2996 688 3030
rect 642 2958 688 2996
rect 642 2924 648 2958
rect 682 2924 688 2958
rect 642 2886 688 2924
rect 642 2852 648 2886
rect 682 2852 688 2886
rect 642 2814 688 2852
rect 642 2780 648 2814
rect 682 2780 688 2814
rect 642 2753 688 2780
rect 1090 4347 1156 4360
rect 1090 4295 1097 4347
rect 1149 4295 1156 4347
rect 1090 4292 1106 4295
rect 1140 4292 1156 4295
rect 1090 4283 1156 4292
rect 1090 4231 1097 4283
rect 1149 4231 1156 4283
rect 1090 4220 1106 4231
rect 1140 4220 1156 4231
rect 1090 4219 1156 4220
rect 1090 4167 1097 4219
rect 1149 4167 1156 4219
rect 1090 4155 1106 4167
rect 1140 4155 1156 4167
rect 1090 4103 1097 4155
rect 1149 4103 1156 4155
rect 1090 4091 1106 4103
rect 1140 4091 1156 4103
rect 1090 4039 1097 4091
rect 1149 4039 1156 4091
rect 1090 4038 1156 4039
rect 1090 4027 1106 4038
rect 1140 4027 1156 4038
rect 1090 3975 1097 4027
rect 1149 3975 1156 4027
rect 1090 3966 1156 3975
rect 1090 3963 1106 3966
rect 1140 3963 1156 3966
rect 1090 3911 1097 3963
rect 1149 3911 1156 3963
rect 1090 3899 1156 3911
rect 1090 3847 1097 3899
rect 1149 3847 1156 3899
rect 1090 3835 1156 3847
rect 1090 3783 1097 3835
rect 1149 3783 1156 3835
rect 1090 3771 1156 3783
rect 1090 3719 1097 3771
rect 1149 3719 1156 3771
rect 1090 3716 1106 3719
rect 1140 3716 1156 3719
rect 1090 3707 1156 3716
rect 1090 3655 1097 3707
rect 1149 3655 1156 3707
rect 1090 3644 1106 3655
rect 1140 3644 1156 3655
rect 1090 3643 1156 3644
rect 1090 3591 1097 3643
rect 1149 3591 1156 3643
rect 1090 3579 1106 3591
rect 1140 3579 1156 3591
rect 1090 3527 1097 3579
rect 1149 3527 1156 3579
rect 1090 3515 1106 3527
rect 1140 3515 1156 3527
rect 1090 3463 1097 3515
rect 1149 3463 1156 3515
rect 1090 3462 1156 3463
rect 1090 3451 1106 3462
rect 1140 3451 1156 3462
rect 1090 3399 1097 3451
rect 1149 3399 1156 3451
rect 1090 3390 1156 3399
rect 1090 3387 1106 3390
rect 1140 3387 1156 3390
rect 1090 3335 1097 3387
rect 1149 3335 1156 3387
rect 1090 3323 1156 3335
rect 1090 3271 1097 3323
rect 1149 3271 1156 3323
rect 1090 3259 1156 3271
rect 1090 3207 1097 3259
rect 1149 3207 1156 3259
rect 1090 3195 1156 3207
rect 1090 3143 1097 3195
rect 1149 3143 1156 3195
rect 1090 3140 1106 3143
rect 1140 3140 1156 3143
rect 1090 3131 1156 3140
rect 1090 3079 1097 3131
rect 1149 3079 1156 3131
rect 1090 3068 1106 3079
rect 1140 3068 1156 3079
rect 1090 3067 1156 3068
rect 1090 3015 1097 3067
rect 1149 3015 1156 3067
rect 1090 3003 1106 3015
rect 1140 3003 1156 3015
rect 1090 2951 1097 3003
rect 1149 2951 1156 3003
rect 1090 2939 1106 2951
rect 1140 2939 1156 2951
rect 1090 2887 1097 2939
rect 1149 2887 1156 2939
rect 1090 2886 1156 2887
rect 1090 2875 1106 2886
rect 1140 2875 1156 2886
rect 1090 2823 1097 2875
rect 1149 2823 1156 2875
rect 1090 2814 1156 2823
rect 1090 2811 1106 2814
rect 1140 2811 1156 2814
rect 1090 2759 1097 2811
rect 1149 2759 1156 2811
rect 1090 2746 1156 2759
rect 1208 4328 1220 4362
rect 1254 4328 1326 4362
rect 1360 4328 1374 4362
rect 1208 4290 1374 4328
rect 1208 4256 1220 4290
rect 1254 4256 1326 4290
rect 1360 4256 1374 4290
rect 1208 4218 1374 4256
rect 1208 4184 1220 4218
rect 1254 4184 1326 4218
rect 1360 4184 1374 4218
rect 1208 4146 1374 4184
rect 1208 4112 1220 4146
rect 1254 4112 1326 4146
rect 1360 4112 1374 4146
rect 1208 4074 1374 4112
rect 1208 4040 1220 4074
rect 1254 4040 1326 4074
rect 1360 4040 1374 4074
rect 1208 4002 1374 4040
rect 1208 3968 1220 4002
rect 1254 3968 1326 4002
rect 1360 3968 1374 4002
rect 1208 3930 1374 3968
rect 1208 3896 1220 3930
rect 1254 3896 1326 3930
rect 1360 3896 1374 3930
rect 1208 3858 1374 3896
rect 1208 3824 1220 3858
rect 1254 3824 1326 3858
rect 1360 3824 1374 3858
rect 1208 3786 1374 3824
rect 1208 3752 1220 3786
rect 1254 3752 1326 3786
rect 1360 3752 1374 3786
rect 1208 3714 1374 3752
rect 1208 3680 1220 3714
rect 1254 3680 1326 3714
rect 1360 3680 1374 3714
rect 1208 3642 1374 3680
rect 1208 3608 1220 3642
rect 1254 3608 1326 3642
rect 1360 3608 1374 3642
rect 1208 3570 1374 3608
rect 1208 3536 1220 3570
rect 1254 3536 1326 3570
rect 1360 3536 1374 3570
rect 1208 3498 1374 3536
rect 1208 3464 1220 3498
rect 1254 3464 1326 3498
rect 1360 3464 1374 3498
rect 1208 3426 1374 3464
rect 1208 3392 1220 3426
rect 1254 3392 1326 3426
rect 1360 3392 1374 3426
rect 1208 3354 1374 3392
rect 1208 3320 1220 3354
rect 1254 3320 1326 3354
rect 1360 3320 1374 3354
rect 1208 3282 1374 3320
rect 1208 3248 1220 3282
rect 1254 3248 1326 3282
rect 1360 3248 1374 3282
rect 1208 3210 1374 3248
rect 1208 3176 1220 3210
rect 1254 3176 1326 3210
rect 1360 3176 1374 3210
rect 1208 3138 1374 3176
rect 1208 3104 1220 3138
rect 1254 3104 1326 3138
rect 1360 3104 1374 3138
rect 1208 3066 1374 3104
rect 1208 3032 1220 3066
rect 1254 3032 1326 3066
rect 1360 3032 1374 3066
rect 1208 2994 1374 3032
rect 1208 2960 1220 2994
rect 1254 2960 1326 2994
rect 1360 2960 1374 2994
rect 1208 2922 1374 2960
rect 1208 2888 1220 2922
rect 1254 2888 1326 2922
rect 1360 2888 1374 2922
rect 1208 2850 1374 2888
rect 1208 2816 1220 2850
rect 1254 2816 1326 2850
rect 1360 2816 1374 2850
rect 1208 2778 1374 2816
rect 1208 2744 1220 2778
rect 1254 2744 1326 2778
rect 1360 2744 1374 2778
rect 1424 4347 1490 4360
rect 1892 4352 1938 4502
rect 1424 4295 1431 4347
rect 1483 4295 1490 4347
rect 1424 4283 1490 4295
rect 1424 4231 1431 4283
rect 1483 4231 1490 4283
rect 1424 4219 1490 4231
rect 1424 4167 1431 4219
rect 1483 4167 1490 4219
rect 1424 4155 1490 4167
rect 1424 4103 1431 4155
rect 1483 4103 1490 4155
rect 1424 4091 1490 4103
rect 1424 4039 1431 4091
rect 1483 4039 1490 4091
rect 1424 4027 1490 4039
rect 1424 3975 1431 4027
rect 1483 3975 1490 4027
rect 1424 3963 1490 3975
rect 1424 3911 1431 3963
rect 1483 3911 1490 3963
rect 1424 3899 1490 3911
rect 1424 3847 1431 3899
rect 1483 3847 1490 3899
rect 1424 3835 1490 3847
rect 1424 3783 1431 3835
rect 1483 3783 1490 3835
rect 1424 3771 1490 3783
rect 1424 3719 1431 3771
rect 1483 3719 1490 3771
rect 1424 3707 1490 3719
rect 1424 3655 1431 3707
rect 1483 3655 1490 3707
rect 1424 3643 1490 3655
rect 1424 3591 1431 3643
rect 1483 3591 1490 3643
rect 1424 3579 1490 3591
rect 1424 3527 1431 3579
rect 1483 3527 1490 3579
rect 1424 3515 1490 3527
rect 1424 3463 1431 3515
rect 1483 3463 1490 3515
rect 1424 3451 1490 3463
rect 1424 3399 1431 3451
rect 1483 3399 1490 3451
rect 1424 3387 1490 3399
rect 1424 3335 1431 3387
rect 1483 3335 1490 3387
rect 1424 3323 1490 3335
rect 1424 3271 1431 3323
rect 1483 3271 1490 3323
rect 1424 3259 1490 3271
rect 1424 3207 1431 3259
rect 1483 3207 1490 3259
rect 1424 3195 1490 3207
rect 1424 3143 1431 3195
rect 1483 3143 1490 3195
rect 1424 3131 1490 3143
rect 1424 3079 1431 3131
rect 1483 3079 1490 3131
rect 1424 3067 1490 3079
rect 1424 3015 1431 3067
rect 1483 3015 1490 3067
rect 1424 3003 1490 3015
rect 1424 2951 1431 3003
rect 1483 2951 1490 3003
rect 1424 2939 1490 2951
rect 1424 2887 1431 2939
rect 1483 2887 1490 2939
rect 1424 2875 1490 2887
rect 1424 2823 1431 2875
rect 1483 2823 1490 2875
rect 1424 2811 1490 2823
rect 1424 2759 1431 2811
rect 1483 2759 1490 2811
rect 1424 2746 1490 2759
rect 2340 4347 2406 4360
rect 2808 4352 2854 4502
rect 2340 4295 2347 4347
rect 2399 4295 2406 4347
rect 2340 4283 2406 4295
rect 2340 4231 2347 4283
rect 2399 4231 2406 4283
rect 2340 4219 2406 4231
rect 2340 4167 2347 4219
rect 2399 4167 2406 4219
rect 2340 4155 2406 4167
rect 2340 4103 2347 4155
rect 2399 4103 2406 4155
rect 2340 4091 2406 4103
rect 2340 4039 2347 4091
rect 2399 4039 2406 4091
rect 2340 4027 2406 4039
rect 2340 3975 2347 4027
rect 2399 3975 2406 4027
rect 2340 3963 2406 3975
rect 2340 3911 2347 3963
rect 2399 3911 2406 3963
rect 2340 3899 2406 3911
rect 2340 3847 2347 3899
rect 2399 3847 2406 3899
rect 2340 3835 2406 3847
rect 2340 3783 2347 3835
rect 2399 3783 2406 3835
rect 2340 3771 2406 3783
rect 2340 3719 2347 3771
rect 2399 3719 2406 3771
rect 2340 3707 2406 3719
rect 2340 3655 2347 3707
rect 2399 3655 2406 3707
rect 2340 3643 2406 3655
rect 2340 3591 2347 3643
rect 2399 3591 2406 3643
rect 2340 3579 2406 3591
rect 2340 3527 2347 3579
rect 2399 3527 2406 3579
rect 2340 3515 2406 3527
rect 2340 3463 2347 3515
rect 2399 3463 2406 3515
rect 2340 3451 2406 3463
rect 2340 3399 2347 3451
rect 2399 3399 2406 3451
rect 2340 3387 2406 3399
rect 2340 3335 2347 3387
rect 2399 3335 2406 3387
rect 2340 3323 2406 3335
rect 2340 3271 2347 3323
rect 2399 3271 2406 3323
rect 2340 3259 2406 3271
rect 2340 3207 2347 3259
rect 2399 3207 2406 3259
rect 2340 3195 2406 3207
rect 2340 3143 2347 3195
rect 2399 3143 2406 3195
rect 2340 3131 2406 3143
rect 2340 3079 2347 3131
rect 2399 3079 2406 3131
rect 2340 3067 2406 3079
rect 2340 3015 2347 3067
rect 2399 3015 2406 3067
rect 2340 3003 2406 3015
rect 2340 2951 2347 3003
rect 2399 2951 2406 3003
rect 2340 2939 2406 2951
rect 2340 2887 2347 2939
rect 2399 2887 2406 2939
rect 2340 2875 2406 2887
rect 2340 2823 2347 2875
rect 2399 2823 2406 2875
rect 2340 2811 2406 2823
rect 2340 2759 2347 2811
rect 2399 2759 2406 2811
rect 2340 2746 2406 2759
rect 3256 4347 3322 4360
rect 3724 4352 3770 4502
rect 3256 4295 3263 4347
rect 3315 4295 3322 4347
rect 3256 4283 3322 4295
rect 3256 4231 3263 4283
rect 3315 4231 3322 4283
rect 3256 4219 3322 4231
rect 3256 4167 3263 4219
rect 3315 4167 3322 4219
rect 3256 4155 3322 4167
rect 3256 4103 3263 4155
rect 3315 4103 3322 4155
rect 3256 4091 3322 4103
rect 3256 4039 3263 4091
rect 3315 4039 3322 4091
rect 3256 4027 3322 4039
rect 3256 3975 3263 4027
rect 3315 3975 3322 4027
rect 3256 3963 3322 3975
rect 3256 3911 3263 3963
rect 3315 3911 3322 3963
rect 3256 3899 3322 3911
rect 3256 3847 3263 3899
rect 3315 3847 3322 3899
rect 3256 3835 3322 3847
rect 3256 3783 3263 3835
rect 3315 3783 3322 3835
rect 3256 3771 3322 3783
rect 3256 3719 3263 3771
rect 3315 3719 3322 3771
rect 3256 3707 3322 3719
rect 3256 3655 3263 3707
rect 3315 3655 3322 3707
rect 3256 3643 3322 3655
rect 3256 3591 3263 3643
rect 3315 3591 3322 3643
rect 3256 3579 3322 3591
rect 3256 3527 3263 3579
rect 3315 3527 3322 3579
rect 3256 3515 3322 3527
rect 3256 3463 3263 3515
rect 3315 3463 3322 3515
rect 3256 3451 3322 3463
rect 3256 3399 3263 3451
rect 3315 3399 3322 3451
rect 3256 3387 3322 3399
rect 3256 3335 3263 3387
rect 3315 3335 3322 3387
rect 3256 3323 3322 3335
rect 3256 3271 3263 3323
rect 3315 3271 3322 3323
rect 3256 3259 3322 3271
rect 3256 3207 3263 3259
rect 3315 3207 3322 3259
rect 3256 3195 3322 3207
rect 3256 3143 3263 3195
rect 3315 3143 3322 3195
rect 3256 3131 3322 3143
rect 3256 3079 3263 3131
rect 3315 3079 3322 3131
rect 3256 3067 3322 3079
rect 3256 3015 3263 3067
rect 3315 3015 3322 3067
rect 3256 3003 3322 3015
rect 3256 2951 3263 3003
rect 3315 2951 3322 3003
rect 3256 2939 3322 2951
rect 3256 2887 3263 2939
rect 3315 2887 3322 2939
rect 3256 2875 3322 2887
rect 3256 2823 3263 2875
rect 3315 2823 3322 2875
rect 3256 2811 3322 2823
rect 3256 2759 3263 2811
rect 3315 2759 3322 2811
rect 3256 2746 3322 2759
rect 836 2660 851 2712
rect 903 2660 918 2712
rect 1208 2706 1374 2744
rect 1208 2672 1220 2706
rect 1254 2672 1326 2706
rect 1360 2672 1374 2706
rect 1208 2652 1374 2672
rect 1638 2660 1653 2712
rect 1705 2660 1720 2712
rect 178 2407 672 2418
rect 178 2064 207 2407
rect 106 2035 207 2064
rect 643 2064 672 2407
rect 1604 2413 2098 2424
rect 818 2083 898 2096
rect 818 2064 833 2083
rect 643 2035 833 2064
rect 106 2031 833 2035
rect 885 2064 898 2083
rect 1604 2064 1633 2413
rect 885 2031 1256 2064
rect 106 1966 1256 2031
rect 1378 2041 1633 2064
rect 2069 2064 2098 2413
rect 2069 2041 2214 2064
rect 1378 2031 2214 2041
rect 1378 1979 1401 2031
rect 1453 1979 2214 2031
rect 1378 1966 2214 1979
rect 10 1665 56 1698
rect 10 1631 16 1665
rect 50 1631 56 1665
rect 10 1330 56 1631
rect 106 1665 152 1966
rect 106 1631 112 1665
rect 146 1631 152 1665
rect 106 1598 152 1631
rect 202 1665 248 1698
rect 202 1631 208 1665
rect 242 1631 248 1665
rect 90 1560 174 1568
rect 90 1559 116 1560
rect 150 1559 174 1560
rect 90 1507 106 1559
rect 158 1507 174 1559
rect 90 1498 174 1507
rect 202 1330 248 1631
rect 298 1665 344 1966
rect 298 1631 304 1665
rect 338 1631 344 1665
rect 298 1598 344 1631
rect 394 1665 440 1698
rect 394 1631 400 1665
rect 434 1631 440 1665
rect 394 1330 440 1631
rect 490 1665 536 1966
rect 490 1631 496 1665
rect 530 1631 536 1665
rect 490 1598 536 1631
rect 586 1665 632 1698
rect 586 1631 592 1665
rect 626 1631 632 1665
rect 586 1330 632 1631
rect 682 1665 728 1966
rect 682 1631 688 1665
rect 722 1631 728 1665
rect 682 1598 728 1631
rect 778 1665 824 1698
rect 778 1631 784 1665
rect 818 1631 824 1665
rect 778 1330 824 1631
rect 874 1665 920 1966
rect 874 1631 880 1665
rect 914 1631 920 1665
rect 874 1598 920 1631
rect 970 1665 1016 1698
rect 970 1631 976 1665
rect 1010 1631 1016 1665
rect 970 1330 1016 1631
rect 1304 1665 1350 1698
rect 1304 1631 1310 1665
rect 1344 1631 1350 1665
rect 1304 1330 1350 1631
rect 1400 1665 1446 1966
rect 1400 1631 1406 1665
rect 1440 1631 1446 1665
rect 1400 1598 1446 1631
rect 1496 1665 1542 1698
rect 1496 1631 1502 1665
rect 1536 1631 1542 1665
rect 1496 1330 1542 1631
rect 1592 1665 1638 1966
rect 1592 1631 1598 1665
rect 1632 1631 1638 1665
rect 1592 1598 1638 1631
rect 1688 1665 1734 1698
rect 1688 1631 1694 1665
rect 1728 1631 1734 1665
rect 1688 1330 1734 1631
rect 1784 1665 1830 1966
rect 1784 1631 1790 1665
rect 1824 1631 1830 1665
rect 1784 1598 1830 1631
rect 1880 1665 1926 1698
rect 1880 1631 1886 1665
rect 1920 1631 1926 1665
rect 1880 1330 1926 1631
rect 1976 1665 2022 1966
rect 1976 1631 1982 1665
rect 2016 1631 2022 1665
rect 1976 1598 2022 1631
rect 2072 1665 2118 1698
rect 2072 1631 2078 1665
rect 2112 1631 2118 1665
rect 2072 1330 2118 1631
rect 2168 1665 2214 1966
rect 2290 1770 2534 1790
rect 2290 1736 2302 1770
rect 2336 1736 2534 1770
rect 2290 1728 2534 1736
rect 2168 1631 2174 1665
rect 2208 1631 2214 1665
rect 2168 1598 2214 1631
rect 2264 1665 2310 1698
rect 2264 1631 2270 1665
rect 2304 1631 2310 1665
rect 2264 1330 2310 1631
rect 10 1243 2310 1330
rect 10 1191 713 1243
rect 765 1233 2310 1243
rect 765 1191 1555 1233
rect 10 1181 1555 1191
rect 1607 1232 2310 1233
rect 1607 1181 2306 1232
rect 10 1103 2306 1181
rect 10 1099 1553 1103
rect 10 1047 717 1099
rect 769 1051 1553 1099
rect 1605 1051 2306 1103
rect 769 1047 2306 1051
rect 10 1032 2306 1047
rect 6 934 2306 1032
rect 6 566 52 934
rect 86 757 170 766
rect 86 705 102 757
rect 154 705 170 757
rect 86 704 114 705
rect 148 704 170 705
rect 86 696 170 704
rect 102 324 148 666
rect 198 566 244 934
rect 294 324 340 666
rect 390 566 436 934
rect 486 324 532 666
rect 582 566 628 934
rect 678 324 724 666
rect 774 566 820 934
rect 870 324 916 666
rect 966 566 1012 934
rect 1300 633 1346 934
rect 1300 599 1306 633
rect 1340 599 1346 633
rect 1300 566 1346 599
rect 1396 633 1442 666
rect 1396 599 1402 633
rect 1436 599 1442 633
rect 1396 324 1442 599
rect 1492 633 1538 934
rect 1492 599 1498 633
rect 1532 599 1538 633
rect 1492 566 1538 599
rect 1588 633 1634 666
rect 1588 599 1594 633
rect 1628 599 1634 633
rect 1588 324 1634 599
rect 1684 633 1730 934
rect 1684 599 1690 633
rect 1724 599 1730 633
rect 1684 566 1730 599
rect 1780 633 1826 666
rect 1780 599 1786 633
rect 1820 599 1826 633
rect 1780 324 1826 599
rect 1876 633 1922 934
rect 1876 599 1882 633
rect 1916 599 1922 633
rect 1876 566 1922 599
rect 1972 633 2018 666
rect 1972 599 1978 633
rect 2012 599 2018 633
rect 1972 324 2018 599
rect 2068 633 2114 934
rect 2068 599 2074 633
rect 2108 599 2114 633
rect 2068 566 2114 599
rect 2164 633 2210 666
rect 2164 599 2170 633
rect 2204 599 2210 633
rect 2164 324 2210 599
rect 2260 633 2306 934
rect 2458 882 2534 1728
rect 2458 830 2470 882
rect 2522 830 2534 882
rect 2458 826 2534 830
rect 2606 1434 2682 1438
rect 2606 1382 2618 1434
rect 2670 1382 2682 1434
rect 2260 599 2266 633
rect 2300 599 2306 633
rect 2260 566 2306 599
rect 2606 536 2682 1382
rect 2284 528 2682 536
rect 2284 494 2296 528
rect 2330 494 2682 528
rect 2284 474 2682 494
rect 102 297 1120 324
rect 102 245 1045 297
rect 1097 245 1120 297
rect 102 226 1120 245
rect 1192 299 2210 324
rect 1192 247 1213 299
rect 1265 247 2210 299
rect 1192 226 2210 247
rect -1160 -563 -1092 -542
rect -1160 -615 -1152 -563
rect -1100 -615 -1092 -563
rect -1160 -627 -1092 -615
rect -1160 -679 -1152 -627
rect -1100 -679 -1092 -627
rect -1160 -691 -1092 -679
rect -1160 -743 -1152 -691
rect -1100 -743 -1092 -691
rect -1160 -755 -1092 -743
rect -1160 -807 -1152 -755
rect -1100 -807 -1092 -755
rect -1160 -819 -1092 -807
rect -1160 -871 -1152 -819
rect -1100 -871 -1092 -819
rect -1160 -883 -1092 -871
rect -1160 -935 -1152 -883
rect -1100 -935 -1092 -883
rect -1160 -947 -1092 -935
rect -1160 -999 -1152 -947
rect -1100 -999 -1092 -947
rect -1160 -1011 -1092 -999
rect -1160 -1063 -1152 -1011
rect -1100 -1063 -1092 -1011
rect -1160 -1075 -1092 -1063
rect -1160 -1127 -1152 -1075
rect -1100 -1127 -1092 -1075
rect -1160 -1139 -1092 -1127
rect -1160 -1191 -1152 -1139
rect -1100 -1191 -1092 -1139
rect -1160 -1203 -1092 -1191
rect -1160 -1255 -1152 -1203
rect -1100 -1255 -1092 -1203
rect -1160 -1267 -1092 -1255
rect -1160 -1319 -1152 -1267
rect -1100 -1319 -1092 -1267
rect -1160 -1331 -1092 -1319
rect -1160 -1383 -1152 -1331
rect -1100 -1383 -1092 -1331
rect -1160 -1395 -1092 -1383
rect -1160 -1447 -1152 -1395
rect -1100 -1447 -1092 -1395
rect -1160 -1459 -1092 -1447
rect -1160 -1511 -1152 -1459
rect -1100 -1511 -1092 -1459
rect -1160 -1523 -1092 -1511
rect -1160 -1575 -1152 -1523
rect -1100 -1575 -1092 -1523
rect -1160 -1587 -1092 -1575
rect -1160 -1639 -1152 -1587
rect -1100 -1639 -1092 -1587
rect -1160 -1651 -1092 -1639
rect -1160 -1703 -1152 -1651
rect -1100 -1703 -1092 -1651
rect -1160 -1715 -1092 -1703
rect -1160 -1767 -1152 -1715
rect -1100 -1767 -1092 -1715
rect -1160 -1779 -1092 -1767
rect -1160 -1831 -1152 -1779
rect -1100 -1831 -1092 -1779
rect -1160 -1843 -1092 -1831
rect -1160 -1895 -1152 -1843
rect -1100 -1895 -1092 -1843
rect -1160 -1907 -1092 -1895
rect -1160 -1959 -1152 -1907
rect -1100 -1959 -1092 -1907
rect -1160 -1971 -1092 -1959
rect -1160 -2023 -1152 -1971
rect -1100 -2023 -1092 -1971
rect -1160 -2035 -1092 -2023
rect -1160 -2087 -1152 -2035
rect -1100 -2087 -1092 -2035
rect -1160 -2099 -1092 -2087
rect -1160 -2151 -1152 -2099
rect -1100 -2151 -1092 -2099
rect -1160 -2163 -1092 -2151
rect -1160 -2215 -1152 -2163
rect -1100 -2215 -1092 -2163
rect -1160 -2227 -1092 -2215
rect -1160 -2279 -1152 -2227
rect -1100 -2279 -1092 -2227
rect -1160 -2291 -1092 -2279
rect -1160 -2343 -1152 -2291
rect -1100 -2343 -1092 -2291
rect -1160 -2355 -1092 -2343
rect -1160 -2407 -1152 -2355
rect -1100 -2407 -1092 -2355
rect -1160 -2419 -1092 -2407
rect -1160 -2471 -1152 -2419
rect -1100 -2471 -1092 -2419
rect -1160 -2483 -1092 -2471
rect -1160 -2535 -1152 -2483
rect -1100 -2535 -1092 -2483
rect -1160 -2547 -1092 -2535
rect -1160 -2599 -1152 -2547
rect -1100 -2599 -1092 -2547
rect -1160 -2611 -1092 -2599
rect -1160 -2663 -1152 -2611
rect -1100 -2663 -1092 -2611
rect -1160 -2675 -1092 -2663
rect -1160 -2727 -1152 -2675
rect -1100 -2727 -1092 -2675
rect -1160 -2739 -1092 -2727
rect -1160 -2791 -1152 -2739
rect -1100 -2791 -1092 -2739
rect -1160 -2803 -1092 -2791
rect -1160 -2855 -1152 -2803
rect -1100 -2855 -1092 -2803
rect -1160 -2867 -1092 -2855
rect -1160 -2919 -1152 -2867
rect -1100 -2919 -1092 -2867
rect -1160 -2931 -1092 -2919
rect -1160 -2983 -1152 -2931
rect -1100 -2983 -1092 -2931
rect -1160 -2995 -1092 -2983
rect -1160 -3047 -1152 -2995
rect -1100 -3047 -1092 -2995
rect -1160 -3059 -1092 -3047
rect -1160 -3111 -1152 -3059
rect -1100 -3111 -1092 -3059
rect -1160 -3123 -1092 -3111
rect -1160 -3175 -1152 -3123
rect -1100 -3175 -1092 -3123
rect -1160 -3196 -1092 -3175
rect -702 -563 -634 -542
rect -702 -615 -694 -563
rect -642 -615 -634 -563
rect -702 -627 -634 -615
rect -702 -679 -694 -627
rect -642 -679 -634 -627
rect -702 -691 -634 -679
rect -702 -743 -694 -691
rect -642 -743 -634 -691
rect -702 -755 -634 -743
rect -702 -807 -694 -755
rect -642 -807 -634 -755
rect -702 -819 -634 -807
rect -702 -871 -694 -819
rect -642 -871 -634 -819
rect -702 -883 -634 -871
rect -702 -935 -694 -883
rect -642 -935 -634 -883
rect -702 -947 -634 -935
rect -702 -999 -694 -947
rect -642 -999 -634 -947
rect -702 -1011 -634 -999
rect -702 -1063 -694 -1011
rect -642 -1063 -634 -1011
rect -702 -1075 -634 -1063
rect -702 -1127 -694 -1075
rect -642 -1127 -634 -1075
rect -702 -1139 -634 -1127
rect -702 -1191 -694 -1139
rect -642 -1191 -634 -1139
rect -702 -1203 -634 -1191
rect -702 -1255 -694 -1203
rect -642 -1255 -634 -1203
rect -702 -1267 -634 -1255
rect -702 -1319 -694 -1267
rect -642 -1319 -634 -1267
rect -702 -1331 -634 -1319
rect -702 -1383 -694 -1331
rect -642 -1383 -634 -1331
rect -702 -1395 -634 -1383
rect -702 -1447 -694 -1395
rect -642 -1447 -634 -1395
rect -702 -1459 -634 -1447
rect -702 -1511 -694 -1459
rect -642 -1511 -634 -1459
rect -702 -1523 -634 -1511
rect -702 -1575 -694 -1523
rect -642 -1575 -634 -1523
rect -702 -1587 -634 -1575
rect -702 -1639 -694 -1587
rect -642 -1639 -634 -1587
rect -702 -1651 -634 -1639
rect -702 -1703 -694 -1651
rect -642 -1703 -634 -1651
rect -702 -1715 -634 -1703
rect -702 -1767 -694 -1715
rect -642 -1767 -634 -1715
rect -702 -1779 -634 -1767
rect -702 -1831 -694 -1779
rect -642 -1831 -634 -1779
rect -702 -1843 -634 -1831
rect -702 -1895 -694 -1843
rect -642 -1895 -634 -1843
rect -702 -1907 -634 -1895
rect -702 -1959 -694 -1907
rect -642 -1959 -634 -1907
rect -702 -1971 -634 -1959
rect -702 -2023 -694 -1971
rect -642 -2023 -634 -1971
rect -702 -2035 -634 -2023
rect -702 -2087 -694 -2035
rect -642 -2087 -634 -2035
rect -702 -2099 -634 -2087
rect -702 -2151 -694 -2099
rect -642 -2151 -634 -2099
rect -702 -2163 -634 -2151
rect -702 -2215 -694 -2163
rect -642 -2215 -634 -2163
rect -702 -2227 -634 -2215
rect -702 -2279 -694 -2227
rect -642 -2279 -634 -2227
rect -702 -2291 -634 -2279
rect -702 -2343 -694 -2291
rect -642 -2343 -634 -2291
rect -702 -2355 -634 -2343
rect -702 -2407 -694 -2355
rect -642 -2407 -634 -2355
rect -702 -2419 -634 -2407
rect -702 -2471 -694 -2419
rect -642 -2471 -634 -2419
rect -702 -2483 -634 -2471
rect -702 -2535 -694 -2483
rect -642 -2535 -634 -2483
rect -702 -2547 -634 -2535
rect -702 -2599 -694 -2547
rect -642 -2599 -634 -2547
rect -702 -2611 -634 -2599
rect -702 -2663 -694 -2611
rect -642 -2663 -634 -2611
rect -702 -2675 -634 -2663
rect -702 -2727 -694 -2675
rect -642 -2727 -634 -2675
rect -702 -2739 -634 -2727
rect -702 -2791 -694 -2739
rect -642 -2791 -634 -2739
rect -702 -2803 -634 -2791
rect -702 -2855 -694 -2803
rect -642 -2855 -634 -2803
rect -702 -2867 -634 -2855
rect -702 -2919 -694 -2867
rect -642 -2919 -634 -2867
rect -702 -2931 -634 -2919
rect -702 -2983 -694 -2931
rect -642 -2983 -634 -2931
rect -702 -2995 -634 -2983
rect -702 -3047 -694 -2995
rect -642 -3047 -634 -2995
rect -702 -3059 -634 -3047
rect -702 -3111 -694 -3059
rect -642 -3111 -634 -3059
rect -702 -3123 -634 -3111
rect -702 -3175 -694 -3123
rect -642 -3175 -634 -3123
rect -702 -3196 -634 -3175
rect -244 -563 -176 -542
rect -244 -615 -236 -563
rect -184 -615 -176 -563
rect -244 -627 -176 -615
rect -244 -679 -236 -627
rect -184 -679 -176 -627
rect -244 -691 -176 -679
rect -244 -743 -236 -691
rect -184 -743 -176 -691
rect -244 -755 -176 -743
rect -244 -807 -236 -755
rect -184 -807 -176 -755
rect -244 -819 -176 -807
rect -244 -871 -236 -819
rect -184 -871 -176 -819
rect -244 -883 -176 -871
rect -244 -935 -236 -883
rect -184 -935 -176 -883
rect -244 -947 -176 -935
rect -244 -999 -236 -947
rect -184 -999 -176 -947
rect -244 -1011 -176 -999
rect -244 -1063 -236 -1011
rect -184 -1063 -176 -1011
rect -244 -1075 -176 -1063
rect -244 -1127 -236 -1075
rect -184 -1127 -176 -1075
rect -244 -1139 -176 -1127
rect -244 -1191 -236 -1139
rect -184 -1191 -176 -1139
rect -244 -1203 -176 -1191
rect -244 -1255 -236 -1203
rect -184 -1255 -176 -1203
rect -244 -1267 -176 -1255
rect -244 -1319 -236 -1267
rect -184 -1319 -176 -1267
rect -244 -1331 -176 -1319
rect -244 -1383 -236 -1331
rect -184 -1383 -176 -1331
rect -244 -1395 -176 -1383
rect -244 -1447 -236 -1395
rect -184 -1447 -176 -1395
rect -244 -1459 -176 -1447
rect -244 -1511 -236 -1459
rect -184 -1511 -176 -1459
rect -244 -1523 -176 -1511
rect -244 -1575 -236 -1523
rect -184 -1575 -176 -1523
rect -244 -1587 -176 -1575
rect -244 -1639 -236 -1587
rect -184 -1639 -176 -1587
rect -244 -1651 -176 -1639
rect -244 -1703 -236 -1651
rect -184 -1703 -176 -1651
rect -244 -1715 -176 -1703
rect -244 -1767 -236 -1715
rect -184 -1767 -176 -1715
rect -244 -1779 -176 -1767
rect -244 -1831 -236 -1779
rect -184 -1831 -176 -1779
rect -244 -1843 -176 -1831
rect -244 -1895 -236 -1843
rect -184 -1895 -176 -1843
rect -244 -1907 -176 -1895
rect -244 -1959 -236 -1907
rect -184 -1959 -176 -1907
rect -244 -1971 -176 -1959
rect -244 -2023 -236 -1971
rect -184 -2023 -176 -1971
rect -244 -2035 -176 -2023
rect -244 -2087 -236 -2035
rect -184 -2087 -176 -2035
rect -244 -2099 -176 -2087
rect -244 -2151 -236 -2099
rect -184 -2151 -176 -2099
rect -244 -2163 -176 -2151
rect -244 -2215 -236 -2163
rect -184 -2215 -176 -2163
rect -244 -2227 -176 -2215
rect -244 -2279 -236 -2227
rect -184 -2279 -176 -2227
rect -244 -2291 -176 -2279
rect -244 -2343 -236 -2291
rect -184 -2343 -176 -2291
rect -244 -2355 -176 -2343
rect -244 -2407 -236 -2355
rect -184 -2407 -176 -2355
rect -244 -2419 -176 -2407
rect -244 -2471 -236 -2419
rect -184 -2471 -176 -2419
rect -244 -2483 -176 -2471
rect -244 -2535 -236 -2483
rect -184 -2535 -176 -2483
rect -244 -2547 -176 -2535
rect -244 -2599 -236 -2547
rect -184 -2599 -176 -2547
rect -244 -2611 -176 -2599
rect -244 -2663 -236 -2611
rect -184 -2663 -176 -2611
rect -244 -2675 -176 -2663
rect -244 -2727 -236 -2675
rect -184 -2727 -176 -2675
rect -244 -2739 -176 -2727
rect -244 -2791 -236 -2739
rect -184 -2791 -176 -2739
rect -244 -2803 -176 -2791
rect -244 -2855 -236 -2803
rect -184 -2855 -176 -2803
rect -244 -2867 -176 -2855
rect -244 -2919 -236 -2867
rect -184 -2919 -176 -2867
rect -244 -2931 -176 -2919
rect -244 -2983 -236 -2931
rect -184 -2983 -176 -2931
rect -244 -2995 -176 -2983
rect -244 -3047 -236 -2995
rect -184 -3047 -176 -2995
rect -244 -3059 -176 -3047
rect -244 -3111 -236 -3059
rect -184 -3111 -176 -3059
rect -244 -3123 -176 -3111
rect -244 -3175 -236 -3123
rect -184 -3175 -176 -3123
rect -244 -3196 -176 -3175
rect 214 -563 282 -542
rect 214 -615 222 -563
rect 274 -615 282 -563
rect 214 -627 282 -615
rect 214 -679 222 -627
rect 274 -679 282 -627
rect 214 -691 282 -679
rect 214 -743 222 -691
rect 274 -743 282 -691
rect 214 -755 282 -743
rect 214 -807 222 -755
rect 274 -807 282 -755
rect 214 -819 282 -807
rect 214 -871 222 -819
rect 274 -871 282 -819
rect 214 -883 282 -871
rect 214 -935 222 -883
rect 274 -935 282 -883
rect 214 -947 282 -935
rect 214 -999 222 -947
rect 274 -999 282 -947
rect 214 -1011 282 -999
rect 214 -1063 222 -1011
rect 274 -1063 282 -1011
rect 214 -1075 282 -1063
rect 214 -1127 222 -1075
rect 274 -1127 282 -1075
rect 214 -1139 282 -1127
rect 214 -1191 222 -1139
rect 274 -1191 282 -1139
rect 214 -1203 282 -1191
rect 214 -1255 222 -1203
rect 274 -1255 282 -1203
rect 214 -1267 282 -1255
rect 214 -1319 222 -1267
rect 274 -1319 282 -1267
rect 214 -1331 282 -1319
rect 214 -1383 222 -1331
rect 274 -1383 282 -1331
rect 214 -1395 282 -1383
rect 214 -1447 222 -1395
rect 274 -1447 282 -1395
rect 214 -1459 282 -1447
rect 214 -1511 222 -1459
rect 274 -1511 282 -1459
rect 214 -1523 282 -1511
rect 214 -1575 222 -1523
rect 274 -1575 282 -1523
rect 214 -1587 282 -1575
rect 214 -1639 222 -1587
rect 274 -1639 282 -1587
rect 214 -1651 282 -1639
rect 214 -1703 222 -1651
rect 274 -1703 282 -1651
rect 214 -1715 282 -1703
rect 214 -1767 222 -1715
rect 274 -1767 282 -1715
rect 214 -1779 282 -1767
rect 214 -1831 222 -1779
rect 274 -1831 282 -1779
rect 214 -1843 282 -1831
rect 214 -1895 222 -1843
rect 274 -1895 282 -1843
rect 214 -1907 282 -1895
rect 214 -1959 222 -1907
rect 274 -1959 282 -1907
rect 214 -1971 282 -1959
rect 214 -2023 222 -1971
rect 274 -2023 282 -1971
rect 214 -2035 282 -2023
rect 214 -2087 222 -2035
rect 274 -2087 282 -2035
rect 214 -2099 282 -2087
rect 214 -2151 222 -2099
rect 274 -2151 282 -2099
rect 214 -2163 282 -2151
rect 214 -2215 222 -2163
rect 274 -2215 282 -2163
rect 214 -2227 282 -2215
rect 214 -2279 222 -2227
rect 274 -2279 282 -2227
rect 214 -2291 282 -2279
rect 214 -2343 222 -2291
rect 274 -2343 282 -2291
rect 214 -2355 282 -2343
rect 214 -2407 222 -2355
rect 274 -2407 282 -2355
rect 214 -2419 282 -2407
rect 214 -2471 222 -2419
rect 274 -2471 282 -2419
rect 214 -2483 282 -2471
rect 214 -2535 222 -2483
rect 274 -2535 282 -2483
rect 214 -2547 282 -2535
rect 214 -2599 222 -2547
rect 274 -2599 282 -2547
rect 214 -2611 282 -2599
rect 214 -2663 222 -2611
rect 274 -2663 282 -2611
rect 214 -2675 282 -2663
rect 214 -2727 222 -2675
rect 274 -2727 282 -2675
rect 214 -2739 282 -2727
rect 214 -2791 222 -2739
rect 274 -2791 282 -2739
rect 214 -2803 282 -2791
rect 214 -2855 222 -2803
rect 274 -2855 282 -2803
rect 214 -2867 282 -2855
rect 214 -2919 222 -2867
rect 274 -2919 282 -2867
rect 214 -2931 282 -2919
rect 214 -2983 222 -2931
rect 274 -2983 282 -2931
rect 214 -2995 282 -2983
rect 214 -3047 222 -2995
rect 274 -3047 282 -2995
rect 214 -3059 282 -3047
rect 214 -3111 222 -3059
rect 274 -3111 282 -3059
rect 214 -3123 282 -3111
rect 214 -3175 222 -3123
rect 274 -3175 282 -3123
rect 214 -3196 282 -3175
rect 672 -563 740 -542
rect 672 -615 680 -563
rect 732 -615 740 -563
rect 672 -627 740 -615
rect 672 -679 680 -627
rect 732 -679 740 -627
rect 672 -691 740 -679
rect 672 -743 680 -691
rect 732 -743 740 -691
rect 672 -755 740 -743
rect 672 -807 680 -755
rect 732 -807 740 -755
rect 672 -819 740 -807
rect 672 -871 680 -819
rect 732 -871 740 -819
rect 672 -883 740 -871
rect 672 -935 680 -883
rect 732 -935 740 -883
rect 672 -947 740 -935
rect 672 -999 680 -947
rect 732 -999 740 -947
rect 672 -1011 740 -999
rect 672 -1063 680 -1011
rect 732 -1063 740 -1011
rect 672 -1075 740 -1063
rect 672 -1127 680 -1075
rect 732 -1127 740 -1075
rect 672 -1139 740 -1127
rect 672 -1191 680 -1139
rect 732 -1191 740 -1139
rect 672 -1203 740 -1191
rect 672 -1255 680 -1203
rect 732 -1255 740 -1203
rect 672 -1267 740 -1255
rect 672 -1319 680 -1267
rect 732 -1319 740 -1267
rect 672 -1331 740 -1319
rect 672 -1383 680 -1331
rect 732 -1383 740 -1331
rect 672 -1395 740 -1383
rect 672 -1447 680 -1395
rect 732 -1447 740 -1395
rect 672 -1459 740 -1447
rect 672 -1511 680 -1459
rect 732 -1511 740 -1459
rect 672 -1523 740 -1511
rect 672 -1575 680 -1523
rect 732 -1575 740 -1523
rect 672 -1587 740 -1575
rect 672 -1639 680 -1587
rect 732 -1639 740 -1587
rect 672 -1651 740 -1639
rect 672 -1703 680 -1651
rect 732 -1703 740 -1651
rect 672 -1715 740 -1703
rect 672 -1767 680 -1715
rect 732 -1767 740 -1715
rect 672 -1779 740 -1767
rect 672 -1831 680 -1779
rect 732 -1831 740 -1779
rect 672 -1843 740 -1831
rect 672 -1895 680 -1843
rect 732 -1895 740 -1843
rect 672 -1907 740 -1895
rect 672 -1959 680 -1907
rect 732 -1959 740 -1907
rect 672 -1971 740 -1959
rect 672 -2023 680 -1971
rect 732 -2023 740 -1971
rect 672 -2035 740 -2023
rect 672 -2087 680 -2035
rect 732 -2087 740 -2035
rect 672 -2099 740 -2087
rect 672 -2151 680 -2099
rect 732 -2151 740 -2099
rect 672 -2163 740 -2151
rect 672 -2215 680 -2163
rect 732 -2215 740 -2163
rect 672 -2227 740 -2215
rect 672 -2279 680 -2227
rect 732 -2279 740 -2227
rect 672 -2291 740 -2279
rect 672 -2343 680 -2291
rect 732 -2343 740 -2291
rect 672 -2355 740 -2343
rect 672 -2407 680 -2355
rect 732 -2407 740 -2355
rect 672 -2419 740 -2407
rect 672 -2471 680 -2419
rect 732 -2471 740 -2419
rect 672 -2483 740 -2471
rect 672 -2535 680 -2483
rect 732 -2535 740 -2483
rect 672 -2547 740 -2535
rect 672 -2599 680 -2547
rect 732 -2599 740 -2547
rect 672 -2611 740 -2599
rect 672 -2663 680 -2611
rect 732 -2663 740 -2611
rect 672 -2675 740 -2663
rect 672 -2727 680 -2675
rect 732 -2727 740 -2675
rect 672 -2739 740 -2727
rect 672 -2791 680 -2739
rect 732 -2791 740 -2739
rect 672 -2803 740 -2791
rect 672 -2855 680 -2803
rect 732 -2855 740 -2803
rect 672 -2867 740 -2855
rect 672 -2919 680 -2867
rect 732 -2919 740 -2867
rect 672 -2931 740 -2919
rect 672 -2983 680 -2931
rect 732 -2983 740 -2931
rect 672 -2995 740 -2983
rect 672 -3047 680 -2995
rect 732 -3047 740 -2995
rect 672 -3059 740 -3047
rect 672 -3111 680 -3059
rect 732 -3111 740 -3059
rect 672 -3123 740 -3111
rect 672 -3175 680 -3123
rect 732 -3175 740 -3123
rect 672 -3196 740 -3175
rect 1130 -563 1198 -542
rect 1130 -615 1138 -563
rect 1190 -615 1198 -563
rect 1130 -627 1198 -615
rect 1130 -679 1138 -627
rect 1190 -679 1198 -627
rect 1130 -691 1198 -679
rect 1130 -743 1138 -691
rect 1190 -743 1198 -691
rect 1130 -755 1198 -743
rect 1130 -807 1138 -755
rect 1190 -807 1198 -755
rect 1130 -819 1198 -807
rect 1130 -871 1138 -819
rect 1190 -871 1198 -819
rect 1130 -883 1198 -871
rect 1130 -935 1138 -883
rect 1190 -935 1198 -883
rect 1130 -947 1198 -935
rect 1130 -999 1138 -947
rect 1190 -999 1198 -947
rect 1130 -1011 1198 -999
rect 1130 -1063 1138 -1011
rect 1190 -1063 1198 -1011
rect 1130 -1075 1198 -1063
rect 1130 -1127 1138 -1075
rect 1190 -1127 1198 -1075
rect 1130 -1139 1198 -1127
rect 1130 -1191 1138 -1139
rect 1190 -1191 1198 -1139
rect 1130 -1203 1198 -1191
rect 1130 -1255 1138 -1203
rect 1190 -1255 1198 -1203
rect 1130 -1267 1198 -1255
rect 1130 -1319 1138 -1267
rect 1190 -1319 1198 -1267
rect 1130 -1331 1198 -1319
rect 1130 -1383 1138 -1331
rect 1190 -1383 1198 -1331
rect 1130 -1395 1198 -1383
rect 1130 -1447 1138 -1395
rect 1190 -1447 1198 -1395
rect 1130 -1459 1198 -1447
rect 1130 -1511 1138 -1459
rect 1190 -1511 1198 -1459
rect 1130 -1523 1198 -1511
rect 1130 -1575 1138 -1523
rect 1190 -1575 1198 -1523
rect 1130 -1587 1198 -1575
rect 1130 -1639 1138 -1587
rect 1190 -1639 1198 -1587
rect 1130 -1651 1198 -1639
rect 1130 -1703 1138 -1651
rect 1190 -1703 1198 -1651
rect 1130 -1715 1198 -1703
rect 1130 -1767 1138 -1715
rect 1190 -1767 1198 -1715
rect 1130 -1779 1198 -1767
rect 1130 -1831 1138 -1779
rect 1190 -1831 1198 -1779
rect 1130 -1843 1198 -1831
rect 1130 -1895 1138 -1843
rect 1190 -1895 1198 -1843
rect 1130 -1907 1198 -1895
rect 1130 -1959 1138 -1907
rect 1190 -1959 1198 -1907
rect 1130 -1971 1198 -1959
rect 1130 -2023 1138 -1971
rect 1190 -2023 1198 -1971
rect 1130 -2035 1198 -2023
rect 1130 -2087 1138 -2035
rect 1190 -2087 1198 -2035
rect 1130 -2099 1198 -2087
rect 1130 -2151 1138 -2099
rect 1190 -2151 1198 -2099
rect 1130 -2163 1198 -2151
rect 1130 -2215 1138 -2163
rect 1190 -2215 1198 -2163
rect 1130 -2227 1198 -2215
rect 1130 -2279 1138 -2227
rect 1190 -2279 1198 -2227
rect 1130 -2291 1198 -2279
rect 1130 -2343 1138 -2291
rect 1190 -2343 1198 -2291
rect 1130 -2355 1198 -2343
rect 1130 -2407 1138 -2355
rect 1190 -2407 1198 -2355
rect 1130 -2419 1198 -2407
rect 1130 -2471 1138 -2419
rect 1190 -2471 1198 -2419
rect 1130 -2483 1198 -2471
rect 1130 -2535 1138 -2483
rect 1190 -2535 1198 -2483
rect 1130 -2547 1198 -2535
rect 1130 -2599 1138 -2547
rect 1190 -2599 1198 -2547
rect 1130 -2611 1198 -2599
rect 1130 -2663 1138 -2611
rect 1190 -2663 1198 -2611
rect 1130 -2675 1198 -2663
rect 1130 -2727 1138 -2675
rect 1190 -2727 1198 -2675
rect 1130 -2739 1198 -2727
rect 1130 -2791 1138 -2739
rect 1190 -2791 1198 -2739
rect 1130 -2803 1198 -2791
rect 1130 -2855 1138 -2803
rect 1190 -2855 1198 -2803
rect 1130 -2867 1198 -2855
rect 1130 -2919 1138 -2867
rect 1190 -2919 1198 -2867
rect 1130 -2931 1198 -2919
rect 1130 -2983 1138 -2931
rect 1190 -2983 1198 -2931
rect 1130 -2995 1198 -2983
rect 1130 -3047 1138 -2995
rect 1190 -3047 1198 -2995
rect 1130 -3059 1198 -3047
rect 1130 -3111 1138 -3059
rect 1190 -3111 1198 -3059
rect 1130 -3123 1198 -3111
rect 1130 -3175 1138 -3123
rect 1190 -3175 1198 -3123
rect 1130 -3196 1198 -3175
rect 1588 -563 1656 -542
rect 1588 -615 1596 -563
rect 1648 -615 1656 -563
rect 1588 -627 1656 -615
rect 1588 -679 1596 -627
rect 1648 -679 1656 -627
rect 1588 -691 1656 -679
rect 1588 -743 1596 -691
rect 1648 -743 1656 -691
rect 1588 -755 1656 -743
rect 1588 -807 1596 -755
rect 1648 -807 1656 -755
rect 1588 -819 1656 -807
rect 1588 -871 1596 -819
rect 1648 -871 1656 -819
rect 1588 -883 1656 -871
rect 1588 -935 1596 -883
rect 1648 -935 1656 -883
rect 1588 -947 1656 -935
rect 1588 -999 1596 -947
rect 1648 -999 1656 -947
rect 1588 -1011 1656 -999
rect 1588 -1063 1596 -1011
rect 1648 -1063 1656 -1011
rect 1588 -1075 1656 -1063
rect 1588 -1127 1596 -1075
rect 1648 -1127 1656 -1075
rect 1588 -1139 1656 -1127
rect 1588 -1191 1596 -1139
rect 1648 -1191 1656 -1139
rect 1588 -1203 1656 -1191
rect 1588 -1255 1596 -1203
rect 1648 -1255 1656 -1203
rect 1588 -1267 1656 -1255
rect 1588 -1319 1596 -1267
rect 1648 -1319 1656 -1267
rect 1588 -1331 1656 -1319
rect 1588 -1383 1596 -1331
rect 1648 -1383 1656 -1331
rect 1588 -1395 1656 -1383
rect 1588 -1447 1596 -1395
rect 1648 -1447 1656 -1395
rect 1588 -1459 1656 -1447
rect 1588 -1511 1596 -1459
rect 1648 -1511 1656 -1459
rect 1588 -1523 1656 -1511
rect 1588 -1575 1596 -1523
rect 1648 -1575 1656 -1523
rect 1588 -1587 1656 -1575
rect 1588 -1639 1596 -1587
rect 1648 -1639 1656 -1587
rect 1588 -1651 1656 -1639
rect 1588 -1703 1596 -1651
rect 1648 -1703 1656 -1651
rect 1588 -1715 1656 -1703
rect 1588 -1767 1596 -1715
rect 1648 -1767 1656 -1715
rect 1588 -1779 1656 -1767
rect 1588 -1831 1596 -1779
rect 1648 -1831 1656 -1779
rect 1588 -1843 1656 -1831
rect 1588 -1895 1596 -1843
rect 1648 -1895 1656 -1843
rect 1588 -1907 1656 -1895
rect 1588 -1959 1596 -1907
rect 1648 -1959 1656 -1907
rect 1588 -1971 1656 -1959
rect 1588 -2023 1596 -1971
rect 1648 -2023 1656 -1971
rect 1588 -2035 1656 -2023
rect 1588 -2087 1596 -2035
rect 1648 -2087 1656 -2035
rect 1588 -2099 1656 -2087
rect 1588 -2151 1596 -2099
rect 1648 -2151 1656 -2099
rect 1588 -2163 1656 -2151
rect 1588 -2215 1596 -2163
rect 1648 -2215 1656 -2163
rect 1588 -2227 1656 -2215
rect 1588 -2279 1596 -2227
rect 1648 -2279 1656 -2227
rect 1588 -2291 1656 -2279
rect 1588 -2343 1596 -2291
rect 1648 -2343 1656 -2291
rect 1588 -2355 1656 -2343
rect 1588 -2407 1596 -2355
rect 1648 -2407 1656 -2355
rect 1588 -2419 1656 -2407
rect 1588 -2471 1596 -2419
rect 1648 -2471 1656 -2419
rect 1588 -2483 1656 -2471
rect 1588 -2535 1596 -2483
rect 1648 -2535 1656 -2483
rect 1588 -2547 1656 -2535
rect 1588 -2599 1596 -2547
rect 1648 -2599 1656 -2547
rect 1588 -2611 1656 -2599
rect 1588 -2663 1596 -2611
rect 1648 -2663 1656 -2611
rect 1588 -2675 1656 -2663
rect 1588 -2727 1596 -2675
rect 1648 -2727 1656 -2675
rect 1588 -2739 1656 -2727
rect 1588 -2791 1596 -2739
rect 1648 -2791 1656 -2739
rect 1588 -2803 1656 -2791
rect 1588 -2855 1596 -2803
rect 1648 -2855 1656 -2803
rect 1588 -2867 1656 -2855
rect 1588 -2919 1596 -2867
rect 1648 -2919 1656 -2867
rect 1588 -2931 1656 -2919
rect 1588 -2983 1596 -2931
rect 1648 -2983 1656 -2931
rect 1588 -2995 1656 -2983
rect 1588 -3047 1596 -2995
rect 1648 -3047 1656 -2995
rect 1588 -3059 1656 -3047
rect 1588 -3111 1596 -3059
rect 1648 -3111 1656 -3059
rect 1588 -3123 1656 -3111
rect 1588 -3175 1596 -3123
rect 1648 -3175 1656 -3123
rect 1588 -3196 1656 -3175
rect 2046 -563 2114 -542
rect 2046 -615 2054 -563
rect 2106 -615 2114 -563
rect 2046 -627 2114 -615
rect 2046 -679 2054 -627
rect 2106 -679 2114 -627
rect 2046 -691 2114 -679
rect 2046 -743 2054 -691
rect 2106 -743 2114 -691
rect 2046 -755 2114 -743
rect 2046 -807 2054 -755
rect 2106 -807 2114 -755
rect 2046 -819 2114 -807
rect 2046 -871 2054 -819
rect 2106 -871 2114 -819
rect 2046 -883 2114 -871
rect 2046 -935 2054 -883
rect 2106 -935 2114 -883
rect 2046 -947 2114 -935
rect 2046 -999 2054 -947
rect 2106 -999 2114 -947
rect 2046 -1011 2114 -999
rect 2046 -1063 2054 -1011
rect 2106 -1063 2114 -1011
rect 2046 -1075 2114 -1063
rect 2046 -1127 2054 -1075
rect 2106 -1127 2114 -1075
rect 2046 -1139 2114 -1127
rect 2046 -1191 2054 -1139
rect 2106 -1191 2114 -1139
rect 2046 -1203 2114 -1191
rect 2046 -1255 2054 -1203
rect 2106 -1255 2114 -1203
rect 2046 -1267 2114 -1255
rect 2046 -1319 2054 -1267
rect 2106 -1319 2114 -1267
rect 2046 -1331 2114 -1319
rect 2046 -1383 2054 -1331
rect 2106 -1383 2114 -1331
rect 2046 -1395 2114 -1383
rect 2046 -1447 2054 -1395
rect 2106 -1447 2114 -1395
rect 2046 -1459 2114 -1447
rect 2046 -1511 2054 -1459
rect 2106 -1511 2114 -1459
rect 2046 -1523 2114 -1511
rect 2046 -1575 2054 -1523
rect 2106 -1575 2114 -1523
rect 2046 -1587 2114 -1575
rect 2046 -1639 2054 -1587
rect 2106 -1639 2114 -1587
rect 2046 -1651 2114 -1639
rect 2046 -1703 2054 -1651
rect 2106 -1703 2114 -1651
rect 2046 -1715 2114 -1703
rect 2046 -1767 2054 -1715
rect 2106 -1767 2114 -1715
rect 2046 -1779 2114 -1767
rect 2046 -1831 2054 -1779
rect 2106 -1831 2114 -1779
rect 2046 -1843 2114 -1831
rect 2046 -1895 2054 -1843
rect 2106 -1895 2114 -1843
rect 2046 -1907 2114 -1895
rect 2046 -1959 2054 -1907
rect 2106 -1959 2114 -1907
rect 2046 -1971 2114 -1959
rect 2046 -2023 2054 -1971
rect 2106 -2023 2114 -1971
rect 2046 -2035 2114 -2023
rect 2046 -2087 2054 -2035
rect 2106 -2087 2114 -2035
rect 2046 -2099 2114 -2087
rect 2046 -2151 2054 -2099
rect 2106 -2151 2114 -2099
rect 2046 -2163 2114 -2151
rect 2046 -2215 2054 -2163
rect 2106 -2215 2114 -2163
rect 2046 -2227 2114 -2215
rect 2046 -2279 2054 -2227
rect 2106 -2279 2114 -2227
rect 2046 -2291 2114 -2279
rect 2046 -2343 2054 -2291
rect 2106 -2343 2114 -2291
rect 2046 -2355 2114 -2343
rect 2046 -2407 2054 -2355
rect 2106 -2407 2114 -2355
rect 2046 -2419 2114 -2407
rect 2046 -2471 2054 -2419
rect 2106 -2471 2114 -2419
rect 2046 -2483 2114 -2471
rect 2046 -2535 2054 -2483
rect 2106 -2535 2114 -2483
rect 2046 -2547 2114 -2535
rect 2046 -2599 2054 -2547
rect 2106 -2599 2114 -2547
rect 2046 -2611 2114 -2599
rect 2046 -2663 2054 -2611
rect 2106 -2663 2114 -2611
rect 2046 -2675 2114 -2663
rect 2046 -2727 2054 -2675
rect 2106 -2727 2114 -2675
rect 2046 -2739 2114 -2727
rect 2046 -2791 2054 -2739
rect 2106 -2791 2114 -2739
rect 2046 -2803 2114 -2791
rect 2046 -2855 2054 -2803
rect 2106 -2855 2114 -2803
rect 2046 -2867 2114 -2855
rect 2046 -2919 2054 -2867
rect 2106 -2919 2114 -2867
rect 2046 -2931 2114 -2919
rect 2046 -2983 2054 -2931
rect 2106 -2983 2114 -2931
rect 2046 -2995 2114 -2983
rect 2046 -3047 2054 -2995
rect 2106 -3047 2114 -2995
rect 2046 -3059 2114 -3047
rect 2046 -3111 2054 -3059
rect 2106 -3111 2114 -3059
rect 2046 -3123 2114 -3111
rect 2046 -3175 2054 -3123
rect 2106 -3175 2114 -3123
rect 2046 -3196 2114 -3175
rect 2504 -563 2572 -542
rect 2504 -615 2512 -563
rect 2564 -615 2572 -563
rect 2504 -627 2572 -615
rect 2504 -679 2512 -627
rect 2564 -679 2572 -627
rect 2504 -691 2572 -679
rect 2504 -743 2512 -691
rect 2564 -743 2572 -691
rect 2504 -755 2572 -743
rect 2504 -807 2512 -755
rect 2564 -807 2572 -755
rect 2504 -819 2572 -807
rect 2504 -871 2512 -819
rect 2564 -871 2572 -819
rect 2504 -883 2572 -871
rect 2504 -935 2512 -883
rect 2564 -935 2572 -883
rect 2504 -947 2572 -935
rect 2504 -999 2512 -947
rect 2564 -999 2572 -947
rect 2504 -1011 2572 -999
rect 2504 -1063 2512 -1011
rect 2564 -1063 2572 -1011
rect 2504 -1075 2572 -1063
rect 2504 -1127 2512 -1075
rect 2564 -1127 2572 -1075
rect 2504 -1139 2572 -1127
rect 2504 -1191 2512 -1139
rect 2564 -1191 2572 -1139
rect 2504 -1203 2572 -1191
rect 2504 -1255 2512 -1203
rect 2564 -1255 2572 -1203
rect 2504 -1267 2572 -1255
rect 2504 -1319 2512 -1267
rect 2564 -1319 2572 -1267
rect 2504 -1331 2572 -1319
rect 2504 -1383 2512 -1331
rect 2564 -1383 2572 -1331
rect 2504 -1395 2572 -1383
rect 2504 -1447 2512 -1395
rect 2564 -1447 2572 -1395
rect 2504 -1459 2572 -1447
rect 2504 -1511 2512 -1459
rect 2564 -1511 2572 -1459
rect 2504 -1523 2572 -1511
rect 2504 -1575 2512 -1523
rect 2564 -1575 2572 -1523
rect 2504 -1587 2572 -1575
rect 2504 -1639 2512 -1587
rect 2564 -1639 2572 -1587
rect 2504 -1651 2572 -1639
rect 2504 -1703 2512 -1651
rect 2564 -1703 2572 -1651
rect 2504 -1715 2572 -1703
rect 2504 -1767 2512 -1715
rect 2564 -1767 2572 -1715
rect 2504 -1779 2572 -1767
rect 2504 -1831 2512 -1779
rect 2564 -1831 2572 -1779
rect 2504 -1843 2572 -1831
rect 2504 -1895 2512 -1843
rect 2564 -1895 2572 -1843
rect 2504 -1907 2572 -1895
rect 2504 -1959 2512 -1907
rect 2564 -1959 2572 -1907
rect 2504 -1971 2572 -1959
rect 2504 -2023 2512 -1971
rect 2564 -2023 2572 -1971
rect 2504 -2035 2572 -2023
rect 2504 -2087 2512 -2035
rect 2564 -2087 2572 -2035
rect 2504 -2099 2572 -2087
rect 2504 -2151 2512 -2099
rect 2564 -2151 2572 -2099
rect 2504 -2163 2572 -2151
rect 2504 -2215 2512 -2163
rect 2564 -2215 2572 -2163
rect 2504 -2227 2572 -2215
rect 2504 -2279 2512 -2227
rect 2564 -2279 2572 -2227
rect 2504 -2291 2572 -2279
rect 2504 -2343 2512 -2291
rect 2564 -2343 2572 -2291
rect 2504 -2355 2572 -2343
rect 2504 -2407 2512 -2355
rect 2564 -2407 2572 -2355
rect 2504 -2419 2572 -2407
rect 2504 -2471 2512 -2419
rect 2564 -2471 2572 -2419
rect 2504 -2483 2572 -2471
rect 2504 -2535 2512 -2483
rect 2564 -2535 2572 -2483
rect 2504 -2547 2572 -2535
rect 2504 -2599 2512 -2547
rect 2564 -2599 2572 -2547
rect 2504 -2611 2572 -2599
rect 2504 -2663 2512 -2611
rect 2564 -2663 2572 -2611
rect 2504 -2675 2572 -2663
rect 2504 -2727 2512 -2675
rect 2564 -2727 2572 -2675
rect 2504 -2739 2572 -2727
rect 2504 -2791 2512 -2739
rect 2564 -2791 2572 -2739
rect 2504 -2803 2572 -2791
rect 2504 -2855 2512 -2803
rect 2564 -2855 2572 -2803
rect 2504 -2867 2572 -2855
rect 2504 -2919 2512 -2867
rect 2564 -2919 2572 -2867
rect 2504 -2931 2572 -2919
rect 2504 -2983 2512 -2931
rect 2564 -2983 2572 -2931
rect 2504 -2995 2572 -2983
rect 2504 -3047 2512 -2995
rect 2564 -3047 2572 -2995
rect 2504 -3059 2572 -3047
rect 2504 -3111 2512 -3059
rect 2564 -3111 2572 -3059
rect 2504 -3123 2572 -3111
rect 2504 -3175 2512 -3123
rect 2564 -3175 2572 -3123
rect 2504 -3196 2572 -3175
rect 2962 -563 3030 -542
rect 2962 -615 2970 -563
rect 3022 -615 3030 -563
rect 2962 -627 3030 -615
rect 2962 -679 2970 -627
rect 3022 -679 3030 -627
rect 2962 -691 3030 -679
rect 2962 -743 2970 -691
rect 3022 -743 3030 -691
rect 2962 -755 3030 -743
rect 2962 -807 2970 -755
rect 3022 -807 3030 -755
rect 2962 -819 3030 -807
rect 2962 -871 2970 -819
rect 3022 -871 3030 -819
rect 2962 -883 3030 -871
rect 2962 -935 2970 -883
rect 3022 -935 3030 -883
rect 2962 -947 3030 -935
rect 2962 -999 2970 -947
rect 3022 -999 3030 -947
rect 2962 -1011 3030 -999
rect 2962 -1063 2970 -1011
rect 3022 -1063 3030 -1011
rect 2962 -1075 3030 -1063
rect 2962 -1127 2970 -1075
rect 3022 -1127 3030 -1075
rect 2962 -1139 3030 -1127
rect 2962 -1191 2970 -1139
rect 3022 -1191 3030 -1139
rect 2962 -1203 3030 -1191
rect 2962 -1255 2970 -1203
rect 3022 -1255 3030 -1203
rect 2962 -1267 3030 -1255
rect 2962 -1319 2970 -1267
rect 3022 -1319 3030 -1267
rect 2962 -1331 3030 -1319
rect 2962 -1383 2970 -1331
rect 3022 -1383 3030 -1331
rect 2962 -1395 3030 -1383
rect 2962 -1447 2970 -1395
rect 3022 -1447 3030 -1395
rect 2962 -1459 3030 -1447
rect 2962 -1511 2970 -1459
rect 3022 -1511 3030 -1459
rect 2962 -1523 3030 -1511
rect 2962 -1575 2970 -1523
rect 3022 -1575 3030 -1523
rect 2962 -1587 3030 -1575
rect 2962 -1639 2970 -1587
rect 3022 -1639 3030 -1587
rect 2962 -1651 3030 -1639
rect 2962 -1703 2970 -1651
rect 3022 -1703 3030 -1651
rect 2962 -1715 3030 -1703
rect 2962 -1767 2970 -1715
rect 3022 -1767 3030 -1715
rect 2962 -1779 3030 -1767
rect 2962 -1831 2970 -1779
rect 3022 -1831 3030 -1779
rect 2962 -1843 3030 -1831
rect 2962 -1895 2970 -1843
rect 3022 -1895 3030 -1843
rect 2962 -1907 3030 -1895
rect 2962 -1959 2970 -1907
rect 3022 -1959 3030 -1907
rect 2962 -1971 3030 -1959
rect 2962 -2023 2970 -1971
rect 3022 -2023 3030 -1971
rect 2962 -2035 3030 -2023
rect 2962 -2087 2970 -2035
rect 3022 -2087 3030 -2035
rect 2962 -2099 3030 -2087
rect 2962 -2151 2970 -2099
rect 3022 -2151 3030 -2099
rect 2962 -2163 3030 -2151
rect 2962 -2215 2970 -2163
rect 3022 -2215 3030 -2163
rect 2962 -2227 3030 -2215
rect 2962 -2279 2970 -2227
rect 3022 -2279 3030 -2227
rect 2962 -2291 3030 -2279
rect 2962 -2343 2970 -2291
rect 3022 -2343 3030 -2291
rect 2962 -2355 3030 -2343
rect 2962 -2407 2970 -2355
rect 3022 -2407 3030 -2355
rect 2962 -2419 3030 -2407
rect 2962 -2471 2970 -2419
rect 3022 -2471 3030 -2419
rect 2962 -2483 3030 -2471
rect 2962 -2535 2970 -2483
rect 3022 -2535 3030 -2483
rect 2962 -2547 3030 -2535
rect 2962 -2599 2970 -2547
rect 3022 -2599 3030 -2547
rect 2962 -2611 3030 -2599
rect 2962 -2663 2970 -2611
rect 3022 -2663 3030 -2611
rect 2962 -2675 3030 -2663
rect 2962 -2727 2970 -2675
rect 3022 -2727 3030 -2675
rect 2962 -2739 3030 -2727
rect 2962 -2791 2970 -2739
rect 3022 -2791 3030 -2739
rect 2962 -2803 3030 -2791
rect 2962 -2855 2970 -2803
rect 3022 -2855 3030 -2803
rect 2962 -2867 3030 -2855
rect 2962 -2919 2970 -2867
rect 3022 -2919 3030 -2867
rect 2962 -2931 3030 -2919
rect 2962 -2983 2970 -2931
rect 3022 -2983 3030 -2931
rect 2962 -2995 3030 -2983
rect 2962 -3047 2970 -2995
rect 3022 -3047 3030 -2995
rect 2962 -3059 3030 -3047
rect 2962 -3111 2970 -3059
rect 3022 -3111 3030 -3059
rect 2962 -3123 3030 -3111
rect 2962 -3175 2970 -3123
rect 3022 -3175 3030 -3123
rect 2962 -3196 3030 -3175
rect 3420 -563 3488 -542
rect 3420 -615 3428 -563
rect 3480 -615 3488 -563
rect 3420 -627 3488 -615
rect 3420 -679 3428 -627
rect 3480 -679 3488 -627
rect 3420 -691 3488 -679
rect 3420 -743 3428 -691
rect 3480 -743 3488 -691
rect 3420 -755 3488 -743
rect 3420 -807 3428 -755
rect 3480 -807 3488 -755
rect 3420 -819 3488 -807
rect 3420 -871 3428 -819
rect 3480 -871 3488 -819
rect 3420 -883 3488 -871
rect 3420 -935 3428 -883
rect 3480 -935 3488 -883
rect 3420 -947 3488 -935
rect 3420 -999 3428 -947
rect 3480 -999 3488 -947
rect 3420 -1011 3488 -999
rect 3420 -1063 3428 -1011
rect 3480 -1063 3488 -1011
rect 3420 -1075 3488 -1063
rect 3420 -1127 3428 -1075
rect 3480 -1127 3488 -1075
rect 3420 -1139 3488 -1127
rect 3420 -1191 3428 -1139
rect 3480 -1191 3488 -1139
rect 3420 -1203 3488 -1191
rect 3420 -1255 3428 -1203
rect 3480 -1255 3488 -1203
rect 3420 -1267 3488 -1255
rect 3420 -1319 3428 -1267
rect 3480 -1319 3488 -1267
rect 3420 -1331 3488 -1319
rect 3420 -1383 3428 -1331
rect 3480 -1383 3488 -1331
rect 3420 -1395 3488 -1383
rect 3420 -1447 3428 -1395
rect 3480 -1447 3488 -1395
rect 3420 -1459 3488 -1447
rect 3420 -1511 3428 -1459
rect 3480 -1511 3488 -1459
rect 3420 -1523 3488 -1511
rect 3420 -1575 3428 -1523
rect 3480 -1575 3488 -1523
rect 3420 -1587 3488 -1575
rect 3420 -1639 3428 -1587
rect 3480 -1639 3488 -1587
rect 3420 -1651 3488 -1639
rect 3420 -1703 3428 -1651
rect 3480 -1703 3488 -1651
rect 3420 -1715 3488 -1703
rect 3420 -1767 3428 -1715
rect 3480 -1767 3488 -1715
rect 3420 -1779 3488 -1767
rect 3420 -1831 3428 -1779
rect 3480 -1831 3488 -1779
rect 3420 -1843 3488 -1831
rect 3420 -1895 3428 -1843
rect 3480 -1895 3488 -1843
rect 3420 -1907 3488 -1895
rect 3420 -1959 3428 -1907
rect 3480 -1959 3488 -1907
rect 3420 -1971 3488 -1959
rect 3420 -2023 3428 -1971
rect 3480 -2023 3488 -1971
rect 3420 -2035 3488 -2023
rect 3420 -2087 3428 -2035
rect 3480 -2087 3488 -2035
rect 3420 -2099 3488 -2087
rect 3420 -2151 3428 -2099
rect 3480 -2151 3488 -2099
rect 3420 -2163 3488 -2151
rect 3420 -2215 3428 -2163
rect 3480 -2215 3488 -2163
rect 3420 -2227 3488 -2215
rect 3420 -2279 3428 -2227
rect 3480 -2279 3488 -2227
rect 3420 -2291 3488 -2279
rect 3420 -2343 3428 -2291
rect 3480 -2343 3488 -2291
rect 3420 -2355 3488 -2343
rect 3420 -2407 3428 -2355
rect 3480 -2407 3488 -2355
rect 3420 -2419 3488 -2407
rect 3420 -2471 3428 -2419
rect 3480 -2471 3488 -2419
rect 3420 -2483 3488 -2471
rect 3420 -2535 3428 -2483
rect 3480 -2535 3488 -2483
rect 3420 -2547 3488 -2535
rect 3420 -2599 3428 -2547
rect 3480 -2599 3488 -2547
rect 3420 -2611 3488 -2599
rect 3420 -2663 3428 -2611
rect 3480 -2663 3488 -2611
rect 3420 -2675 3488 -2663
rect 3420 -2727 3428 -2675
rect 3480 -2727 3488 -2675
rect 3420 -2739 3488 -2727
rect 3420 -2791 3428 -2739
rect 3480 -2791 3488 -2739
rect 3420 -2803 3488 -2791
rect 3420 -2855 3428 -2803
rect 3480 -2855 3488 -2803
rect 3420 -2867 3488 -2855
rect 3420 -2919 3428 -2867
rect 3480 -2919 3488 -2867
rect 3420 -2931 3488 -2919
rect 3420 -2983 3428 -2931
rect 3480 -2983 3488 -2931
rect 3420 -2995 3488 -2983
rect 3420 -3047 3428 -2995
rect 3480 -3047 3488 -2995
rect 3420 -3059 3488 -3047
rect 3420 -3111 3428 -3059
rect 3480 -3111 3488 -3059
rect 3420 -3123 3488 -3111
rect 3420 -3175 3428 -3123
rect 3480 -3175 3488 -3123
rect 3420 -3196 3488 -3175
rect -950 -3224 -845 -3209
rect -1401 -3228 -845 -3224
rect -1401 -3262 -915 -3228
rect -881 -3262 -845 -3228
rect -1401 -3277 -845 -3262
rect -1401 -3292 -935 -3277
rect -691 -3324 -645 -3196
rect 225 -3324 271 -3196
rect 1141 -3324 1187 -3196
rect 2057 -3326 2103 -3196
rect 2973 -3326 3019 -3196
<< via1 >>
rect -1200 6574 -1148 6605
rect -1200 6553 -1191 6574
rect -1191 6553 -1157 6574
rect -1157 6553 -1148 6574
rect -1136 6574 -1084 6605
rect -1136 6553 -1119 6574
rect -1119 6553 -1085 6574
rect -1085 6553 -1084 6574
rect -1072 6574 -1020 6605
rect -1008 6574 -956 6605
rect -944 6574 -892 6605
rect -880 6574 -828 6605
rect -816 6574 -764 6605
rect -752 6574 -700 6605
rect -1072 6553 -1047 6574
rect -1047 6553 -1020 6574
rect -1008 6553 -975 6574
rect -975 6553 -956 6574
rect -944 6553 -941 6574
rect -941 6553 -903 6574
rect -903 6553 -892 6574
rect -880 6553 -869 6574
rect -869 6553 -831 6574
rect -831 6553 -828 6574
rect -816 6553 -797 6574
rect -797 6553 -764 6574
rect -752 6553 -725 6574
rect -725 6553 -700 6574
rect -688 6574 -636 6605
rect -688 6553 -687 6574
rect -687 6553 -653 6574
rect -653 6553 -636 6574
rect -624 6574 -572 6605
rect -624 6553 -615 6574
rect -615 6553 -581 6574
rect -581 6553 -572 6574
rect -560 6574 -508 6605
rect -560 6553 -543 6574
rect -543 6553 -509 6574
rect -509 6553 -508 6574
rect -496 6574 -444 6605
rect -432 6574 -380 6605
rect -368 6574 -316 6605
rect -304 6574 -252 6605
rect -240 6574 -188 6605
rect -176 6574 -124 6605
rect -496 6553 -471 6574
rect -471 6553 -444 6574
rect -432 6553 -399 6574
rect -399 6553 -380 6574
rect -368 6553 -365 6574
rect -365 6553 -327 6574
rect -327 6553 -316 6574
rect -304 6553 -293 6574
rect -293 6553 -255 6574
rect -255 6553 -252 6574
rect -240 6553 -221 6574
rect -221 6553 -188 6574
rect -176 6553 -149 6574
rect -149 6553 -124 6574
rect -112 6574 -60 6605
rect -112 6553 -111 6574
rect -111 6553 -77 6574
rect -77 6553 -60 6574
rect -48 6574 4 6605
rect -48 6553 -39 6574
rect -39 6553 -5 6574
rect -5 6553 4 6574
rect 16 6574 68 6605
rect 16 6553 33 6574
rect 33 6553 67 6574
rect 67 6553 68 6574
rect 80 6574 132 6605
rect 144 6574 196 6605
rect 208 6574 260 6605
rect 272 6574 324 6605
rect 336 6574 388 6605
rect 400 6574 452 6605
rect 80 6553 105 6574
rect 105 6553 132 6574
rect 144 6553 177 6574
rect 177 6553 196 6574
rect 208 6553 211 6574
rect 211 6553 249 6574
rect 249 6553 260 6574
rect 272 6553 283 6574
rect 283 6553 321 6574
rect 321 6553 324 6574
rect 336 6553 355 6574
rect 355 6553 388 6574
rect 400 6553 427 6574
rect 427 6553 452 6574
rect 464 6574 516 6605
rect 464 6553 465 6574
rect 465 6553 499 6574
rect 499 6553 516 6574
rect 528 6574 580 6605
rect 528 6553 537 6574
rect 537 6553 571 6574
rect 571 6553 580 6574
rect 592 6574 644 6605
rect 592 6553 609 6574
rect 609 6553 643 6574
rect 643 6553 644 6574
rect 656 6574 708 6605
rect 720 6574 772 6605
rect 784 6574 836 6605
rect 848 6574 900 6605
rect 912 6574 964 6605
rect 976 6574 1028 6605
rect 656 6553 681 6574
rect 681 6553 708 6574
rect 720 6553 753 6574
rect 753 6553 772 6574
rect 784 6553 787 6574
rect 787 6553 825 6574
rect 825 6553 836 6574
rect 848 6553 859 6574
rect 859 6553 897 6574
rect 897 6553 900 6574
rect 912 6553 931 6574
rect 931 6553 964 6574
rect 976 6553 1003 6574
rect 1003 6553 1028 6574
rect 1040 6574 1092 6605
rect 1040 6553 1041 6574
rect 1041 6553 1075 6574
rect 1075 6553 1092 6574
rect 1104 6574 1156 6605
rect 1104 6553 1113 6574
rect 1113 6553 1147 6574
rect 1147 6553 1156 6574
rect 1168 6553 1220 6605
rect 1232 6553 1284 6605
rect 1296 6553 1348 6605
rect 1360 6553 1412 6605
rect 1424 6574 1476 6605
rect 1424 6553 1433 6574
rect 1433 6553 1467 6574
rect 1467 6553 1476 6574
rect 1488 6574 1540 6605
rect 1488 6553 1505 6574
rect 1505 6553 1539 6574
rect 1539 6553 1540 6574
rect 1552 6574 1604 6605
rect 1616 6574 1668 6605
rect 1680 6574 1732 6605
rect 1744 6574 1796 6605
rect 1808 6574 1860 6605
rect 1872 6574 1924 6605
rect 1552 6553 1577 6574
rect 1577 6553 1604 6574
rect 1616 6553 1649 6574
rect 1649 6553 1668 6574
rect 1680 6553 1683 6574
rect 1683 6553 1721 6574
rect 1721 6553 1732 6574
rect 1744 6553 1755 6574
rect 1755 6553 1793 6574
rect 1793 6553 1796 6574
rect 1808 6553 1827 6574
rect 1827 6553 1860 6574
rect 1872 6553 1899 6574
rect 1899 6553 1924 6574
rect 1936 6574 1988 6605
rect 1936 6553 1937 6574
rect 1937 6553 1971 6574
rect 1971 6553 1988 6574
rect 2000 6574 2052 6605
rect 2000 6553 2009 6574
rect 2009 6553 2043 6574
rect 2043 6553 2052 6574
rect 2064 6574 2116 6605
rect 2064 6553 2081 6574
rect 2081 6553 2115 6574
rect 2115 6553 2116 6574
rect 2128 6574 2180 6605
rect 2192 6574 2244 6605
rect 2256 6574 2308 6605
rect 2320 6574 2372 6605
rect 2384 6574 2436 6605
rect 2448 6574 2500 6605
rect 2128 6553 2153 6574
rect 2153 6553 2180 6574
rect 2192 6553 2225 6574
rect 2225 6553 2244 6574
rect 2256 6553 2259 6574
rect 2259 6553 2297 6574
rect 2297 6553 2308 6574
rect 2320 6553 2331 6574
rect 2331 6553 2369 6574
rect 2369 6553 2372 6574
rect 2384 6553 2403 6574
rect 2403 6553 2436 6574
rect 2448 6553 2475 6574
rect 2475 6553 2500 6574
rect 2512 6574 2564 6605
rect 2512 6553 2513 6574
rect 2513 6553 2547 6574
rect 2547 6553 2564 6574
rect 2576 6574 2628 6605
rect 2576 6553 2585 6574
rect 2585 6553 2619 6574
rect 2619 6553 2628 6574
rect 2640 6574 2692 6605
rect 2640 6553 2657 6574
rect 2657 6553 2691 6574
rect 2691 6553 2692 6574
rect 2704 6574 2756 6605
rect 2768 6574 2820 6605
rect 2832 6574 2884 6605
rect 2896 6574 2948 6605
rect 2960 6574 3012 6605
rect 3024 6574 3076 6605
rect 2704 6553 2729 6574
rect 2729 6553 2756 6574
rect 2768 6553 2801 6574
rect 2801 6553 2820 6574
rect 2832 6553 2835 6574
rect 2835 6553 2873 6574
rect 2873 6553 2884 6574
rect 2896 6553 2907 6574
rect 2907 6553 2945 6574
rect 2945 6553 2948 6574
rect 2960 6553 2979 6574
rect 2979 6553 3012 6574
rect 3024 6553 3051 6574
rect 3051 6553 3076 6574
rect 3088 6574 3140 6605
rect 3088 6553 3089 6574
rect 3089 6553 3123 6574
rect 3123 6553 3140 6574
rect 3152 6574 3204 6605
rect 3152 6553 3161 6574
rect 3161 6553 3195 6574
rect 3195 6553 3204 6574
rect 3216 6574 3268 6605
rect 3216 6553 3233 6574
rect 3233 6553 3267 6574
rect 3267 6553 3268 6574
rect 3280 6574 3332 6605
rect 3344 6574 3396 6605
rect 3408 6574 3460 6605
rect 3472 6574 3524 6605
rect 3536 6574 3588 6605
rect 3600 6574 3652 6605
rect 3280 6553 3305 6574
rect 3305 6553 3332 6574
rect 3344 6553 3377 6574
rect 3377 6553 3396 6574
rect 3408 6553 3411 6574
rect 3411 6553 3449 6574
rect 3449 6553 3460 6574
rect 3472 6553 3483 6574
rect 3483 6553 3521 6574
rect 3521 6553 3524 6574
rect 3536 6553 3555 6574
rect 3555 6553 3588 6574
rect 3600 6553 3627 6574
rect 3627 6553 3652 6574
rect 3664 6574 3716 6605
rect 3664 6553 3665 6574
rect 3665 6553 3699 6574
rect 3699 6553 3716 6574
rect 3728 6574 3780 6605
rect 3728 6553 3737 6574
rect 3737 6553 3771 6574
rect 3771 6553 3780 6574
rect -735 6364 -683 6385
rect -735 6333 -726 6364
rect -726 6333 -692 6364
rect -692 6333 -683 6364
rect -735 6292 -683 6321
rect -735 6269 -726 6292
rect -726 6269 -692 6292
rect -692 6269 -683 6292
rect -735 6220 -683 6257
rect -735 6205 -726 6220
rect -726 6205 -692 6220
rect -692 6205 -683 6220
rect -735 6186 -726 6193
rect -726 6186 -692 6193
rect -692 6186 -683 6193
rect -735 6148 -683 6186
rect -735 6141 -726 6148
rect -726 6141 -692 6148
rect -692 6141 -683 6148
rect -735 6114 -726 6129
rect -726 6114 -692 6129
rect -692 6114 -683 6129
rect -735 6077 -683 6114
rect -735 6042 -726 6065
rect -726 6042 -692 6065
rect -692 6042 -683 6065
rect -735 6013 -683 6042
rect -735 5970 -726 6001
rect -726 5970 -692 6001
rect -692 5970 -683 6001
rect -735 5949 -683 5970
rect -735 5932 -683 5937
rect -735 5898 -726 5932
rect -726 5898 -692 5932
rect -692 5898 -683 5932
rect -735 5885 -683 5898
rect -735 5860 -683 5873
rect -735 5826 -726 5860
rect -726 5826 -692 5860
rect -692 5826 -683 5860
rect -735 5821 -683 5826
rect -735 5788 -683 5809
rect -735 5757 -726 5788
rect -726 5757 -692 5788
rect -692 5757 -683 5788
rect -735 5716 -683 5745
rect -735 5693 -726 5716
rect -726 5693 -692 5716
rect -692 5693 -683 5716
rect -735 5644 -683 5681
rect -735 5629 -726 5644
rect -726 5629 -692 5644
rect -692 5629 -683 5644
rect -735 5610 -726 5617
rect -726 5610 -692 5617
rect -692 5610 -683 5617
rect -735 5572 -683 5610
rect -735 5565 -726 5572
rect -726 5565 -692 5572
rect -692 5565 -683 5572
rect -735 5538 -726 5553
rect -726 5538 -692 5553
rect -692 5538 -683 5553
rect -735 5501 -683 5538
rect -735 5466 -726 5489
rect -726 5466 -692 5489
rect -692 5466 -683 5489
rect -735 5437 -683 5466
rect -735 5394 -726 5425
rect -726 5394 -692 5425
rect -692 5394 -683 5425
rect -735 5373 -683 5394
rect -735 5356 -683 5361
rect -735 5322 -726 5356
rect -726 5322 -692 5356
rect -692 5322 -683 5356
rect -735 5309 -683 5322
rect -735 5284 -683 5297
rect -735 5250 -726 5284
rect -726 5250 -692 5284
rect -692 5250 -683 5284
rect -735 5245 -683 5250
rect -735 5212 -683 5233
rect -735 5181 -726 5212
rect -726 5181 -692 5212
rect -692 5181 -683 5212
rect -735 5140 -683 5169
rect -735 5117 -726 5140
rect -726 5117 -692 5140
rect -692 5117 -683 5140
rect -735 5068 -683 5105
rect -735 5053 -726 5068
rect -726 5053 -692 5068
rect -692 5053 -683 5068
rect -735 5034 -726 5041
rect -726 5034 -692 5041
rect -692 5034 -683 5041
rect -735 4996 -683 5034
rect -735 4989 -726 4996
rect -726 4989 -692 4996
rect -692 4989 -683 4996
rect -735 4962 -726 4977
rect -726 4962 -692 4977
rect -692 4962 -683 4977
rect -735 4925 -683 4962
rect -735 4890 -726 4913
rect -726 4890 -692 4913
rect -692 4890 -683 4913
rect -735 4861 -683 4890
rect -735 4818 -726 4849
rect -726 4818 -692 4849
rect -692 4818 -683 4849
rect -735 4797 -683 4818
rect 181 6364 233 6385
rect 181 6333 190 6364
rect 190 6333 224 6364
rect 224 6333 233 6364
rect 181 6292 233 6321
rect 181 6269 190 6292
rect 190 6269 224 6292
rect 224 6269 233 6292
rect 181 6220 233 6257
rect 181 6205 190 6220
rect 190 6205 224 6220
rect 224 6205 233 6220
rect 181 6186 190 6193
rect 190 6186 224 6193
rect 224 6186 233 6193
rect 181 6148 233 6186
rect 181 6141 190 6148
rect 190 6141 224 6148
rect 224 6141 233 6148
rect 181 6114 190 6129
rect 190 6114 224 6129
rect 224 6114 233 6129
rect 181 6077 233 6114
rect 181 6042 190 6065
rect 190 6042 224 6065
rect 224 6042 233 6065
rect 181 6013 233 6042
rect 181 5970 190 6001
rect 190 5970 224 6001
rect 224 5970 233 6001
rect 181 5949 233 5970
rect 181 5932 233 5937
rect 181 5898 190 5932
rect 190 5898 224 5932
rect 224 5898 233 5932
rect 181 5885 233 5898
rect 181 5860 233 5873
rect 181 5826 190 5860
rect 190 5826 224 5860
rect 224 5826 233 5860
rect 181 5821 233 5826
rect 181 5788 233 5809
rect 181 5757 190 5788
rect 190 5757 224 5788
rect 224 5757 233 5788
rect 181 5716 233 5745
rect 181 5693 190 5716
rect 190 5693 224 5716
rect 224 5693 233 5716
rect 181 5644 233 5681
rect 181 5629 190 5644
rect 190 5629 224 5644
rect 224 5629 233 5644
rect 181 5610 190 5617
rect 190 5610 224 5617
rect 224 5610 233 5617
rect 181 5572 233 5610
rect 181 5565 190 5572
rect 190 5565 224 5572
rect 224 5565 233 5572
rect 181 5538 190 5553
rect 190 5538 224 5553
rect 224 5538 233 5553
rect 181 5501 233 5538
rect 181 5466 190 5489
rect 190 5466 224 5489
rect 224 5466 233 5489
rect 181 5437 233 5466
rect 181 5394 190 5425
rect 190 5394 224 5425
rect 224 5394 233 5425
rect 181 5373 233 5394
rect 181 5356 233 5361
rect 181 5322 190 5356
rect 190 5322 224 5356
rect 224 5322 233 5356
rect 181 5309 233 5322
rect 181 5284 233 5297
rect 181 5250 190 5284
rect 190 5250 224 5284
rect 224 5250 233 5284
rect 181 5245 233 5250
rect 181 5212 233 5233
rect 181 5181 190 5212
rect 190 5181 224 5212
rect 224 5181 233 5212
rect 181 5140 233 5169
rect 181 5117 190 5140
rect 190 5117 224 5140
rect 224 5117 233 5140
rect 181 5068 233 5105
rect 181 5053 190 5068
rect 190 5053 224 5068
rect 224 5053 233 5068
rect 181 5034 190 5041
rect 190 5034 224 5041
rect 224 5034 233 5041
rect 181 4996 233 5034
rect 181 4989 190 4996
rect 190 4989 224 4996
rect 224 4989 233 4996
rect 181 4962 190 4977
rect 190 4962 224 4977
rect 224 4962 233 4977
rect 181 4925 233 4962
rect 181 4890 190 4913
rect 190 4890 224 4913
rect 224 4890 233 4913
rect 181 4861 233 4890
rect 181 4818 190 4849
rect 190 4818 224 4849
rect 224 4818 233 4849
rect 181 4797 233 4818
rect 1097 6364 1149 6385
rect 1097 6333 1106 6364
rect 1106 6333 1140 6364
rect 1140 6333 1149 6364
rect 1097 6292 1149 6321
rect 1097 6269 1106 6292
rect 1106 6269 1140 6292
rect 1140 6269 1149 6292
rect 1097 6220 1149 6257
rect 1097 6205 1106 6220
rect 1106 6205 1140 6220
rect 1140 6205 1149 6220
rect 1097 6186 1106 6193
rect 1106 6186 1140 6193
rect 1140 6186 1149 6193
rect 1097 6148 1149 6186
rect 1097 6141 1106 6148
rect 1106 6141 1140 6148
rect 1140 6141 1149 6148
rect 1097 6114 1106 6129
rect 1106 6114 1140 6129
rect 1140 6114 1149 6129
rect 1097 6077 1149 6114
rect 1097 6042 1106 6065
rect 1106 6042 1140 6065
rect 1140 6042 1149 6065
rect 1097 6013 1149 6042
rect 1097 5970 1106 6001
rect 1106 5970 1140 6001
rect 1140 5970 1149 6001
rect 1097 5949 1149 5970
rect 1097 5932 1149 5937
rect 1097 5898 1106 5932
rect 1106 5898 1140 5932
rect 1140 5898 1149 5932
rect 1097 5885 1149 5898
rect 1097 5860 1149 5873
rect 1097 5826 1106 5860
rect 1106 5826 1140 5860
rect 1140 5826 1149 5860
rect 1097 5821 1149 5826
rect 1097 5788 1149 5809
rect 1097 5757 1106 5788
rect 1106 5757 1140 5788
rect 1140 5757 1149 5788
rect 1097 5716 1149 5745
rect 1097 5693 1106 5716
rect 1106 5693 1140 5716
rect 1140 5693 1149 5716
rect 1097 5644 1149 5681
rect 1097 5629 1106 5644
rect 1106 5629 1140 5644
rect 1140 5629 1149 5644
rect 1097 5610 1106 5617
rect 1106 5610 1140 5617
rect 1140 5610 1149 5617
rect 1097 5572 1149 5610
rect 1097 5565 1106 5572
rect 1106 5565 1140 5572
rect 1140 5565 1149 5572
rect 1097 5538 1106 5553
rect 1106 5538 1140 5553
rect 1140 5538 1149 5553
rect 1097 5501 1149 5538
rect 1097 5466 1106 5489
rect 1106 5466 1140 5489
rect 1140 5466 1149 5489
rect 1097 5437 1149 5466
rect 1097 5394 1106 5425
rect 1106 5394 1140 5425
rect 1140 5394 1149 5425
rect 1097 5373 1149 5394
rect 1097 5356 1149 5361
rect 1097 5322 1106 5356
rect 1106 5322 1140 5356
rect 1140 5322 1149 5356
rect 1097 5309 1149 5322
rect 1097 5284 1149 5297
rect 1097 5250 1106 5284
rect 1106 5250 1140 5284
rect 1140 5250 1149 5284
rect 1097 5245 1149 5250
rect 1097 5212 1149 5233
rect 1097 5181 1106 5212
rect 1106 5181 1140 5212
rect 1140 5181 1149 5212
rect 1097 5140 1149 5169
rect 1097 5117 1106 5140
rect 1106 5117 1140 5140
rect 1140 5117 1149 5140
rect 1097 5068 1149 5105
rect 1097 5053 1106 5068
rect 1106 5053 1140 5068
rect 1140 5053 1149 5068
rect 1097 5034 1106 5041
rect 1106 5034 1140 5041
rect 1140 5034 1149 5041
rect 1097 4996 1149 5034
rect 1097 4989 1106 4996
rect 1106 4989 1140 4996
rect 1140 4989 1149 4996
rect 1097 4962 1106 4977
rect 1106 4962 1140 4977
rect 1140 4962 1149 4977
rect 1097 4925 1149 4962
rect 1097 4890 1106 4913
rect 1106 4890 1140 4913
rect 1140 4890 1149 4913
rect 1097 4861 1149 4890
rect 1097 4818 1106 4849
rect 1106 4818 1140 4849
rect 1140 4818 1149 4849
rect 1097 4797 1149 4818
rect 1431 6333 1483 6385
rect 1431 6269 1483 6321
rect 1431 6205 1483 6257
rect 1431 6141 1483 6193
rect 1431 6077 1483 6129
rect 1431 6013 1483 6065
rect 1431 5949 1483 6001
rect 1431 5885 1483 5937
rect 1431 5821 1483 5873
rect 1431 5757 1483 5809
rect 1431 5693 1483 5745
rect 1431 5629 1483 5681
rect 1431 5565 1483 5617
rect 1431 5501 1483 5553
rect 1431 5437 1483 5489
rect 1431 5373 1483 5425
rect 1431 5309 1483 5361
rect 1431 5245 1483 5297
rect 1431 5181 1483 5233
rect 1431 5117 1483 5169
rect 1431 5053 1483 5105
rect 1431 4989 1483 5041
rect 1431 4925 1483 4977
rect 1431 4861 1483 4913
rect 1431 4797 1483 4849
rect 2347 6333 2399 6385
rect 2347 6269 2399 6321
rect 2347 6205 2399 6257
rect 2347 6141 2399 6193
rect 2347 6077 2399 6129
rect 2347 6013 2399 6065
rect 2347 5949 2399 6001
rect 2347 5885 2399 5937
rect 2347 5821 2399 5873
rect 2347 5757 2399 5809
rect 2347 5693 2399 5745
rect 2347 5629 2399 5681
rect 2347 5565 2399 5617
rect 2347 5501 2399 5553
rect 2347 5437 2399 5489
rect 2347 5373 2399 5425
rect 2347 5309 2399 5361
rect 2347 5245 2399 5297
rect 2347 5181 2399 5233
rect 2347 5117 2399 5169
rect 2347 5053 2399 5105
rect 2347 4989 2399 5041
rect 2347 4925 2399 4977
rect 2347 4861 2399 4913
rect 2347 4797 2399 4849
rect 3263 6333 3315 6385
rect 3263 6269 3315 6321
rect 3263 6205 3315 6257
rect 3263 6141 3315 6193
rect 3263 6077 3315 6129
rect 3263 6013 3315 6065
rect 3263 5949 3315 6001
rect 3263 5885 3315 5937
rect 3263 5821 3315 5873
rect 3263 5757 3315 5809
rect 3263 5693 3315 5745
rect 3263 5629 3315 5681
rect 3263 5565 3315 5617
rect 3263 5501 3315 5553
rect 3263 5437 3315 5489
rect 3263 5373 3315 5425
rect 3263 5309 3315 5361
rect 3263 5245 3315 5297
rect 3263 5181 3315 5233
rect 3263 5117 3315 5169
rect 3263 5053 3315 5105
rect 3263 4989 3315 5041
rect 3263 4925 3315 4977
rect 3263 4861 3315 4913
rect 3263 4797 3315 4849
rect -735 4326 -683 4347
rect -735 4295 -726 4326
rect -726 4295 -692 4326
rect -692 4295 -683 4326
rect -735 4254 -683 4283
rect -735 4231 -726 4254
rect -726 4231 -692 4254
rect -692 4231 -683 4254
rect -735 4182 -683 4219
rect -735 4167 -726 4182
rect -726 4167 -692 4182
rect -692 4167 -683 4182
rect -735 4148 -726 4155
rect -726 4148 -692 4155
rect -692 4148 -683 4155
rect -735 4110 -683 4148
rect -735 4103 -726 4110
rect -726 4103 -692 4110
rect -692 4103 -683 4110
rect -735 4076 -726 4091
rect -726 4076 -692 4091
rect -692 4076 -683 4091
rect -735 4039 -683 4076
rect -735 4004 -726 4027
rect -726 4004 -692 4027
rect -692 4004 -683 4027
rect -735 3975 -683 4004
rect -735 3932 -726 3963
rect -726 3932 -692 3963
rect -692 3932 -683 3963
rect -735 3911 -683 3932
rect -735 3894 -683 3899
rect -735 3860 -726 3894
rect -726 3860 -692 3894
rect -692 3860 -683 3894
rect -735 3847 -683 3860
rect -735 3822 -683 3835
rect -735 3788 -726 3822
rect -726 3788 -692 3822
rect -692 3788 -683 3822
rect -735 3783 -683 3788
rect -735 3750 -683 3771
rect -735 3719 -726 3750
rect -726 3719 -692 3750
rect -692 3719 -683 3750
rect -735 3678 -683 3707
rect -735 3655 -726 3678
rect -726 3655 -692 3678
rect -692 3655 -683 3678
rect -735 3606 -683 3643
rect -735 3591 -726 3606
rect -726 3591 -692 3606
rect -692 3591 -683 3606
rect -735 3572 -726 3579
rect -726 3572 -692 3579
rect -692 3572 -683 3579
rect -735 3534 -683 3572
rect -735 3527 -726 3534
rect -726 3527 -692 3534
rect -692 3527 -683 3534
rect -735 3500 -726 3515
rect -726 3500 -692 3515
rect -692 3500 -683 3515
rect -735 3463 -683 3500
rect -735 3428 -726 3451
rect -726 3428 -692 3451
rect -692 3428 -683 3451
rect -735 3399 -683 3428
rect -735 3356 -726 3387
rect -726 3356 -692 3387
rect -692 3356 -683 3387
rect -735 3335 -683 3356
rect -735 3318 -683 3323
rect -735 3284 -726 3318
rect -726 3284 -692 3318
rect -692 3284 -683 3318
rect -735 3271 -683 3284
rect -735 3246 -683 3259
rect -735 3212 -726 3246
rect -726 3212 -692 3246
rect -692 3212 -683 3246
rect -735 3207 -683 3212
rect -735 3174 -683 3195
rect -735 3143 -726 3174
rect -726 3143 -692 3174
rect -692 3143 -683 3174
rect -735 3102 -683 3131
rect -735 3079 -726 3102
rect -726 3079 -692 3102
rect -692 3079 -683 3102
rect -735 3030 -683 3067
rect -735 3015 -726 3030
rect -726 3015 -692 3030
rect -692 3015 -683 3030
rect -735 2996 -726 3003
rect -726 2996 -692 3003
rect -692 2996 -683 3003
rect -735 2958 -683 2996
rect -735 2951 -726 2958
rect -726 2951 -692 2958
rect -692 2951 -683 2958
rect -735 2924 -726 2939
rect -726 2924 -692 2939
rect -692 2924 -683 2939
rect -735 2887 -683 2924
rect -735 2852 -726 2875
rect -726 2852 -692 2875
rect -692 2852 -683 2875
rect -735 2823 -683 2852
rect -735 2780 -726 2811
rect -726 2780 -692 2811
rect -692 2780 -683 2811
rect -735 2759 -683 2780
rect 181 4326 233 4347
rect 181 4295 190 4326
rect 190 4295 224 4326
rect 224 4295 233 4326
rect 181 4254 233 4283
rect 181 4231 190 4254
rect 190 4231 224 4254
rect 224 4231 233 4254
rect 181 4182 233 4219
rect 181 4167 190 4182
rect 190 4167 224 4182
rect 224 4167 233 4182
rect 181 4148 190 4155
rect 190 4148 224 4155
rect 224 4148 233 4155
rect 181 4110 233 4148
rect 181 4103 190 4110
rect 190 4103 224 4110
rect 224 4103 233 4110
rect 181 4076 190 4091
rect 190 4076 224 4091
rect 224 4076 233 4091
rect 181 4039 233 4076
rect 181 4004 190 4027
rect 190 4004 224 4027
rect 224 4004 233 4027
rect 181 3975 233 4004
rect 181 3932 190 3963
rect 190 3932 224 3963
rect 224 3932 233 3963
rect 181 3911 233 3932
rect 181 3894 233 3899
rect 181 3860 190 3894
rect 190 3860 224 3894
rect 224 3860 233 3894
rect 181 3847 233 3860
rect 181 3822 233 3835
rect 181 3788 190 3822
rect 190 3788 224 3822
rect 224 3788 233 3822
rect 181 3783 233 3788
rect 181 3750 233 3771
rect 181 3719 190 3750
rect 190 3719 224 3750
rect 224 3719 233 3750
rect 181 3678 233 3707
rect 181 3655 190 3678
rect 190 3655 224 3678
rect 224 3655 233 3678
rect 181 3606 233 3643
rect 181 3591 190 3606
rect 190 3591 224 3606
rect 224 3591 233 3606
rect 181 3572 190 3579
rect 190 3572 224 3579
rect 224 3572 233 3579
rect 181 3534 233 3572
rect 181 3527 190 3534
rect 190 3527 224 3534
rect 224 3527 233 3534
rect 181 3500 190 3515
rect 190 3500 224 3515
rect 224 3500 233 3515
rect 181 3463 233 3500
rect 181 3428 190 3451
rect 190 3428 224 3451
rect 224 3428 233 3451
rect 181 3399 233 3428
rect 181 3356 190 3387
rect 190 3356 224 3387
rect 224 3356 233 3387
rect 181 3335 233 3356
rect 181 3318 233 3323
rect 181 3284 190 3318
rect 190 3284 224 3318
rect 224 3284 233 3318
rect 181 3271 233 3284
rect 181 3246 233 3259
rect 181 3212 190 3246
rect 190 3212 224 3246
rect 224 3212 233 3246
rect 181 3207 233 3212
rect 181 3174 233 3195
rect 181 3143 190 3174
rect 190 3143 224 3174
rect 224 3143 233 3174
rect 181 3102 233 3131
rect 181 3079 190 3102
rect 190 3079 224 3102
rect 224 3079 233 3102
rect 181 3030 233 3067
rect 181 3015 190 3030
rect 190 3015 224 3030
rect 224 3015 233 3030
rect 181 2996 190 3003
rect 190 2996 224 3003
rect 224 2996 233 3003
rect 181 2958 233 2996
rect 181 2951 190 2958
rect 190 2951 224 2958
rect 224 2951 233 2958
rect 181 2924 190 2939
rect 190 2924 224 2939
rect 224 2924 233 2939
rect 181 2887 233 2924
rect 181 2852 190 2875
rect 190 2852 224 2875
rect 224 2852 233 2875
rect 181 2823 233 2852
rect 181 2780 190 2811
rect 190 2780 224 2811
rect 224 2780 233 2811
rect 181 2759 233 2780
rect 1097 4326 1149 4347
rect 1097 4295 1106 4326
rect 1106 4295 1140 4326
rect 1140 4295 1149 4326
rect 1097 4254 1149 4283
rect 1097 4231 1106 4254
rect 1106 4231 1140 4254
rect 1140 4231 1149 4254
rect 1097 4182 1149 4219
rect 1097 4167 1106 4182
rect 1106 4167 1140 4182
rect 1140 4167 1149 4182
rect 1097 4148 1106 4155
rect 1106 4148 1140 4155
rect 1140 4148 1149 4155
rect 1097 4110 1149 4148
rect 1097 4103 1106 4110
rect 1106 4103 1140 4110
rect 1140 4103 1149 4110
rect 1097 4076 1106 4091
rect 1106 4076 1140 4091
rect 1140 4076 1149 4091
rect 1097 4039 1149 4076
rect 1097 4004 1106 4027
rect 1106 4004 1140 4027
rect 1140 4004 1149 4027
rect 1097 3975 1149 4004
rect 1097 3932 1106 3963
rect 1106 3932 1140 3963
rect 1140 3932 1149 3963
rect 1097 3911 1149 3932
rect 1097 3894 1149 3899
rect 1097 3860 1106 3894
rect 1106 3860 1140 3894
rect 1140 3860 1149 3894
rect 1097 3847 1149 3860
rect 1097 3822 1149 3835
rect 1097 3788 1106 3822
rect 1106 3788 1140 3822
rect 1140 3788 1149 3822
rect 1097 3783 1149 3788
rect 1097 3750 1149 3771
rect 1097 3719 1106 3750
rect 1106 3719 1140 3750
rect 1140 3719 1149 3750
rect 1097 3678 1149 3707
rect 1097 3655 1106 3678
rect 1106 3655 1140 3678
rect 1140 3655 1149 3678
rect 1097 3606 1149 3643
rect 1097 3591 1106 3606
rect 1106 3591 1140 3606
rect 1140 3591 1149 3606
rect 1097 3572 1106 3579
rect 1106 3572 1140 3579
rect 1140 3572 1149 3579
rect 1097 3534 1149 3572
rect 1097 3527 1106 3534
rect 1106 3527 1140 3534
rect 1140 3527 1149 3534
rect 1097 3500 1106 3515
rect 1106 3500 1140 3515
rect 1140 3500 1149 3515
rect 1097 3463 1149 3500
rect 1097 3428 1106 3451
rect 1106 3428 1140 3451
rect 1140 3428 1149 3451
rect 1097 3399 1149 3428
rect 1097 3356 1106 3387
rect 1106 3356 1140 3387
rect 1140 3356 1149 3387
rect 1097 3335 1149 3356
rect 1097 3318 1149 3323
rect 1097 3284 1106 3318
rect 1106 3284 1140 3318
rect 1140 3284 1149 3318
rect 1097 3271 1149 3284
rect 1097 3246 1149 3259
rect 1097 3212 1106 3246
rect 1106 3212 1140 3246
rect 1140 3212 1149 3246
rect 1097 3207 1149 3212
rect 1097 3174 1149 3195
rect 1097 3143 1106 3174
rect 1106 3143 1140 3174
rect 1140 3143 1149 3174
rect 1097 3102 1149 3131
rect 1097 3079 1106 3102
rect 1106 3079 1140 3102
rect 1140 3079 1149 3102
rect 1097 3030 1149 3067
rect 1097 3015 1106 3030
rect 1106 3015 1140 3030
rect 1140 3015 1149 3030
rect 1097 2996 1106 3003
rect 1106 2996 1140 3003
rect 1140 2996 1149 3003
rect 1097 2958 1149 2996
rect 1097 2951 1106 2958
rect 1106 2951 1140 2958
rect 1140 2951 1149 2958
rect 1097 2924 1106 2939
rect 1106 2924 1140 2939
rect 1140 2924 1149 2939
rect 1097 2887 1149 2924
rect 1097 2852 1106 2875
rect 1106 2852 1140 2875
rect 1140 2852 1149 2875
rect 1097 2823 1149 2852
rect 1097 2780 1106 2811
rect 1106 2780 1140 2811
rect 1140 2780 1149 2811
rect 1097 2759 1149 2780
rect 1431 4295 1483 4347
rect 1431 4231 1483 4283
rect 1431 4167 1483 4219
rect 1431 4103 1483 4155
rect 1431 4039 1483 4091
rect 1431 3975 1483 4027
rect 1431 3911 1483 3963
rect 1431 3847 1483 3899
rect 1431 3783 1483 3835
rect 1431 3719 1483 3771
rect 1431 3655 1483 3707
rect 1431 3591 1483 3643
rect 1431 3527 1483 3579
rect 1431 3463 1483 3515
rect 1431 3399 1483 3451
rect 1431 3335 1483 3387
rect 1431 3271 1483 3323
rect 1431 3207 1483 3259
rect 1431 3143 1483 3195
rect 1431 3079 1483 3131
rect 1431 3015 1483 3067
rect 1431 2951 1483 3003
rect 1431 2887 1483 2939
rect 1431 2823 1483 2875
rect 1431 2759 1483 2811
rect 2347 4295 2399 4347
rect 2347 4231 2399 4283
rect 2347 4167 2399 4219
rect 2347 4103 2399 4155
rect 2347 4039 2399 4091
rect 2347 3975 2399 4027
rect 2347 3911 2399 3963
rect 2347 3847 2399 3899
rect 2347 3783 2399 3835
rect 2347 3719 2399 3771
rect 2347 3655 2399 3707
rect 2347 3591 2399 3643
rect 2347 3527 2399 3579
rect 2347 3463 2399 3515
rect 2347 3399 2399 3451
rect 2347 3335 2399 3387
rect 2347 3271 2399 3323
rect 2347 3207 2399 3259
rect 2347 3143 2399 3195
rect 2347 3079 2399 3131
rect 2347 3015 2399 3067
rect 2347 2951 2399 3003
rect 2347 2887 2399 2939
rect 2347 2823 2399 2875
rect 2347 2759 2399 2811
rect 3263 4295 3315 4347
rect 3263 4231 3315 4283
rect 3263 4167 3315 4219
rect 3263 4103 3315 4155
rect 3263 4039 3315 4091
rect 3263 3975 3315 4027
rect 3263 3911 3315 3963
rect 3263 3847 3315 3899
rect 3263 3783 3315 3835
rect 3263 3719 3315 3771
rect 3263 3655 3315 3707
rect 3263 3591 3315 3643
rect 3263 3527 3315 3579
rect 3263 3463 3315 3515
rect 3263 3399 3315 3451
rect 3263 3335 3315 3387
rect 3263 3271 3315 3323
rect 3263 3207 3315 3259
rect 3263 3143 3315 3195
rect 3263 3079 3315 3131
rect 3263 3015 3315 3067
rect 3263 2951 3315 3003
rect 3263 2887 3315 2939
rect 3263 2823 3315 2875
rect 3263 2759 3315 2811
rect 851 2706 903 2712
rect 851 2672 860 2706
rect 860 2672 894 2706
rect 894 2672 903 2706
rect 851 2660 903 2672
rect 1653 2706 1705 2712
rect 1653 2672 1655 2706
rect 1655 2672 1689 2706
rect 1689 2672 1705 2706
rect 1653 2660 1705 2672
rect 207 2035 643 2407
rect 833 2031 885 2083
rect 1633 2041 2069 2413
rect 1401 1979 1453 2031
rect 106 1526 116 1559
rect 116 1526 150 1559
rect 150 1526 158 1559
rect 106 1507 158 1526
rect 713 1191 765 1243
rect 1555 1181 1607 1233
rect 717 1047 769 1099
rect 1553 1051 1605 1103
rect 102 738 154 757
rect 102 705 114 738
rect 114 705 148 738
rect 148 705 154 738
rect 2470 830 2522 882
rect 2618 1382 2670 1434
rect 1045 245 1097 297
rect 1213 247 1265 299
rect -1152 -615 -1100 -563
rect -1152 -679 -1100 -627
rect -1152 -743 -1100 -691
rect -1152 -807 -1100 -755
rect -1152 -871 -1100 -819
rect -1152 -935 -1100 -883
rect -1152 -999 -1100 -947
rect -1152 -1063 -1100 -1011
rect -1152 -1127 -1100 -1075
rect -1152 -1191 -1100 -1139
rect -1152 -1255 -1100 -1203
rect -1152 -1319 -1100 -1267
rect -1152 -1383 -1100 -1331
rect -1152 -1447 -1100 -1395
rect -1152 -1511 -1100 -1459
rect -1152 -1575 -1100 -1523
rect -1152 -1639 -1100 -1587
rect -1152 -1703 -1100 -1651
rect -1152 -1767 -1100 -1715
rect -1152 -1831 -1100 -1779
rect -1152 -1895 -1100 -1843
rect -1152 -1959 -1100 -1907
rect -1152 -2023 -1100 -1971
rect -1152 -2087 -1100 -2035
rect -1152 -2151 -1100 -2099
rect -1152 -2215 -1100 -2163
rect -1152 -2279 -1100 -2227
rect -1152 -2343 -1100 -2291
rect -1152 -2407 -1100 -2355
rect -1152 -2471 -1100 -2419
rect -1152 -2535 -1100 -2483
rect -1152 -2599 -1100 -2547
rect -1152 -2663 -1100 -2611
rect -1152 -2727 -1100 -2675
rect -1152 -2791 -1100 -2739
rect -1152 -2855 -1100 -2803
rect -1152 -2919 -1100 -2867
rect -1152 -2983 -1100 -2931
rect -1152 -3047 -1100 -2995
rect -1152 -3111 -1100 -3059
rect -1152 -3175 -1100 -3123
rect -694 -615 -642 -563
rect -694 -679 -642 -627
rect -694 -743 -642 -691
rect -694 -807 -642 -755
rect -694 -871 -642 -819
rect -694 -935 -642 -883
rect -694 -999 -642 -947
rect -694 -1063 -642 -1011
rect -694 -1127 -642 -1075
rect -694 -1191 -642 -1139
rect -694 -1255 -642 -1203
rect -694 -1319 -642 -1267
rect -694 -1383 -642 -1331
rect -694 -1447 -642 -1395
rect -694 -1511 -642 -1459
rect -694 -1575 -642 -1523
rect -694 -1639 -642 -1587
rect -694 -1703 -642 -1651
rect -694 -1767 -642 -1715
rect -694 -1831 -642 -1779
rect -694 -1895 -642 -1843
rect -694 -1959 -642 -1907
rect -694 -2023 -642 -1971
rect -694 -2087 -642 -2035
rect -694 -2151 -642 -2099
rect -694 -2215 -642 -2163
rect -694 -2279 -642 -2227
rect -694 -2343 -642 -2291
rect -694 -2407 -642 -2355
rect -694 -2471 -642 -2419
rect -694 -2535 -642 -2483
rect -694 -2599 -642 -2547
rect -694 -2663 -642 -2611
rect -694 -2727 -642 -2675
rect -694 -2791 -642 -2739
rect -694 -2855 -642 -2803
rect -694 -2919 -642 -2867
rect -694 -2983 -642 -2931
rect -694 -3047 -642 -2995
rect -694 -3111 -642 -3059
rect -694 -3175 -642 -3123
rect -236 -615 -184 -563
rect -236 -679 -184 -627
rect -236 -743 -184 -691
rect -236 -807 -184 -755
rect -236 -871 -184 -819
rect -236 -935 -184 -883
rect -236 -999 -184 -947
rect -236 -1063 -184 -1011
rect -236 -1127 -184 -1075
rect -236 -1191 -184 -1139
rect -236 -1255 -184 -1203
rect -236 -1319 -184 -1267
rect -236 -1383 -184 -1331
rect -236 -1447 -184 -1395
rect -236 -1511 -184 -1459
rect -236 -1575 -184 -1523
rect -236 -1639 -184 -1587
rect -236 -1703 -184 -1651
rect -236 -1767 -184 -1715
rect -236 -1831 -184 -1779
rect -236 -1895 -184 -1843
rect -236 -1959 -184 -1907
rect -236 -2023 -184 -1971
rect -236 -2087 -184 -2035
rect -236 -2151 -184 -2099
rect -236 -2215 -184 -2163
rect -236 -2279 -184 -2227
rect -236 -2343 -184 -2291
rect -236 -2407 -184 -2355
rect -236 -2471 -184 -2419
rect -236 -2535 -184 -2483
rect -236 -2599 -184 -2547
rect -236 -2663 -184 -2611
rect -236 -2727 -184 -2675
rect -236 -2791 -184 -2739
rect -236 -2855 -184 -2803
rect -236 -2919 -184 -2867
rect -236 -2983 -184 -2931
rect -236 -3047 -184 -2995
rect -236 -3111 -184 -3059
rect -236 -3175 -184 -3123
rect 222 -615 274 -563
rect 222 -679 274 -627
rect 222 -743 274 -691
rect 222 -807 274 -755
rect 222 -871 274 -819
rect 222 -935 274 -883
rect 222 -999 274 -947
rect 222 -1063 274 -1011
rect 222 -1127 274 -1075
rect 222 -1191 274 -1139
rect 222 -1255 274 -1203
rect 222 -1319 274 -1267
rect 222 -1383 274 -1331
rect 222 -1447 274 -1395
rect 222 -1511 274 -1459
rect 222 -1575 274 -1523
rect 222 -1639 274 -1587
rect 222 -1703 274 -1651
rect 222 -1767 274 -1715
rect 222 -1831 274 -1779
rect 222 -1895 274 -1843
rect 222 -1959 274 -1907
rect 222 -2023 274 -1971
rect 222 -2087 274 -2035
rect 222 -2151 274 -2099
rect 222 -2215 274 -2163
rect 222 -2279 274 -2227
rect 222 -2343 274 -2291
rect 222 -2407 274 -2355
rect 222 -2471 274 -2419
rect 222 -2535 274 -2483
rect 222 -2599 274 -2547
rect 222 -2663 274 -2611
rect 222 -2727 274 -2675
rect 222 -2791 274 -2739
rect 222 -2855 274 -2803
rect 222 -2919 274 -2867
rect 222 -2983 274 -2931
rect 222 -3047 274 -2995
rect 222 -3111 274 -3059
rect 222 -3175 274 -3123
rect 680 -615 732 -563
rect 680 -679 732 -627
rect 680 -743 732 -691
rect 680 -807 732 -755
rect 680 -871 732 -819
rect 680 -935 732 -883
rect 680 -999 732 -947
rect 680 -1063 732 -1011
rect 680 -1127 732 -1075
rect 680 -1191 732 -1139
rect 680 -1255 732 -1203
rect 680 -1319 732 -1267
rect 680 -1383 732 -1331
rect 680 -1447 732 -1395
rect 680 -1511 732 -1459
rect 680 -1575 732 -1523
rect 680 -1639 732 -1587
rect 680 -1703 732 -1651
rect 680 -1767 732 -1715
rect 680 -1831 732 -1779
rect 680 -1895 732 -1843
rect 680 -1959 732 -1907
rect 680 -2023 732 -1971
rect 680 -2087 732 -2035
rect 680 -2151 732 -2099
rect 680 -2215 732 -2163
rect 680 -2279 732 -2227
rect 680 -2343 732 -2291
rect 680 -2407 732 -2355
rect 680 -2471 732 -2419
rect 680 -2535 732 -2483
rect 680 -2599 732 -2547
rect 680 -2663 732 -2611
rect 680 -2727 732 -2675
rect 680 -2791 732 -2739
rect 680 -2855 732 -2803
rect 680 -2919 732 -2867
rect 680 -2983 732 -2931
rect 680 -3047 732 -2995
rect 680 -3111 732 -3059
rect 680 -3175 732 -3123
rect 1138 -615 1190 -563
rect 1138 -679 1190 -627
rect 1138 -743 1190 -691
rect 1138 -807 1190 -755
rect 1138 -871 1190 -819
rect 1138 -935 1190 -883
rect 1138 -999 1190 -947
rect 1138 -1063 1190 -1011
rect 1138 -1127 1190 -1075
rect 1138 -1191 1190 -1139
rect 1138 -1255 1190 -1203
rect 1138 -1319 1190 -1267
rect 1138 -1383 1190 -1331
rect 1138 -1447 1190 -1395
rect 1138 -1511 1190 -1459
rect 1138 -1575 1190 -1523
rect 1138 -1639 1190 -1587
rect 1138 -1703 1190 -1651
rect 1138 -1767 1190 -1715
rect 1138 -1831 1190 -1779
rect 1138 -1895 1190 -1843
rect 1138 -1959 1190 -1907
rect 1138 -2023 1190 -1971
rect 1138 -2087 1190 -2035
rect 1138 -2151 1190 -2099
rect 1138 -2215 1190 -2163
rect 1138 -2279 1190 -2227
rect 1138 -2343 1190 -2291
rect 1138 -2407 1190 -2355
rect 1138 -2471 1190 -2419
rect 1138 -2535 1190 -2483
rect 1138 -2599 1190 -2547
rect 1138 -2663 1190 -2611
rect 1138 -2727 1190 -2675
rect 1138 -2791 1190 -2739
rect 1138 -2855 1190 -2803
rect 1138 -2919 1190 -2867
rect 1138 -2983 1190 -2931
rect 1138 -3047 1190 -2995
rect 1138 -3111 1190 -3059
rect 1138 -3175 1190 -3123
rect 1596 -615 1648 -563
rect 1596 -679 1648 -627
rect 1596 -743 1648 -691
rect 1596 -807 1648 -755
rect 1596 -871 1648 -819
rect 1596 -935 1648 -883
rect 1596 -999 1648 -947
rect 1596 -1063 1648 -1011
rect 1596 -1127 1648 -1075
rect 1596 -1191 1648 -1139
rect 1596 -1255 1648 -1203
rect 1596 -1319 1648 -1267
rect 1596 -1383 1648 -1331
rect 1596 -1447 1648 -1395
rect 1596 -1511 1648 -1459
rect 1596 -1575 1648 -1523
rect 1596 -1639 1648 -1587
rect 1596 -1703 1648 -1651
rect 1596 -1767 1648 -1715
rect 1596 -1831 1648 -1779
rect 1596 -1895 1648 -1843
rect 1596 -1959 1648 -1907
rect 1596 -2023 1648 -1971
rect 1596 -2087 1648 -2035
rect 1596 -2151 1648 -2099
rect 1596 -2215 1648 -2163
rect 1596 -2279 1648 -2227
rect 1596 -2343 1648 -2291
rect 1596 -2407 1648 -2355
rect 1596 -2471 1648 -2419
rect 1596 -2535 1648 -2483
rect 1596 -2599 1648 -2547
rect 1596 -2663 1648 -2611
rect 1596 -2727 1648 -2675
rect 1596 -2791 1648 -2739
rect 1596 -2855 1648 -2803
rect 1596 -2919 1648 -2867
rect 1596 -2983 1648 -2931
rect 1596 -3047 1648 -2995
rect 1596 -3111 1648 -3059
rect 1596 -3175 1648 -3123
rect 2054 -615 2106 -563
rect 2054 -679 2106 -627
rect 2054 -743 2106 -691
rect 2054 -807 2106 -755
rect 2054 -871 2106 -819
rect 2054 -935 2106 -883
rect 2054 -999 2106 -947
rect 2054 -1063 2106 -1011
rect 2054 -1127 2106 -1075
rect 2054 -1191 2106 -1139
rect 2054 -1255 2106 -1203
rect 2054 -1319 2106 -1267
rect 2054 -1383 2106 -1331
rect 2054 -1447 2106 -1395
rect 2054 -1511 2106 -1459
rect 2054 -1575 2106 -1523
rect 2054 -1639 2106 -1587
rect 2054 -1703 2106 -1651
rect 2054 -1767 2106 -1715
rect 2054 -1831 2106 -1779
rect 2054 -1895 2106 -1843
rect 2054 -1959 2106 -1907
rect 2054 -2023 2106 -1971
rect 2054 -2087 2106 -2035
rect 2054 -2151 2106 -2099
rect 2054 -2215 2106 -2163
rect 2054 -2279 2106 -2227
rect 2054 -2343 2106 -2291
rect 2054 -2407 2106 -2355
rect 2054 -2471 2106 -2419
rect 2054 -2535 2106 -2483
rect 2054 -2599 2106 -2547
rect 2054 -2663 2106 -2611
rect 2054 -2727 2106 -2675
rect 2054 -2791 2106 -2739
rect 2054 -2855 2106 -2803
rect 2054 -2919 2106 -2867
rect 2054 -2983 2106 -2931
rect 2054 -3047 2106 -2995
rect 2054 -3111 2106 -3059
rect 2054 -3175 2106 -3123
rect 2512 -615 2564 -563
rect 2512 -679 2564 -627
rect 2512 -743 2564 -691
rect 2512 -807 2564 -755
rect 2512 -871 2564 -819
rect 2512 -935 2564 -883
rect 2512 -999 2564 -947
rect 2512 -1063 2564 -1011
rect 2512 -1127 2564 -1075
rect 2512 -1191 2564 -1139
rect 2512 -1255 2564 -1203
rect 2512 -1319 2564 -1267
rect 2512 -1383 2564 -1331
rect 2512 -1447 2564 -1395
rect 2512 -1511 2564 -1459
rect 2512 -1575 2564 -1523
rect 2512 -1639 2564 -1587
rect 2512 -1703 2564 -1651
rect 2512 -1767 2564 -1715
rect 2512 -1831 2564 -1779
rect 2512 -1895 2564 -1843
rect 2512 -1959 2564 -1907
rect 2512 -2023 2564 -1971
rect 2512 -2087 2564 -2035
rect 2512 -2151 2564 -2099
rect 2512 -2215 2564 -2163
rect 2512 -2279 2564 -2227
rect 2512 -2343 2564 -2291
rect 2512 -2407 2564 -2355
rect 2512 -2471 2564 -2419
rect 2512 -2535 2564 -2483
rect 2512 -2599 2564 -2547
rect 2512 -2663 2564 -2611
rect 2512 -2727 2564 -2675
rect 2512 -2791 2564 -2739
rect 2512 -2855 2564 -2803
rect 2512 -2919 2564 -2867
rect 2512 -2983 2564 -2931
rect 2512 -3047 2564 -2995
rect 2512 -3111 2564 -3059
rect 2512 -3175 2564 -3123
rect 2970 -615 3022 -563
rect 2970 -679 3022 -627
rect 2970 -743 3022 -691
rect 2970 -807 3022 -755
rect 2970 -871 3022 -819
rect 2970 -935 3022 -883
rect 2970 -999 3022 -947
rect 2970 -1063 3022 -1011
rect 2970 -1127 3022 -1075
rect 2970 -1191 3022 -1139
rect 2970 -1255 3022 -1203
rect 2970 -1319 3022 -1267
rect 2970 -1383 3022 -1331
rect 2970 -1447 3022 -1395
rect 2970 -1511 3022 -1459
rect 2970 -1575 3022 -1523
rect 2970 -1639 3022 -1587
rect 2970 -1703 3022 -1651
rect 2970 -1767 3022 -1715
rect 2970 -1831 3022 -1779
rect 2970 -1895 3022 -1843
rect 2970 -1959 3022 -1907
rect 2970 -2023 3022 -1971
rect 2970 -2087 3022 -2035
rect 2970 -2151 3022 -2099
rect 2970 -2215 3022 -2163
rect 2970 -2279 3022 -2227
rect 2970 -2343 3022 -2291
rect 2970 -2407 3022 -2355
rect 2970 -2471 3022 -2419
rect 2970 -2535 3022 -2483
rect 2970 -2599 3022 -2547
rect 2970 -2663 3022 -2611
rect 2970 -2727 3022 -2675
rect 2970 -2791 3022 -2739
rect 2970 -2855 3022 -2803
rect 2970 -2919 3022 -2867
rect 2970 -2983 3022 -2931
rect 2970 -3047 3022 -2995
rect 2970 -3111 3022 -3059
rect 2970 -3175 3022 -3123
rect 3428 -615 3480 -563
rect 3428 -679 3480 -627
rect 3428 -743 3480 -691
rect 3428 -807 3480 -755
rect 3428 -871 3480 -819
rect 3428 -935 3480 -883
rect 3428 -999 3480 -947
rect 3428 -1063 3480 -1011
rect 3428 -1127 3480 -1075
rect 3428 -1191 3480 -1139
rect 3428 -1255 3480 -1203
rect 3428 -1319 3480 -1267
rect 3428 -1383 3480 -1331
rect 3428 -1447 3480 -1395
rect 3428 -1511 3480 -1459
rect 3428 -1575 3480 -1523
rect 3428 -1639 3480 -1587
rect 3428 -1703 3480 -1651
rect 3428 -1767 3480 -1715
rect 3428 -1831 3480 -1779
rect 3428 -1895 3480 -1843
rect 3428 -1959 3480 -1907
rect 3428 -2023 3480 -1971
rect 3428 -2087 3480 -2035
rect 3428 -2151 3480 -2099
rect 3428 -2215 3480 -2163
rect 3428 -2279 3480 -2227
rect 3428 -2343 3480 -2291
rect 3428 -2407 3480 -2355
rect 3428 -2471 3480 -2419
rect 3428 -2535 3480 -2483
rect 3428 -2599 3480 -2547
rect 3428 -2663 3480 -2611
rect 3428 -2727 3480 -2675
rect 3428 -2791 3480 -2739
rect 3428 -2855 3480 -2803
rect 3428 -2919 3480 -2867
rect 3428 -2983 3480 -2931
rect 3428 -3047 3480 -2995
rect 3428 -3111 3480 -3059
rect 3428 -3175 3480 -3123
<< metal2 >>
rect -1202 6605 3782 6620
rect -1202 6553 -1200 6605
rect -1148 6553 -1136 6605
rect -1084 6553 -1072 6605
rect -1020 6553 -1008 6605
rect -956 6553 -944 6605
rect -892 6553 -880 6605
rect -828 6553 -816 6605
rect -764 6553 -752 6605
rect -700 6553 -688 6605
rect -636 6553 -624 6605
rect -572 6553 -560 6605
rect -508 6553 -496 6605
rect -444 6553 -432 6605
rect -380 6553 -368 6605
rect -316 6553 -304 6605
rect -252 6553 -240 6605
rect -188 6553 -176 6605
rect -124 6553 -112 6605
rect -60 6553 -48 6605
rect 4 6553 16 6605
rect 68 6553 80 6605
rect 132 6553 144 6605
rect 196 6553 208 6605
rect 260 6553 272 6605
rect 324 6553 336 6605
rect 388 6553 400 6605
rect 452 6553 464 6605
rect 516 6553 528 6605
rect 580 6553 592 6605
rect 644 6553 656 6605
rect 708 6553 720 6605
rect 772 6553 784 6605
rect 836 6553 848 6605
rect 900 6553 912 6605
rect 964 6553 976 6605
rect 1028 6553 1040 6605
rect 1092 6553 1104 6605
rect 1156 6553 1168 6605
rect 1220 6553 1232 6605
rect 1284 6553 1296 6605
rect 1348 6553 1360 6605
rect 1412 6553 1424 6605
rect 1476 6553 1488 6605
rect 1540 6553 1552 6605
rect 1604 6553 1616 6605
rect 1668 6553 1680 6605
rect 1732 6553 1744 6605
rect 1796 6553 1808 6605
rect 1860 6553 1872 6605
rect 1924 6553 1936 6605
rect 1988 6553 2000 6605
rect 2052 6553 2064 6605
rect 2116 6553 2128 6605
rect 2180 6553 2192 6605
rect 2244 6553 2256 6605
rect 2308 6553 2320 6605
rect 2372 6553 2384 6605
rect 2436 6553 2448 6605
rect 2500 6553 2512 6605
rect 2564 6553 2576 6605
rect 2628 6553 2640 6605
rect 2692 6553 2704 6605
rect 2756 6553 2768 6605
rect 2820 6553 2832 6605
rect 2884 6553 2896 6605
rect 2948 6553 2960 6605
rect 3012 6553 3024 6605
rect 3076 6553 3088 6605
rect 3140 6553 3152 6605
rect 3204 6553 3216 6605
rect 3268 6553 3280 6605
rect 3332 6553 3344 6605
rect 3396 6553 3408 6605
rect 3460 6553 3472 6605
rect 3524 6553 3536 6605
rect 3588 6553 3600 6605
rect 3652 6553 3664 6605
rect 3716 6553 3728 6605
rect 3780 6553 3782 6605
rect -1202 6538 3782 6553
rect -742 6385 -676 6398
rect -742 6333 -735 6385
rect -683 6333 -676 6385
rect -742 6321 -676 6333
rect -742 6269 -735 6321
rect -683 6269 -676 6321
rect -742 6257 -676 6269
rect -742 6205 -735 6257
rect -683 6205 -676 6257
rect -742 6193 -676 6205
rect -742 6141 -735 6193
rect -683 6141 -676 6193
rect -742 6129 -676 6141
rect -742 6077 -735 6129
rect -683 6077 -676 6129
rect -742 6065 -676 6077
rect -742 6013 -735 6065
rect -683 6013 -676 6065
rect -742 6001 -676 6013
rect -742 5949 -735 6001
rect -683 5949 -676 6001
rect -742 5937 -676 5949
rect -742 5885 -735 5937
rect -683 5885 -676 5937
rect -742 5873 -676 5885
rect -742 5821 -735 5873
rect -683 5821 -676 5873
rect -742 5809 -676 5821
rect -742 5757 -735 5809
rect -683 5757 -676 5809
rect -742 5745 -676 5757
rect -742 5693 -735 5745
rect -683 5693 -676 5745
rect -742 5681 -676 5693
rect -742 5629 -735 5681
rect -683 5629 -676 5681
rect -742 5617 -676 5629
rect -742 5565 -735 5617
rect -683 5565 -676 5617
rect -742 5553 -676 5565
rect -742 5501 -735 5553
rect -683 5501 -676 5553
rect -742 5489 -676 5501
rect -742 5437 -735 5489
rect -683 5437 -676 5489
rect -742 5425 -676 5437
rect -742 5373 -735 5425
rect -683 5373 -676 5425
rect -742 5361 -676 5373
rect -742 5309 -735 5361
rect -683 5309 -676 5361
rect -742 5297 -676 5309
rect -742 5245 -735 5297
rect -683 5245 -676 5297
rect -742 5233 -676 5245
rect -742 5181 -735 5233
rect -683 5181 -676 5233
rect -742 5169 -676 5181
rect -742 5117 -735 5169
rect -683 5117 -676 5169
rect -742 5105 -676 5117
rect -742 5053 -735 5105
rect -683 5053 -676 5105
rect -742 5041 -676 5053
rect -742 4989 -735 5041
rect -683 4989 -676 5041
rect -742 4977 -676 4989
rect -742 4925 -735 4977
rect -683 4925 -676 4977
rect -742 4913 -676 4925
rect -742 4861 -735 4913
rect -683 4861 -676 4913
rect -742 4849 -676 4861
rect -742 4797 -735 4849
rect -683 4797 -676 4849
rect -742 4347 -676 4797
rect -742 4295 -735 4347
rect -683 4295 -676 4347
rect -742 4283 -676 4295
rect -742 4231 -735 4283
rect -683 4231 -676 4283
rect -742 4219 -676 4231
rect -742 4167 -735 4219
rect -683 4167 -676 4219
rect -742 4155 -676 4167
rect -742 4103 -735 4155
rect -683 4103 -676 4155
rect -742 4091 -676 4103
rect -742 4039 -735 4091
rect -683 4039 -676 4091
rect -742 4027 -676 4039
rect -742 3975 -735 4027
rect -683 3975 -676 4027
rect -742 3963 -676 3975
rect -742 3911 -735 3963
rect -683 3911 -676 3963
rect -742 3899 -676 3911
rect -742 3847 -735 3899
rect -683 3847 -676 3899
rect -742 3835 -676 3847
rect -742 3783 -735 3835
rect -683 3783 -676 3835
rect -742 3771 -676 3783
rect -742 3719 -735 3771
rect -683 3719 -676 3771
rect -742 3707 -676 3719
rect -742 3655 -735 3707
rect -683 3655 -676 3707
rect -742 3643 -676 3655
rect -742 3591 -735 3643
rect -683 3591 -676 3643
rect -742 3579 -676 3591
rect -742 3527 -735 3579
rect -683 3527 -676 3579
rect -742 3515 -676 3527
rect -742 3463 -735 3515
rect -683 3463 -676 3515
rect -742 3451 -676 3463
rect -742 3399 -735 3451
rect -683 3399 -676 3451
rect -742 3387 -676 3399
rect -742 3335 -735 3387
rect -683 3335 -676 3387
rect -742 3323 -676 3335
rect -742 3271 -735 3323
rect -683 3271 -676 3323
rect -742 3259 -676 3271
rect -742 3207 -735 3259
rect -683 3207 -676 3259
rect -742 3195 -676 3207
rect -742 3143 -735 3195
rect -683 3143 -676 3195
rect -742 3131 -676 3143
rect -742 3079 -735 3131
rect -683 3079 -676 3131
rect -742 3067 -676 3079
rect -742 3015 -735 3067
rect -683 3015 -676 3067
rect -742 3003 -676 3015
rect -742 2951 -735 3003
rect -683 2951 -676 3003
rect -742 2939 -676 2951
rect -742 2887 -735 2939
rect -683 2887 -676 2939
rect -742 2875 -676 2887
rect -742 2823 -735 2875
rect -683 2823 -676 2875
rect -742 2811 -676 2823
rect -742 2759 -735 2811
rect -683 2759 -676 2811
rect -742 2474 -676 2759
rect 174 6385 240 6398
rect 174 6333 181 6385
rect 233 6333 240 6385
rect 174 6321 240 6333
rect 174 6269 181 6321
rect 233 6269 240 6321
rect 174 6257 240 6269
rect 174 6205 181 6257
rect 233 6205 240 6257
rect 174 6193 240 6205
rect 174 6141 181 6193
rect 233 6141 240 6193
rect 174 6129 240 6141
rect 174 6077 181 6129
rect 233 6077 240 6129
rect 174 6065 240 6077
rect 174 6013 181 6065
rect 233 6013 240 6065
rect 174 6001 240 6013
rect 174 5949 181 6001
rect 233 5949 240 6001
rect 174 5937 240 5949
rect 174 5885 181 5937
rect 233 5885 240 5937
rect 174 5873 240 5885
rect 174 5821 181 5873
rect 233 5821 240 5873
rect 174 5809 240 5821
rect 174 5757 181 5809
rect 233 5757 240 5809
rect 174 5745 240 5757
rect 174 5693 181 5745
rect 233 5693 240 5745
rect 174 5681 240 5693
rect 174 5629 181 5681
rect 233 5629 240 5681
rect 174 5617 240 5629
rect 174 5565 181 5617
rect 233 5565 240 5617
rect 174 5553 240 5565
rect 174 5501 181 5553
rect 233 5501 240 5553
rect 174 5489 240 5501
rect 174 5437 181 5489
rect 233 5437 240 5489
rect 174 5425 240 5437
rect 174 5373 181 5425
rect 233 5373 240 5425
rect 174 5361 240 5373
rect 174 5309 181 5361
rect 233 5309 240 5361
rect 174 5297 240 5309
rect 174 5245 181 5297
rect 233 5245 240 5297
rect 174 5233 240 5245
rect 174 5181 181 5233
rect 233 5181 240 5233
rect 174 5169 240 5181
rect 174 5117 181 5169
rect 233 5117 240 5169
rect 174 5105 240 5117
rect 174 5053 181 5105
rect 233 5053 240 5105
rect 174 5041 240 5053
rect 174 4989 181 5041
rect 233 4989 240 5041
rect 174 4977 240 4989
rect 174 4925 181 4977
rect 233 4925 240 4977
rect 174 4913 240 4925
rect 174 4861 181 4913
rect 233 4861 240 4913
rect 174 4849 240 4861
rect 174 4797 181 4849
rect 233 4797 240 4849
rect 174 4347 240 4797
rect 174 4295 181 4347
rect 233 4295 240 4347
rect 174 4283 240 4295
rect 174 4231 181 4283
rect 233 4231 240 4283
rect 174 4219 240 4231
rect 174 4167 181 4219
rect 233 4167 240 4219
rect 174 4155 240 4167
rect 174 4103 181 4155
rect 233 4103 240 4155
rect 174 4091 240 4103
rect 174 4039 181 4091
rect 233 4039 240 4091
rect 174 4027 240 4039
rect 174 3975 181 4027
rect 233 3975 240 4027
rect 174 3963 240 3975
rect 174 3911 181 3963
rect 233 3911 240 3963
rect 174 3899 240 3911
rect 174 3847 181 3899
rect 233 3847 240 3899
rect 174 3835 240 3847
rect 174 3783 181 3835
rect 233 3783 240 3835
rect 174 3771 240 3783
rect 174 3719 181 3771
rect 233 3719 240 3771
rect 174 3707 240 3719
rect 174 3655 181 3707
rect 233 3655 240 3707
rect 174 3643 240 3655
rect 174 3591 181 3643
rect 233 3591 240 3643
rect 174 3579 240 3591
rect 174 3527 181 3579
rect 233 3527 240 3579
rect 174 3515 240 3527
rect 174 3463 181 3515
rect 233 3463 240 3515
rect 174 3451 240 3463
rect 174 3399 181 3451
rect 233 3399 240 3451
rect 174 3387 240 3399
rect 174 3335 181 3387
rect 233 3335 240 3387
rect 174 3323 240 3335
rect 174 3271 181 3323
rect 233 3271 240 3323
rect 174 3259 240 3271
rect 174 3207 181 3259
rect 233 3207 240 3259
rect 174 3195 240 3207
rect 174 3143 181 3195
rect 233 3143 240 3195
rect 174 3131 240 3143
rect 174 3079 181 3131
rect 233 3079 240 3131
rect 174 3067 240 3079
rect 174 3015 181 3067
rect 233 3015 240 3067
rect 174 3003 240 3015
rect 174 2951 181 3003
rect 233 2951 240 3003
rect 174 2939 240 2951
rect 174 2887 181 2939
rect 233 2887 240 2939
rect 174 2875 240 2887
rect 174 2823 181 2875
rect 233 2823 240 2875
rect 174 2811 240 2823
rect 174 2759 181 2811
rect 233 2759 240 2811
rect 174 2474 240 2759
rect 1090 6385 1156 6398
rect 1090 6333 1097 6385
rect 1149 6333 1156 6385
rect 1090 6321 1156 6333
rect 1090 6269 1097 6321
rect 1149 6269 1156 6321
rect 1090 6257 1156 6269
rect 1090 6205 1097 6257
rect 1149 6205 1156 6257
rect 1090 6193 1156 6205
rect 1090 6141 1097 6193
rect 1149 6141 1156 6193
rect 1090 6129 1156 6141
rect 1090 6077 1097 6129
rect 1149 6077 1156 6129
rect 1090 6065 1156 6077
rect 1090 6013 1097 6065
rect 1149 6013 1156 6065
rect 1090 6001 1156 6013
rect 1090 5949 1097 6001
rect 1149 5949 1156 6001
rect 1090 5937 1156 5949
rect 1090 5885 1097 5937
rect 1149 5885 1156 5937
rect 1090 5873 1156 5885
rect 1090 5821 1097 5873
rect 1149 5821 1156 5873
rect 1090 5809 1156 5821
rect 1090 5757 1097 5809
rect 1149 5757 1156 5809
rect 1090 5745 1156 5757
rect 1090 5693 1097 5745
rect 1149 5693 1156 5745
rect 1090 5681 1156 5693
rect 1090 5629 1097 5681
rect 1149 5629 1156 5681
rect 1090 5617 1156 5629
rect 1090 5565 1097 5617
rect 1149 5565 1156 5617
rect 1090 5553 1156 5565
rect 1090 5501 1097 5553
rect 1149 5501 1156 5553
rect 1090 5489 1156 5501
rect 1090 5437 1097 5489
rect 1149 5437 1156 5489
rect 1090 5425 1156 5437
rect 1090 5373 1097 5425
rect 1149 5373 1156 5425
rect 1090 5361 1156 5373
rect 1090 5309 1097 5361
rect 1149 5309 1156 5361
rect 1090 5297 1156 5309
rect 1090 5245 1097 5297
rect 1149 5245 1156 5297
rect 1090 5233 1156 5245
rect 1090 5181 1097 5233
rect 1149 5181 1156 5233
rect 1090 5169 1156 5181
rect 1090 5117 1097 5169
rect 1149 5117 1156 5169
rect 1090 5105 1156 5117
rect 1090 5053 1097 5105
rect 1149 5053 1156 5105
rect 1090 5041 1156 5053
rect 1090 4989 1097 5041
rect 1149 4989 1156 5041
rect 1090 4977 1156 4989
rect 1090 4925 1097 4977
rect 1149 4925 1156 4977
rect 1090 4913 1156 4925
rect 1090 4861 1097 4913
rect 1149 4861 1156 4913
rect 1090 4849 1156 4861
rect 1090 4797 1097 4849
rect 1149 4797 1156 4849
rect 1090 4347 1156 4797
rect 1090 4295 1097 4347
rect 1149 4295 1156 4347
rect 1090 4283 1156 4295
rect 1090 4231 1097 4283
rect 1149 4231 1156 4283
rect 1090 4219 1156 4231
rect 1090 4167 1097 4219
rect 1149 4167 1156 4219
rect 1090 4155 1156 4167
rect 1090 4103 1097 4155
rect 1149 4103 1156 4155
rect 1090 4091 1156 4103
rect 1090 4039 1097 4091
rect 1149 4039 1156 4091
rect 1090 4027 1156 4039
rect 1090 3975 1097 4027
rect 1149 3975 1156 4027
rect 1090 3963 1156 3975
rect 1090 3911 1097 3963
rect 1149 3911 1156 3963
rect 1090 3899 1156 3911
rect 1090 3847 1097 3899
rect 1149 3847 1156 3899
rect 1090 3835 1156 3847
rect 1090 3783 1097 3835
rect 1149 3783 1156 3835
rect 1090 3771 1156 3783
rect 1090 3719 1097 3771
rect 1149 3719 1156 3771
rect 1090 3707 1156 3719
rect 1090 3655 1097 3707
rect 1149 3655 1156 3707
rect 1090 3643 1156 3655
rect 1090 3591 1097 3643
rect 1149 3591 1156 3643
rect 1090 3579 1156 3591
rect 1090 3527 1097 3579
rect 1149 3527 1156 3579
rect 1090 3515 1156 3527
rect 1090 3463 1097 3515
rect 1149 3463 1156 3515
rect 1090 3451 1156 3463
rect 1090 3399 1097 3451
rect 1149 3399 1156 3451
rect 1090 3387 1156 3399
rect 1090 3335 1097 3387
rect 1149 3335 1156 3387
rect 1090 3323 1156 3335
rect 1090 3271 1097 3323
rect 1149 3271 1156 3323
rect 1090 3259 1156 3271
rect 1090 3207 1097 3259
rect 1149 3207 1156 3259
rect 1090 3195 1156 3207
rect 1090 3143 1097 3195
rect 1149 3143 1156 3195
rect 1090 3131 1156 3143
rect 1090 3079 1097 3131
rect 1149 3079 1156 3131
rect 1090 3067 1156 3079
rect 1090 3015 1097 3067
rect 1149 3015 1156 3067
rect 1090 3003 1156 3015
rect 1090 2951 1097 3003
rect 1149 2951 1156 3003
rect 1090 2939 1156 2951
rect 1090 2887 1097 2939
rect 1149 2887 1156 2939
rect 1090 2875 1156 2887
rect 1090 2823 1097 2875
rect 1149 2823 1156 2875
rect 1090 2811 1156 2823
rect 1090 2759 1097 2811
rect 1149 2759 1156 2811
rect 836 2714 918 2732
rect 836 2658 849 2714
rect 905 2658 918 2714
rect 836 2640 918 2658
rect 1090 2474 1156 2759
rect -742 2407 1156 2474
rect -742 2396 207 2407
rect 188 2035 207 2396
rect 643 2396 1156 2407
rect 1424 6385 1490 6398
rect 1424 6333 1431 6385
rect 1483 6333 1490 6385
rect 1424 6321 1490 6333
rect 1424 6269 1431 6321
rect 1483 6269 1490 6321
rect 1424 6257 1490 6269
rect 1424 6205 1431 6257
rect 1483 6205 1490 6257
rect 1424 6193 1490 6205
rect 1424 6141 1431 6193
rect 1483 6141 1490 6193
rect 1424 6129 1490 6141
rect 1424 6077 1431 6129
rect 1483 6077 1490 6129
rect 1424 6065 1490 6077
rect 1424 6013 1431 6065
rect 1483 6013 1490 6065
rect 1424 6001 1490 6013
rect 1424 5949 1431 6001
rect 1483 5949 1490 6001
rect 1424 5937 1490 5949
rect 1424 5885 1431 5937
rect 1483 5885 1490 5937
rect 1424 5873 1490 5885
rect 1424 5821 1431 5873
rect 1483 5821 1490 5873
rect 1424 5809 1490 5821
rect 1424 5757 1431 5809
rect 1483 5757 1490 5809
rect 1424 5745 1490 5757
rect 1424 5693 1431 5745
rect 1483 5693 1490 5745
rect 1424 5681 1490 5693
rect 1424 5629 1431 5681
rect 1483 5629 1490 5681
rect 1424 5617 1490 5629
rect 1424 5565 1431 5617
rect 1483 5565 1490 5617
rect 1424 5553 1490 5565
rect 1424 5501 1431 5553
rect 1483 5501 1490 5553
rect 1424 5489 1490 5501
rect 1424 5437 1431 5489
rect 1483 5437 1490 5489
rect 1424 5425 1490 5437
rect 1424 5373 1431 5425
rect 1483 5373 1490 5425
rect 1424 5361 1490 5373
rect 1424 5309 1431 5361
rect 1483 5309 1490 5361
rect 1424 5297 1490 5309
rect 1424 5245 1431 5297
rect 1483 5245 1490 5297
rect 1424 5233 1490 5245
rect 1424 5181 1431 5233
rect 1483 5181 1490 5233
rect 1424 5169 1490 5181
rect 1424 5117 1431 5169
rect 1483 5117 1490 5169
rect 1424 5105 1490 5117
rect 1424 5053 1431 5105
rect 1483 5053 1490 5105
rect 1424 5041 1490 5053
rect 1424 4989 1431 5041
rect 1483 4989 1490 5041
rect 1424 4977 1490 4989
rect 1424 4925 1431 4977
rect 1483 4925 1490 4977
rect 1424 4913 1490 4925
rect 1424 4861 1431 4913
rect 1483 4861 1490 4913
rect 1424 4849 1490 4861
rect 1424 4797 1431 4849
rect 1483 4797 1490 4849
rect 1424 4347 1490 4797
rect 1424 4295 1431 4347
rect 1483 4295 1490 4347
rect 1424 4283 1490 4295
rect 1424 4231 1431 4283
rect 1483 4231 1490 4283
rect 1424 4219 1490 4231
rect 1424 4167 1431 4219
rect 1483 4167 1490 4219
rect 1424 4155 1490 4167
rect 1424 4103 1431 4155
rect 1483 4103 1490 4155
rect 1424 4091 1490 4103
rect 1424 4039 1431 4091
rect 1483 4039 1490 4091
rect 1424 4027 1490 4039
rect 1424 3975 1431 4027
rect 1483 3975 1490 4027
rect 1424 3963 1490 3975
rect 1424 3911 1431 3963
rect 1483 3911 1490 3963
rect 1424 3899 1490 3911
rect 1424 3847 1431 3899
rect 1483 3847 1490 3899
rect 1424 3835 1490 3847
rect 1424 3783 1431 3835
rect 1483 3783 1490 3835
rect 1424 3771 1490 3783
rect 1424 3719 1431 3771
rect 1483 3719 1490 3771
rect 1424 3707 1490 3719
rect 1424 3655 1431 3707
rect 1483 3655 1490 3707
rect 1424 3643 1490 3655
rect 1424 3591 1431 3643
rect 1483 3591 1490 3643
rect 1424 3579 1490 3591
rect 1424 3527 1431 3579
rect 1483 3527 1490 3579
rect 1424 3515 1490 3527
rect 1424 3463 1431 3515
rect 1483 3463 1490 3515
rect 1424 3451 1490 3463
rect 1424 3399 1431 3451
rect 1483 3399 1490 3451
rect 1424 3387 1490 3399
rect 1424 3335 1431 3387
rect 1483 3335 1490 3387
rect 1424 3323 1490 3335
rect 1424 3271 1431 3323
rect 1483 3271 1490 3323
rect 1424 3259 1490 3271
rect 1424 3207 1431 3259
rect 1483 3207 1490 3259
rect 1424 3195 1490 3207
rect 1424 3143 1431 3195
rect 1483 3143 1490 3195
rect 1424 3131 1490 3143
rect 1424 3079 1431 3131
rect 1483 3079 1490 3131
rect 1424 3067 1490 3079
rect 1424 3015 1431 3067
rect 1483 3015 1490 3067
rect 1424 3003 1490 3015
rect 1424 2951 1431 3003
rect 1483 2951 1490 3003
rect 1424 2939 1490 2951
rect 1424 2887 1431 2939
rect 1483 2887 1490 2939
rect 1424 2875 1490 2887
rect 1424 2823 1431 2875
rect 1483 2823 1490 2875
rect 1424 2811 1490 2823
rect 1424 2759 1431 2811
rect 1483 2759 1490 2811
rect 1424 2474 1490 2759
rect 2340 6385 2406 6398
rect 2340 6333 2347 6385
rect 2399 6333 2406 6385
rect 2340 6321 2406 6333
rect 2340 6269 2347 6321
rect 2399 6269 2406 6321
rect 2340 6257 2406 6269
rect 2340 6205 2347 6257
rect 2399 6205 2406 6257
rect 2340 6193 2406 6205
rect 2340 6141 2347 6193
rect 2399 6141 2406 6193
rect 2340 6129 2406 6141
rect 2340 6077 2347 6129
rect 2399 6077 2406 6129
rect 2340 6065 2406 6077
rect 2340 6013 2347 6065
rect 2399 6013 2406 6065
rect 2340 6001 2406 6013
rect 2340 5949 2347 6001
rect 2399 5949 2406 6001
rect 2340 5937 2406 5949
rect 2340 5885 2347 5937
rect 2399 5885 2406 5937
rect 2340 5873 2406 5885
rect 2340 5821 2347 5873
rect 2399 5821 2406 5873
rect 2340 5809 2406 5821
rect 2340 5757 2347 5809
rect 2399 5757 2406 5809
rect 2340 5745 2406 5757
rect 2340 5693 2347 5745
rect 2399 5693 2406 5745
rect 2340 5681 2406 5693
rect 2340 5629 2347 5681
rect 2399 5629 2406 5681
rect 2340 5617 2406 5629
rect 2340 5565 2347 5617
rect 2399 5565 2406 5617
rect 2340 5553 2406 5565
rect 2340 5501 2347 5553
rect 2399 5501 2406 5553
rect 2340 5489 2406 5501
rect 2340 5437 2347 5489
rect 2399 5437 2406 5489
rect 2340 5425 2406 5437
rect 2340 5373 2347 5425
rect 2399 5373 2406 5425
rect 2340 5361 2406 5373
rect 2340 5309 2347 5361
rect 2399 5309 2406 5361
rect 2340 5297 2406 5309
rect 2340 5245 2347 5297
rect 2399 5245 2406 5297
rect 2340 5233 2406 5245
rect 2340 5181 2347 5233
rect 2399 5181 2406 5233
rect 2340 5169 2406 5181
rect 2340 5117 2347 5169
rect 2399 5117 2406 5169
rect 2340 5105 2406 5117
rect 2340 5053 2347 5105
rect 2399 5053 2406 5105
rect 2340 5041 2406 5053
rect 2340 4989 2347 5041
rect 2399 4989 2406 5041
rect 2340 4977 2406 4989
rect 2340 4925 2347 4977
rect 2399 4925 2406 4977
rect 2340 4913 2406 4925
rect 2340 4861 2347 4913
rect 2399 4861 2406 4913
rect 2340 4849 2406 4861
rect 2340 4797 2347 4849
rect 2399 4797 2406 4849
rect 2340 4347 2406 4797
rect 2340 4295 2347 4347
rect 2399 4295 2406 4347
rect 2340 4283 2406 4295
rect 2340 4231 2347 4283
rect 2399 4231 2406 4283
rect 2340 4219 2406 4231
rect 2340 4167 2347 4219
rect 2399 4167 2406 4219
rect 2340 4155 2406 4167
rect 2340 4103 2347 4155
rect 2399 4103 2406 4155
rect 2340 4091 2406 4103
rect 2340 4039 2347 4091
rect 2399 4039 2406 4091
rect 2340 4027 2406 4039
rect 2340 3975 2347 4027
rect 2399 3975 2406 4027
rect 2340 3963 2406 3975
rect 2340 3911 2347 3963
rect 2399 3911 2406 3963
rect 2340 3899 2406 3911
rect 2340 3847 2347 3899
rect 2399 3847 2406 3899
rect 2340 3835 2406 3847
rect 2340 3783 2347 3835
rect 2399 3783 2406 3835
rect 2340 3771 2406 3783
rect 2340 3719 2347 3771
rect 2399 3719 2406 3771
rect 2340 3707 2406 3719
rect 2340 3655 2347 3707
rect 2399 3655 2406 3707
rect 2340 3643 2406 3655
rect 2340 3591 2347 3643
rect 2399 3591 2406 3643
rect 2340 3579 2406 3591
rect 2340 3527 2347 3579
rect 2399 3527 2406 3579
rect 2340 3515 2406 3527
rect 2340 3463 2347 3515
rect 2399 3463 2406 3515
rect 2340 3451 2406 3463
rect 2340 3399 2347 3451
rect 2399 3399 2406 3451
rect 2340 3387 2406 3399
rect 2340 3335 2347 3387
rect 2399 3335 2406 3387
rect 2340 3323 2406 3335
rect 2340 3271 2347 3323
rect 2399 3271 2406 3323
rect 2340 3259 2406 3271
rect 2340 3207 2347 3259
rect 2399 3207 2406 3259
rect 2340 3195 2406 3207
rect 2340 3143 2347 3195
rect 2399 3143 2406 3195
rect 2340 3131 2406 3143
rect 2340 3079 2347 3131
rect 2399 3079 2406 3131
rect 2340 3067 2406 3079
rect 2340 3015 2347 3067
rect 2399 3015 2406 3067
rect 2340 3003 2406 3015
rect 2340 2951 2347 3003
rect 2399 2951 2406 3003
rect 2340 2939 2406 2951
rect 2340 2887 2347 2939
rect 2399 2887 2406 2939
rect 2340 2875 2406 2887
rect 2340 2823 2347 2875
rect 2399 2823 2406 2875
rect 2340 2811 2406 2823
rect 2340 2759 2347 2811
rect 2399 2759 2406 2811
rect 1638 2714 1720 2732
rect 1638 2658 1651 2714
rect 1707 2658 1720 2714
rect 1638 2640 1720 2658
rect 2340 2474 2406 2759
rect 3256 6385 3322 6398
rect 3256 6333 3263 6385
rect 3315 6333 3322 6385
rect 3256 6321 3322 6333
rect 3256 6269 3263 6321
rect 3315 6269 3322 6321
rect 3256 6257 3322 6269
rect 3256 6205 3263 6257
rect 3315 6205 3322 6257
rect 3256 6193 3322 6205
rect 3256 6141 3263 6193
rect 3315 6141 3322 6193
rect 3256 6129 3322 6141
rect 3256 6077 3263 6129
rect 3315 6077 3322 6129
rect 3256 6065 3322 6077
rect 3256 6013 3263 6065
rect 3315 6013 3322 6065
rect 3256 6001 3322 6013
rect 3256 5949 3263 6001
rect 3315 5949 3322 6001
rect 3256 5937 3322 5949
rect 3256 5885 3263 5937
rect 3315 5885 3322 5937
rect 3256 5873 3322 5885
rect 3256 5821 3263 5873
rect 3315 5821 3322 5873
rect 3256 5809 3322 5821
rect 3256 5757 3263 5809
rect 3315 5757 3322 5809
rect 3256 5745 3322 5757
rect 3256 5693 3263 5745
rect 3315 5693 3322 5745
rect 3256 5681 3322 5693
rect 3256 5629 3263 5681
rect 3315 5629 3322 5681
rect 3256 5617 3322 5629
rect 3256 5565 3263 5617
rect 3315 5565 3322 5617
rect 3256 5553 3322 5565
rect 3256 5501 3263 5553
rect 3315 5501 3322 5553
rect 3256 5489 3322 5501
rect 3256 5437 3263 5489
rect 3315 5437 3322 5489
rect 3256 5425 3322 5437
rect 3256 5373 3263 5425
rect 3315 5373 3322 5425
rect 3256 5361 3322 5373
rect 3256 5309 3263 5361
rect 3315 5309 3322 5361
rect 3256 5297 3322 5309
rect 3256 5245 3263 5297
rect 3315 5245 3322 5297
rect 3256 5233 3322 5245
rect 3256 5181 3263 5233
rect 3315 5181 3322 5233
rect 3256 5169 3322 5181
rect 3256 5117 3263 5169
rect 3315 5117 3322 5169
rect 3256 5105 3322 5117
rect 3256 5053 3263 5105
rect 3315 5053 3322 5105
rect 3256 5041 3322 5053
rect 3256 4989 3263 5041
rect 3315 4989 3322 5041
rect 3256 4977 3322 4989
rect 3256 4925 3263 4977
rect 3315 4925 3322 4977
rect 3256 4913 3322 4925
rect 3256 4861 3263 4913
rect 3315 4861 3322 4913
rect 3256 4849 3322 4861
rect 3256 4797 3263 4849
rect 3315 4797 3322 4849
rect 3256 4347 3322 4797
rect 3256 4295 3263 4347
rect 3315 4295 3322 4347
rect 3256 4283 3322 4295
rect 3256 4231 3263 4283
rect 3315 4231 3322 4283
rect 3256 4219 3322 4231
rect 3256 4167 3263 4219
rect 3315 4167 3322 4219
rect 3256 4155 3322 4167
rect 3256 4103 3263 4155
rect 3315 4103 3322 4155
rect 3256 4091 3322 4103
rect 3256 4039 3263 4091
rect 3315 4039 3322 4091
rect 3256 4027 3322 4039
rect 3256 3975 3263 4027
rect 3315 3975 3322 4027
rect 3256 3963 3322 3975
rect 3256 3911 3263 3963
rect 3315 3911 3322 3963
rect 3256 3899 3322 3911
rect 3256 3847 3263 3899
rect 3315 3847 3322 3899
rect 3256 3835 3322 3847
rect 3256 3783 3263 3835
rect 3315 3783 3322 3835
rect 3256 3771 3322 3783
rect 3256 3719 3263 3771
rect 3315 3719 3322 3771
rect 3256 3707 3322 3719
rect 3256 3655 3263 3707
rect 3315 3655 3322 3707
rect 3256 3643 3322 3655
rect 3256 3591 3263 3643
rect 3315 3591 3322 3643
rect 3256 3579 3322 3591
rect 3256 3527 3263 3579
rect 3315 3527 3322 3579
rect 3256 3515 3322 3527
rect 3256 3463 3263 3515
rect 3315 3463 3322 3515
rect 3256 3451 3322 3463
rect 3256 3399 3263 3451
rect 3315 3399 3322 3451
rect 3256 3387 3322 3399
rect 3256 3335 3263 3387
rect 3315 3335 3322 3387
rect 3256 3323 3322 3335
rect 3256 3271 3263 3323
rect 3315 3271 3322 3323
rect 3256 3259 3322 3271
rect 3256 3207 3263 3259
rect 3315 3207 3322 3259
rect 3256 3195 3322 3207
rect 3256 3143 3263 3195
rect 3315 3143 3322 3195
rect 3256 3131 3322 3143
rect 3256 3079 3263 3131
rect 3315 3079 3322 3131
rect 3256 3067 3322 3079
rect 3256 3015 3263 3067
rect 3315 3015 3322 3067
rect 3256 3003 3322 3015
rect 3256 2951 3263 3003
rect 3315 2951 3322 3003
rect 3256 2939 3322 2951
rect 3256 2887 3263 2939
rect 3315 2887 3322 2939
rect 3256 2875 3322 2887
rect 3256 2823 3263 2875
rect 3315 2823 3322 2875
rect 3256 2811 3322 2823
rect 3256 2759 3263 2811
rect 3315 2759 3322 2811
rect 3256 2474 3322 2759
rect 1424 2413 3322 2474
rect 1424 2396 1633 2413
rect 643 2035 662 2396
rect 188 2014 662 2035
rect 818 2085 898 2096
rect 818 2029 831 2085
rect 887 2029 898 2085
rect 818 2016 898 2029
rect 1378 2031 1474 2054
rect 1378 1979 1401 2031
rect 1453 1979 1474 2031
rect 1614 2041 1633 2396
rect 2069 2396 3322 2413
rect 2069 2041 2088 2396
rect 1614 2020 2088 2041
rect 1378 1950 1474 1979
rect 1016 1925 1474 1950
rect 1016 1869 1039 1925
rect 1095 1869 1474 1925
rect 1016 1852 1474 1869
rect 100 1559 164 1578
rect 100 1507 106 1559
rect 158 1507 164 1559
rect 100 1438 164 1507
rect 2616 1438 2672 1448
rect 100 1434 2708 1438
rect 100 1382 2618 1434
rect 2670 1382 2708 1434
rect 100 1378 2708 1382
rect 2616 1368 2672 1378
rect 650 1245 826 1298
rect 650 1189 711 1245
rect 767 1189 826 1245
rect 650 1101 826 1189
rect 650 1045 715 1101
rect 771 1045 826 1101
rect 650 1002 826 1045
rect 1494 1235 1670 1298
rect 1494 1179 1553 1235
rect 1609 1179 1670 1235
rect 1494 1105 1670 1179
rect 1494 1049 1551 1105
rect 1607 1049 1670 1105
rect 1494 1002 1670 1049
rect 2468 886 2524 896
rect 96 882 2704 886
rect 96 830 2470 882
rect 2522 830 2704 882
rect 96 826 2704 830
rect 96 757 160 826
rect 2468 816 2524 826
rect 96 705 102 757
rect 154 705 160 757
rect 96 686 160 705
rect 1020 299 1120 324
rect 1020 243 1043 299
rect 1099 243 1120 299
rect 1020 226 1120 243
rect 1192 301 1292 324
rect 1192 245 1211 301
rect 1267 245 1292 301
rect 1192 226 1292 245
rect -1142 0 3470 40
rect -1142 -60 -1104 0
rect -1160 -216 -1104 -60
rect 3432 -60 3470 0
rect 3432 -216 3488 -60
rect -1160 -264 3488 -216
rect -1160 -563 -1092 -264
rect -1160 -615 -1152 -563
rect -1100 -615 -1092 -563
rect -1160 -627 -1092 -615
rect -1160 -679 -1152 -627
rect -1100 -679 -1092 -627
rect -1160 -691 -1092 -679
rect -1160 -743 -1152 -691
rect -1100 -743 -1092 -691
rect -1160 -755 -1092 -743
rect -1160 -807 -1152 -755
rect -1100 -807 -1092 -755
rect -1160 -819 -1092 -807
rect -1160 -871 -1152 -819
rect -1100 -871 -1092 -819
rect -1160 -883 -1092 -871
rect -1160 -935 -1152 -883
rect -1100 -935 -1092 -883
rect -1160 -947 -1092 -935
rect -1160 -999 -1152 -947
rect -1100 -999 -1092 -947
rect -1160 -1011 -1092 -999
rect -1160 -1063 -1152 -1011
rect -1100 -1063 -1092 -1011
rect -1160 -1075 -1092 -1063
rect -1160 -1127 -1152 -1075
rect -1100 -1127 -1092 -1075
rect -1160 -1139 -1092 -1127
rect -1160 -1191 -1152 -1139
rect -1100 -1191 -1092 -1139
rect -1160 -1203 -1092 -1191
rect -1160 -1255 -1152 -1203
rect -1100 -1255 -1092 -1203
rect -1160 -1267 -1092 -1255
rect -1160 -1319 -1152 -1267
rect -1100 -1319 -1092 -1267
rect -1160 -1331 -1092 -1319
rect -1160 -1383 -1152 -1331
rect -1100 -1383 -1092 -1331
rect -1160 -1395 -1092 -1383
rect -1160 -1447 -1152 -1395
rect -1100 -1447 -1092 -1395
rect -1160 -1459 -1092 -1447
rect -1160 -1511 -1152 -1459
rect -1100 -1511 -1092 -1459
rect -1160 -1523 -1092 -1511
rect -1160 -1575 -1152 -1523
rect -1100 -1575 -1092 -1523
rect -1160 -1587 -1092 -1575
rect -1160 -1639 -1152 -1587
rect -1100 -1639 -1092 -1587
rect -1160 -1651 -1092 -1639
rect -1160 -1703 -1152 -1651
rect -1100 -1703 -1092 -1651
rect -1160 -1715 -1092 -1703
rect -1160 -1767 -1152 -1715
rect -1100 -1767 -1092 -1715
rect -1160 -1779 -1092 -1767
rect -1160 -1831 -1152 -1779
rect -1100 -1831 -1092 -1779
rect -1160 -1843 -1092 -1831
rect -1160 -1895 -1152 -1843
rect -1100 -1895 -1092 -1843
rect -1160 -1907 -1092 -1895
rect -1160 -1959 -1152 -1907
rect -1100 -1959 -1092 -1907
rect -1160 -1971 -1092 -1959
rect -1160 -2023 -1152 -1971
rect -1100 -2023 -1092 -1971
rect -1160 -2035 -1092 -2023
rect -1160 -2087 -1152 -2035
rect -1100 -2087 -1092 -2035
rect -1160 -2099 -1092 -2087
rect -1160 -2151 -1152 -2099
rect -1100 -2151 -1092 -2099
rect -1160 -2163 -1092 -2151
rect -1160 -2215 -1152 -2163
rect -1100 -2215 -1092 -2163
rect -1160 -2227 -1092 -2215
rect -1160 -2279 -1152 -2227
rect -1100 -2279 -1092 -2227
rect -1160 -2291 -1092 -2279
rect -1160 -2343 -1152 -2291
rect -1100 -2343 -1092 -2291
rect -1160 -2355 -1092 -2343
rect -1160 -2407 -1152 -2355
rect -1100 -2407 -1092 -2355
rect -1160 -2419 -1092 -2407
rect -1160 -2471 -1152 -2419
rect -1100 -2471 -1092 -2419
rect -1160 -2483 -1092 -2471
rect -1160 -2535 -1152 -2483
rect -1100 -2535 -1092 -2483
rect -1160 -2547 -1092 -2535
rect -1160 -2599 -1152 -2547
rect -1100 -2599 -1092 -2547
rect -1160 -2611 -1092 -2599
rect -1160 -2663 -1152 -2611
rect -1100 -2663 -1092 -2611
rect -1160 -2675 -1092 -2663
rect -1160 -2727 -1152 -2675
rect -1100 -2727 -1092 -2675
rect -1160 -2739 -1092 -2727
rect -1160 -2791 -1152 -2739
rect -1100 -2791 -1092 -2739
rect -1160 -2803 -1092 -2791
rect -1160 -2855 -1152 -2803
rect -1100 -2855 -1092 -2803
rect -1160 -2867 -1092 -2855
rect -1160 -2919 -1152 -2867
rect -1100 -2919 -1092 -2867
rect -1160 -2931 -1092 -2919
rect -1160 -2983 -1152 -2931
rect -1100 -2983 -1092 -2931
rect -1160 -2995 -1092 -2983
rect -1160 -3047 -1152 -2995
rect -1100 -3047 -1092 -2995
rect -1160 -3059 -1092 -3047
rect -1160 -3111 -1152 -3059
rect -1100 -3111 -1092 -3059
rect -1160 -3123 -1092 -3111
rect -1160 -3175 -1152 -3123
rect -1100 -3175 -1092 -3123
rect -1160 -3196 -1092 -3175
rect -702 -563 -634 -542
rect -702 -615 -694 -563
rect -642 -615 -634 -563
rect -702 -627 -634 -615
rect -702 -679 -694 -627
rect -642 -679 -634 -627
rect -702 -691 -634 -679
rect -702 -743 -694 -691
rect -642 -743 -634 -691
rect -702 -755 -634 -743
rect -702 -807 -694 -755
rect -642 -807 -634 -755
rect -702 -819 -634 -807
rect -702 -871 -694 -819
rect -642 -871 -634 -819
rect -702 -883 -634 -871
rect -702 -935 -694 -883
rect -642 -935 -634 -883
rect -702 -947 -634 -935
rect -702 -999 -694 -947
rect -642 -999 -634 -947
rect -702 -1011 -634 -999
rect -702 -1063 -694 -1011
rect -642 -1063 -634 -1011
rect -702 -1075 -634 -1063
rect -702 -1127 -694 -1075
rect -642 -1127 -634 -1075
rect -702 -1139 -634 -1127
rect -702 -1191 -694 -1139
rect -642 -1191 -634 -1139
rect -702 -1203 -634 -1191
rect -702 -1255 -694 -1203
rect -642 -1255 -634 -1203
rect -702 -1267 -634 -1255
rect -702 -1319 -694 -1267
rect -642 -1319 -634 -1267
rect -702 -1331 -634 -1319
rect -702 -1383 -694 -1331
rect -642 -1383 -634 -1331
rect -702 -1395 -634 -1383
rect -702 -1447 -694 -1395
rect -642 -1447 -634 -1395
rect -702 -1459 -634 -1447
rect -702 -1511 -694 -1459
rect -642 -1511 -634 -1459
rect -702 -1523 -634 -1511
rect -702 -1575 -694 -1523
rect -642 -1575 -634 -1523
rect -702 -1587 -634 -1575
rect -702 -1639 -694 -1587
rect -642 -1639 -634 -1587
rect -702 -1651 -634 -1639
rect -702 -1703 -694 -1651
rect -642 -1703 -634 -1651
rect -702 -1715 -634 -1703
rect -702 -1767 -694 -1715
rect -642 -1767 -634 -1715
rect -702 -1779 -634 -1767
rect -702 -1831 -694 -1779
rect -642 -1831 -634 -1779
rect -702 -1843 -634 -1831
rect -702 -1895 -694 -1843
rect -642 -1895 -634 -1843
rect -702 -1907 -634 -1895
rect -702 -1959 -694 -1907
rect -642 -1959 -634 -1907
rect -702 -1971 -634 -1959
rect -702 -2023 -694 -1971
rect -642 -2023 -634 -1971
rect -702 -2035 -634 -2023
rect -702 -2087 -694 -2035
rect -642 -2087 -634 -2035
rect -702 -2099 -634 -2087
rect -702 -2151 -694 -2099
rect -642 -2151 -634 -2099
rect -702 -2163 -634 -2151
rect -702 -2215 -694 -2163
rect -642 -2215 -634 -2163
rect -702 -2227 -634 -2215
rect -702 -2279 -694 -2227
rect -642 -2279 -634 -2227
rect -702 -2291 -634 -2279
rect -702 -2343 -694 -2291
rect -642 -2343 -634 -2291
rect -702 -2355 -634 -2343
rect -702 -2407 -694 -2355
rect -642 -2407 -634 -2355
rect -702 -2419 -634 -2407
rect -702 -2471 -694 -2419
rect -642 -2471 -634 -2419
rect -702 -2483 -634 -2471
rect -702 -2535 -694 -2483
rect -642 -2535 -634 -2483
rect -702 -2547 -634 -2535
rect -702 -2599 -694 -2547
rect -642 -2599 -634 -2547
rect -702 -2611 -634 -2599
rect -702 -2663 -694 -2611
rect -642 -2663 -634 -2611
rect -702 -2675 -634 -2663
rect -702 -2727 -694 -2675
rect -642 -2727 -634 -2675
rect -702 -2739 -634 -2727
rect -702 -2791 -694 -2739
rect -642 -2791 -634 -2739
rect -702 -2803 -634 -2791
rect -702 -2855 -694 -2803
rect -642 -2855 -634 -2803
rect -702 -2867 -634 -2855
rect -702 -2919 -694 -2867
rect -642 -2919 -634 -2867
rect -702 -2931 -634 -2919
rect -702 -2983 -694 -2931
rect -642 -2983 -634 -2931
rect -702 -2995 -634 -2983
rect -702 -3047 -694 -2995
rect -642 -3047 -634 -2995
rect -702 -3059 -634 -3047
rect -702 -3111 -694 -3059
rect -642 -3111 -634 -3059
rect -702 -3123 -634 -3111
rect -702 -3175 -694 -3123
rect -642 -3175 -634 -3123
rect -702 -3472 -634 -3175
rect -244 -563 -176 -264
rect -244 -615 -236 -563
rect -184 -615 -176 -563
rect -244 -627 -176 -615
rect -244 -679 -236 -627
rect -184 -679 -176 -627
rect -244 -691 -176 -679
rect -244 -743 -236 -691
rect -184 -743 -176 -691
rect -244 -755 -176 -743
rect -244 -807 -236 -755
rect -184 -807 -176 -755
rect -244 -819 -176 -807
rect -244 -871 -236 -819
rect -184 -871 -176 -819
rect -244 -883 -176 -871
rect -244 -935 -236 -883
rect -184 -935 -176 -883
rect -244 -947 -176 -935
rect -244 -999 -236 -947
rect -184 -999 -176 -947
rect -244 -1011 -176 -999
rect -244 -1063 -236 -1011
rect -184 -1063 -176 -1011
rect -244 -1075 -176 -1063
rect -244 -1127 -236 -1075
rect -184 -1127 -176 -1075
rect -244 -1139 -176 -1127
rect -244 -1191 -236 -1139
rect -184 -1191 -176 -1139
rect -244 -1203 -176 -1191
rect -244 -1255 -236 -1203
rect -184 -1255 -176 -1203
rect -244 -1267 -176 -1255
rect -244 -1319 -236 -1267
rect -184 -1319 -176 -1267
rect -244 -1331 -176 -1319
rect -244 -1383 -236 -1331
rect -184 -1383 -176 -1331
rect -244 -1395 -176 -1383
rect -244 -1447 -236 -1395
rect -184 -1447 -176 -1395
rect -244 -1459 -176 -1447
rect -244 -1511 -236 -1459
rect -184 -1511 -176 -1459
rect -244 -1523 -176 -1511
rect -244 -1575 -236 -1523
rect -184 -1575 -176 -1523
rect -244 -1587 -176 -1575
rect -244 -1639 -236 -1587
rect -184 -1639 -176 -1587
rect -244 -1651 -176 -1639
rect -244 -1703 -236 -1651
rect -184 -1703 -176 -1651
rect -244 -1715 -176 -1703
rect -244 -1767 -236 -1715
rect -184 -1767 -176 -1715
rect -244 -1779 -176 -1767
rect -244 -1831 -236 -1779
rect -184 -1831 -176 -1779
rect -244 -1843 -176 -1831
rect -244 -1895 -236 -1843
rect -184 -1895 -176 -1843
rect -244 -1907 -176 -1895
rect -244 -1959 -236 -1907
rect -184 -1959 -176 -1907
rect -244 -1971 -176 -1959
rect -244 -2023 -236 -1971
rect -184 -2023 -176 -1971
rect -244 -2035 -176 -2023
rect -244 -2087 -236 -2035
rect -184 -2087 -176 -2035
rect -244 -2099 -176 -2087
rect -244 -2151 -236 -2099
rect -184 -2151 -176 -2099
rect -244 -2163 -176 -2151
rect -244 -2215 -236 -2163
rect -184 -2215 -176 -2163
rect -244 -2227 -176 -2215
rect -244 -2279 -236 -2227
rect -184 -2279 -176 -2227
rect -244 -2291 -176 -2279
rect -244 -2343 -236 -2291
rect -184 -2343 -176 -2291
rect -244 -2355 -176 -2343
rect -244 -2407 -236 -2355
rect -184 -2407 -176 -2355
rect -244 -2419 -176 -2407
rect -244 -2471 -236 -2419
rect -184 -2471 -176 -2419
rect -244 -2483 -176 -2471
rect -244 -2535 -236 -2483
rect -184 -2535 -176 -2483
rect -244 -2547 -176 -2535
rect -244 -2599 -236 -2547
rect -184 -2599 -176 -2547
rect -244 -2611 -176 -2599
rect -244 -2663 -236 -2611
rect -184 -2663 -176 -2611
rect -244 -2675 -176 -2663
rect -244 -2727 -236 -2675
rect -184 -2727 -176 -2675
rect -244 -2739 -176 -2727
rect -244 -2791 -236 -2739
rect -184 -2791 -176 -2739
rect -244 -2803 -176 -2791
rect -244 -2855 -236 -2803
rect -184 -2855 -176 -2803
rect -244 -2867 -176 -2855
rect -244 -2919 -236 -2867
rect -184 -2919 -176 -2867
rect -244 -2931 -176 -2919
rect -244 -2983 -236 -2931
rect -184 -2983 -176 -2931
rect -244 -2995 -176 -2983
rect -244 -3047 -236 -2995
rect -184 -3047 -176 -2995
rect -244 -3059 -176 -3047
rect -244 -3111 -236 -3059
rect -184 -3111 -176 -3059
rect -244 -3123 -176 -3111
rect -244 -3175 -236 -3123
rect -184 -3175 -176 -3123
rect -244 -3196 -176 -3175
rect 214 -563 282 -542
rect 214 -615 222 -563
rect 274 -615 282 -563
rect 214 -627 282 -615
rect 214 -679 222 -627
rect 274 -679 282 -627
rect 214 -691 282 -679
rect 214 -743 222 -691
rect 274 -743 282 -691
rect 214 -755 282 -743
rect 214 -807 222 -755
rect 274 -807 282 -755
rect 214 -819 282 -807
rect 214 -871 222 -819
rect 274 -871 282 -819
rect 214 -883 282 -871
rect 214 -935 222 -883
rect 274 -935 282 -883
rect 214 -947 282 -935
rect 214 -999 222 -947
rect 274 -999 282 -947
rect 214 -1011 282 -999
rect 214 -1063 222 -1011
rect 274 -1063 282 -1011
rect 214 -1075 282 -1063
rect 214 -1127 222 -1075
rect 274 -1127 282 -1075
rect 214 -1139 282 -1127
rect 214 -1191 222 -1139
rect 274 -1191 282 -1139
rect 214 -1203 282 -1191
rect 214 -1255 222 -1203
rect 274 -1255 282 -1203
rect 214 -1267 282 -1255
rect 214 -1319 222 -1267
rect 274 -1319 282 -1267
rect 214 -1331 282 -1319
rect 214 -1383 222 -1331
rect 274 -1383 282 -1331
rect 214 -1395 282 -1383
rect 214 -1447 222 -1395
rect 274 -1447 282 -1395
rect 214 -1459 282 -1447
rect 214 -1511 222 -1459
rect 274 -1511 282 -1459
rect 214 -1523 282 -1511
rect 214 -1575 222 -1523
rect 274 -1575 282 -1523
rect 214 -1587 282 -1575
rect 214 -1639 222 -1587
rect 274 -1639 282 -1587
rect 214 -1651 282 -1639
rect 214 -1703 222 -1651
rect 274 -1703 282 -1651
rect 214 -1715 282 -1703
rect 214 -1767 222 -1715
rect 274 -1767 282 -1715
rect 214 -1779 282 -1767
rect 214 -1831 222 -1779
rect 274 -1831 282 -1779
rect 214 -1843 282 -1831
rect 214 -1895 222 -1843
rect 274 -1895 282 -1843
rect 214 -1907 282 -1895
rect 214 -1959 222 -1907
rect 274 -1959 282 -1907
rect 214 -1971 282 -1959
rect 214 -2023 222 -1971
rect 274 -2023 282 -1971
rect 214 -2035 282 -2023
rect 214 -2087 222 -2035
rect 274 -2087 282 -2035
rect 214 -2099 282 -2087
rect 214 -2151 222 -2099
rect 274 -2151 282 -2099
rect 214 -2163 282 -2151
rect 214 -2215 222 -2163
rect 274 -2215 282 -2163
rect 214 -2227 282 -2215
rect 214 -2279 222 -2227
rect 274 -2279 282 -2227
rect 214 -2291 282 -2279
rect 214 -2343 222 -2291
rect 274 -2343 282 -2291
rect 214 -2355 282 -2343
rect 214 -2407 222 -2355
rect 274 -2407 282 -2355
rect 214 -2419 282 -2407
rect 214 -2471 222 -2419
rect 274 -2471 282 -2419
rect 214 -2483 282 -2471
rect 214 -2535 222 -2483
rect 274 -2535 282 -2483
rect 214 -2547 282 -2535
rect 214 -2599 222 -2547
rect 274 -2599 282 -2547
rect 214 -2611 282 -2599
rect 214 -2663 222 -2611
rect 274 -2663 282 -2611
rect 214 -2675 282 -2663
rect 214 -2727 222 -2675
rect 274 -2727 282 -2675
rect 214 -2739 282 -2727
rect 214 -2791 222 -2739
rect 274 -2791 282 -2739
rect 214 -2803 282 -2791
rect 214 -2855 222 -2803
rect 274 -2855 282 -2803
rect 214 -2867 282 -2855
rect 214 -2919 222 -2867
rect 274 -2919 282 -2867
rect 214 -2931 282 -2919
rect 214 -2983 222 -2931
rect 274 -2983 282 -2931
rect 214 -2995 282 -2983
rect 214 -3047 222 -2995
rect 274 -3047 282 -2995
rect 214 -3059 282 -3047
rect 214 -3111 222 -3059
rect 274 -3111 282 -3059
rect 214 -3123 282 -3111
rect 214 -3175 222 -3123
rect 274 -3175 282 -3123
rect 214 -3472 282 -3175
rect 672 -563 740 -264
rect 672 -615 680 -563
rect 732 -615 740 -563
rect 672 -627 740 -615
rect 672 -679 680 -627
rect 732 -679 740 -627
rect 672 -691 740 -679
rect 672 -743 680 -691
rect 732 -743 740 -691
rect 672 -755 740 -743
rect 672 -807 680 -755
rect 732 -807 740 -755
rect 672 -819 740 -807
rect 672 -871 680 -819
rect 732 -871 740 -819
rect 672 -883 740 -871
rect 672 -935 680 -883
rect 732 -935 740 -883
rect 672 -947 740 -935
rect 672 -999 680 -947
rect 732 -999 740 -947
rect 672 -1011 740 -999
rect 672 -1063 680 -1011
rect 732 -1063 740 -1011
rect 672 -1075 740 -1063
rect 672 -1127 680 -1075
rect 732 -1127 740 -1075
rect 672 -1139 740 -1127
rect 672 -1191 680 -1139
rect 732 -1191 740 -1139
rect 672 -1203 740 -1191
rect 672 -1255 680 -1203
rect 732 -1255 740 -1203
rect 672 -1267 740 -1255
rect 672 -1319 680 -1267
rect 732 -1319 740 -1267
rect 672 -1331 740 -1319
rect 672 -1383 680 -1331
rect 732 -1383 740 -1331
rect 672 -1395 740 -1383
rect 672 -1447 680 -1395
rect 732 -1447 740 -1395
rect 672 -1459 740 -1447
rect 672 -1511 680 -1459
rect 732 -1511 740 -1459
rect 672 -1523 740 -1511
rect 672 -1575 680 -1523
rect 732 -1575 740 -1523
rect 672 -1587 740 -1575
rect 672 -1639 680 -1587
rect 732 -1639 740 -1587
rect 672 -1651 740 -1639
rect 672 -1703 680 -1651
rect 732 -1703 740 -1651
rect 672 -1715 740 -1703
rect 672 -1767 680 -1715
rect 732 -1767 740 -1715
rect 672 -1779 740 -1767
rect 672 -1831 680 -1779
rect 732 -1831 740 -1779
rect 672 -1843 740 -1831
rect 672 -1895 680 -1843
rect 732 -1895 740 -1843
rect 672 -1907 740 -1895
rect 672 -1959 680 -1907
rect 732 -1959 740 -1907
rect 672 -1971 740 -1959
rect 672 -2023 680 -1971
rect 732 -2023 740 -1971
rect 672 -2035 740 -2023
rect 672 -2087 680 -2035
rect 732 -2087 740 -2035
rect 672 -2099 740 -2087
rect 672 -2151 680 -2099
rect 732 -2151 740 -2099
rect 672 -2163 740 -2151
rect 672 -2215 680 -2163
rect 732 -2215 740 -2163
rect 672 -2227 740 -2215
rect 672 -2279 680 -2227
rect 732 -2279 740 -2227
rect 672 -2291 740 -2279
rect 672 -2343 680 -2291
rect 732 -2343 740 -2291
rect 672 -2355 740 -2343
rect 672 -2407 680 -2355
rect 732 -2407 740 -2355
rect 672 -2419 740 -2407
rect 672 -2471 680 -2419
rect 732 -2471 740 -2419
rect 672 -2483 740 -2471
rect 672 -2535 680 -2483
rect 732 -2535 740 -2483
rect 672 -2547 740 -2535
rect 672 -2599 680 -2547
rect 732 -2599 740 -2547
rect 672 -2611 740 -2599
rect 672 -2663 680 -2611
rect 732 -2663 740 -2611
rect 672 -2675 740 -2663
rect 672 -2727 680 -2675
rect 732 -2727 740 -2675
rect 672 -2739 740 -2727
rect 672 -2791 680 -2739
rect 732 -2791 740 -2739
rect 672 -2803 740 -2791
rect 672 -2855 680 -2803
rect 732 -2855 740 -2803
rect 672 -2867 740 -2855
rect 672 -2919 680 -2867
rect 732 -2919 740 -2867
rect 672 -2931 740 -2919
rect 672 -2983 680 -2931
rect 732 -2983 740 -2931
rect 672 -2995 740 -2983
rect 672 -3047 680 -2995
rect 732 -3047 740 -2995
rect 672 -3059 740 -3047
rect 672 -3111 680 -3059
rect 732 -3111 740 -3059
rect 672 -3123 740 -3111
rect 672 -3175 680 -3123
rect 732 -3175 740 -3123
rect 672 -3196 740 -3175
rect 1130 -563 1198 -542
rect 1130 -615 1138 -563
rect 1190 -615 1198 -563
rect 1130 -627 1198 -615
rect 1130 -679 1138 -627
rect 1190 -679 1198 -627
rect 1130 -691 1198 -679
rect 1130 -743 1138 -691
rect 1190 -743 1198 -691
rect 1130 -755 1198 -743
rect 1130 -807 1138 -755
rect 1190 -807 1198 -755
rect 1130 -819 1198 -807
rect 1130 -871 1138 -819
rect 1190 -871 1198 -819
rect 1130 -883 1198 -871
rect 1130 -935 1138 -883
rect 1190 -935 1198 -883
rect 1130 -947 1198 -935
rect 1130 -999 1138 -947
rect 1190 -999 1198 -947
rect 1130 -1011 1198 -999
rect 1130 -1063 1138 -1011
rect 1190 -1063 1198 -1011
rect 1130 -1075 1198 -1063
rect 1130 -1127 1138 -1075
rect 1190 -1127 1198 -1075
rect 1130 -1139 1198 -1127
rect 1130 -1191 1138 -1139
rect 1190 -1191 1198 -1139
rect 1130 -1203 1198 -1191
rect 1130 -1255 1138 -1203
rect 1190 -1255 1198 -1203
rect 1130 -1267 1198 -1255
rect 1130 -1319 1138 -1267
rect 1190 -1319 1198 -1267
rect 1130 -1331 1198 -1319
rect 1130 -1383 1138 -1331
rect 1190 -1383 1198 -1331
rect 1130 -1395 1198 -1383
rect 1130 -1447 1138 -1395
rect 1190 -1447 1198 -1395
rect 1130 -1459 1198 -1447
rect 1130 -1511 1138 -1459
rect 1190 -1511 1198 -1459
rect 1130 -1523 1198 -1511
rect 1130 -1575 1138 -1523
rect 1190 -1575 1198 -1523
rect 1130 -1587 1198 -1575
rect 1130 -1639 1138 -1587
rect 1190 -1639 1198 -1587
rect 1130 -1651 1198 -1639
rect 1130 -1703 1138 -1651
rect 1190 -1703 1198 -1651
rect 1130 -1715 1198 -1703
rect 1130 -1767 1138 -1715
rect 1190 -1767 1198 -1715
rect 1130 -1779 1198 -1767
rect 1130 -1831 1138 -1779
rect 1190 -1831 1198 -1779
rect 1130 -1843 1198 -1831
rect 1130 -1895 1138 -1843
rect 1190 -1895 1198 -1843
rect 1130 -1907 1198 -1895
rect 1130 -1959 1138 -1907
rect 1190 -1959 1198 -1907
rect 1130 -1971 1198 -1959
rect 1130 -2023 1138 -1971
rect 1190 -2023 1198 -1971
rect 1130 -2035 1198 -2023
rect 1130 -2087 1138 -2035
rect 1190 -2087 1198 -2035
rect 1130 -2099 1198 -2087
rect 1130 -2151 1138 -2099
rect 1190 -2151 1198 -2099
rect 1130 -2163 1198 -2151
rect 1130 -2215 1138 -2163
rect 1190 -2215 1198 -2163
rect 1130 -2227 1198 -2215
rect 1130 -2279 1138 -2227
rect 1190 -2279 1198 -2227
rect 1130 -2291 1198 -2279
rect 1130 -2343 1138 -2291
rect 1190 -2343 1198 -2291
rect 1130 -2355 1198 -2343
rect 1130 -2407 1138 -2355
rect 1190 -2407 1198 -2355
rect 1130 -2419 1198 -2407
rect 1130 -2471 1138 -2419
rect 1190 -2471 1198 -2419
rect 1130 -2483 1198 -2471
rect 1130 -2535 1138 -2483
rect 1190 -2535 1198 -2483
rect 1130 -2547 1198 -2535
rect 1130 -2599 1138 -2547
rect 1190 -2599 1198 -2547
rect 1130 -2611 1198 -2599
rect 1130 -2663 1138 -2611
rect 1190 -2663 1198 -2611
rect 1130 -2675 1198 -2663
rect 1130 -2727 1138 -2675
rect 1190 -2727 1198 -2675
rect 1130 -2739 1198 -2727
rect 1130 -2791 1138 -2739
rect 1190 -2791 1198 -2739
rect 1130 -2803 1198 -2791
rect 1130 -2855 1138 -2803
rect 1190 -2855 1198 -2803
rect 1130 -2867 1198 -2855
rect 1130 -2919 1138 -2867
rect 1190 -2919 1198 -2867
rect 1130 -2931 1198 -2919
rect 1130 -2983 1138 -2931
rect 1190 -2983 1198 -2931
rect 1130 -2995 1198 -2983
rect 1130 -3047 1138 -2995
rect 1190 -3047 1198 -2995
rect 1130 -3059 1198 -3047
rect 1130 -3111 1138 -3059
rect 1190 -3111 1198 -3059
rect 1130 -3123 1198 -3111
rect 1130 -3175 1138 -3123
rect 1190 -3175 1198 -3123
rect 1130 -3472 1198 -3175
rect 1588 -563 1656 -264
rect 1588 -615 1596 -563
rect 1648 -615 1656 -563
rect 1588 -627 1656 -615
rect 1588 -679 1596 -627
rect 1648 -679 1656 -627
rect 1588 -691 1656 -679
rect 1588 -743 1596 -691
rect 1648 -743 1656 -691
rect 1588 -755 1656 -743
rect 1588 -807 1596 -755
rect 1648 -807 1656 -755
rect 1588 -819 1656 -807
rect 1588 -871 1596 -819
rect 1648 -871 1656 -819
rect 1588 -883 1656 -871
rect 1588 -935 1596 -883
rect 1648 -935 1656 -883
rect 1588 -947 1656 -935
rect 1588 -999 1596 -947
rect 1648 -999 1656 -947
rect 1588 -1011 1656 -999
rect 1588 -1063 1596 -1011
rect 1648 -1063 1656 -1011
rect 1588 -1075 1656 -1063
rect 1588 -1127 1596 -1075
rect 1648 -1127 1656 -1075
rect 1588 -1139 1656 -1127
rect 1588 -1191 1596 -1139
rect 1648 -1191 1656 -1139
rect 1588 -1203 1656 -1191
rect 1588 -1255 1596 -1203
rect 1648 -1255 1656 -1203
rect 1588 -1267 1656 -1255
rect 1588 -1319 1596 -1267
rect 1648 -1319 1656 -1267
rect 1588 -1331 1656 -1319
rect 1588 -1383 1596 -1331
rect 1648 -1383 1656 -1331
rect 1588 -1395 1656 -1383
rect 1588 -1447 1596 -1395
rect 1648 -1447 1656 -1395
rect 1588 -1459 1656 -1447
rect 1588 -1511 1596 -1459
rect 1648 -1511 1656 -1459
rect 1588 -1523 1656 -1511
rect 1588 -1575 1596 -1523
rect 1648 -1575 1656 -1523
rect 1588 -1587 1656 -1575
rect 1588 -1639 1596 -1587
rect 1648 -1639 1656 -1587
rect 1588 -1651 1656 -1639
rect 1588 -1703 1596 -1651
rect 1648 -1703 1656 -1651
rect 1588 -1715 1656 -1703
rect 1588 -1767 1596 -1715
rect 1648 -1767 1656 -1715
rect 1588 -1779 1656 -1767
rect 1588 -1831 1596 -1779
rect 1648 -1831 1656 -1779
rect 1588 -1843 1656 -1831
rect 1588 -1895 1596 -1843
rect 1648 -1895 1656 -1843
rect 1588 -1907 1656 -1895
rect 1588 -1959 1596 -1907
rect 1648 -1959 1656 -1907
rect 1588 -1971 1656 -1959
rect 1588 -2023 1596 -1971
rect 1648 -2023 1656 -1971
rect 1588 -2035 1656 -2023
rect 1588 -2087 1596 -2035
rect 1648 -2087 1656 -2035
rect 1588 -2099 1656 -2087
rect 1588 -2151 1596 -2099
rect 1648 -2151 1656 -2099
rect 1588 -2163 1656 -2151
rect 1588 -2215 1596 -2163
rect 1648 -2215 1656 -2163
rect 1588 -2227 1656 -2215
rect 1588 -2279 1596 -2227
rect 1648 -2279 1656 -2227
rect 1588 -2291 1656 -2279
rect 1588 -2343 1596 -2291
rect 1648 -2343 1656 -2291
rect 1588 -2355 1656 -2343
rect 1588 -2407 1596 -2355
rect 1648 -2407 1656 -2355
rect 1588 -2419 1656 -2407
rect 1588 -2471 1596 -2419
rect 1648 -2471 1656 -2419
rect 1588 -2483 1656 -2471
rect 1588 -2535 1596 -2483
rect 1648 -2535 1656 -2483
rect 1588 -2547 1656 -2535
rect 1588 -2599 1596 -2547
rect 1648 -2599 1656 -2547
rect 1588 -2611 1656 -2599
rect 1588 -2663 1596 -2611
rect 1648 -2663 1656 -2611
rect 1588 -2675 1656 -2663
rect 1588 -2727 1596 -2675
rect 1648 -2727 1656 -2675
rect 1588 -2739 1656 -2727
rect 1588 -2791 1596 -2739
rect 1648 -2791 1656 -2739
rect 1588 -2803 1656 -2791
rect 1588 -2855 1596 -2803
rect 1648 -2855 1656 -2803
rect 1588 -2867 1656 -2855
rect 1588 -2919 1596 -2867
rect 1648 -2919 1656 -2867
rect 1588 -2931 1656 -2919
rect 1588 -2983 1596 -2931
rect 1648 -2983 1656 -2931
rect 1588 -2995 1656 -2983
rect 1588 -3047 1596 -2995
rect 1648 -3047 1656 -2995
rect 1588 -3059 1656 -3047
rect 1588 -3111 1596 -3059
rect 1648 -3111 1656 -3059
rect 1588 -3123 1656 -3111
rect 1588 -3175 1596 -3123
rect 1648 -3175 1656 -3123
rect 1588 -3196 1656 -3175
rect 2046 -563 2114 -542
rect 2046 -615 2054 -563
rect 2106 -615 2114 -563
rect 2046 -627 2114 -615
rect 2046 -679 2054 -627
rect 2106 -679 2114 -627
rect 2046 -691 2114 -679
rect 2046 -743 2054 -691
rect 2106 -743 2114 -691
rect 2046 -755 2114 -743
rect 2046 -807 2054 -755
rect 2106 -807 2114 -755
rect 2046 -819 2114 -807
rect 2046 -871 2054 -819
rect 2106 -871 2114 -819
rect 2046 -883 2114 -871
rect 2046 -935 2054 -883
rect 2106 -935 2114 -883
rect 2046 -947 2114 -935
rect 2046 -999 2054 -947
rect 2106 -999 2114 -947
rect 2046 -1011 2114 -999
rect 2046 -1063 2054 -1011
rect 2106 -1063 2114 -1011
rect 2046 -1075 2114 -1063
rect 2046 -1127 2054 -1075
rect 2106 -1127 2114 -1075
rect 2046 -1139 2114 -1127
rect 2046 -1191 2054 -1139
rect 2106 -1191 2114 -1139
rect 2046 -1203 2114 -1191
rect 2046 -1255 2054 -1203
rect 2106 -1255 2114 -1203
rect 2046 -1267 2114 -1255
rect 2046 -1319 2054 -1267
rect 2106 -1319 2114 -1267
rect 2046 -1331 2114 -1319
rect 2046 -1383 2054 -1331
rect 2106 -1383 2114 -1331
rect 2046 -1395 2114 -1383
rect 2046 -1447 2054 -1395
rect 2106 -1447 2114 -1395
rect 2046 -1459 2114 -1447
rect 2046 -1511 2054 -1459
rect 2106 -1511 2114 -1459
rect 2046 -1523 2114 -1511
rect 2046 -1575 2054 -1523
rect 2106 -1575 2114 -1523
rect 2046 -1587 2114 -1575
rect 2046 -1639 2054 -1587
rect 2106 -1639 2114 -1587
rect 2046 -1651 2114 -1639
rect 2046 -1703 2054 -1651
rect 2106 -1703 2114 -1651
rect 2046 -1715 2114 -1703
rect 2046 -1767 2054 -1715
rect 2106 -1767 2114 -1715
rect 2046 -1779 2114 -1767
rect 2046 -1831 2054 -1779
rect 2106 -1831 2114 -1779
rect 2046 -1843 2114 -1831
rect 2046 -1895 2054 -1843
rect 2106 -1895 2114 -1843
rect 2046 -1907 2114 -1895
rect 2046 -1959 2054 -1907
rect 2106 -1959 2114 -1907
rect 2046 -1971 2114 -1959
rect 2046 -2023 2054 -1971
rect 2106 -2023 2114 -1971
rect 2046 -2035 2114 -2023
rect 2046 -2087 2054 -2035
rect 2106 -2087 2114 -2035
rect 2046 -2099 2114 -2087
rect 2046 -2151 2054 -2099
rect 2106 -2151 2114 -2099
rect 2046 -2163 2114 -2151
rect 2046 -2215 2054 -2163
rect 2106 -2215 2114 -2163
rect 2046 -2227 2114 -2215
rect 2046 -2279 2054 -2227
rect 2106 -2279 2114 -2227
rect 2046 -2291 2114 -2279
rect 2046 -2343 2054 -2291
rect 2106 -2343 2114 -2291
rect 2046 -2355 2114 -2343
rect 2046 -2407 2054 -2355
rect 2106 -2407 2114 -2355
rect 2046 -2419 2114 -2407
rect 2046 -2471 2054 -2419
rect 2106 -2471 2114 -2419
rect 2046 -2483 2114 -2471
rect 2046 -2535 2054 -2483
rect 2106 -2535 2114 -2483
rect 2046 -2547 2114 -2535
rect 2046 -2599 2054 -2547
rect 2106 -2599 2114 -2547
rect 2046 -2611 2114 -2599
rect 2046 -2663 2054 -2611
rect 2106 -2663 2114 -2611
rect 2046 -2675 2114 -2663
rect 2046 -2727 2054 -2675
rect 2106 -2727 2114 -2675
rect 2046 -2739 2114 -2727
rect 2046 -2791 2054 -2739
rect 2106 -2791 2114 -2739
rect 2046 -2803 2114 -2791
rect 2046 -2855 2054 -2803
rect 2106 -2855 2114 -2803
rect 2046 -2867 2114 -2855
rect 2046 -2919 2054 -2867
rect 2106 -2919 2114 -2867
rect 2046 -2931 2114 -2919
rect 2046 -2983 2054 -2931
rect 2106 -2983 2114 -2931
rect 2046 -2995 2114 -2983
rect 2046 -3047 2054 -2995
rect 2106 -3047 2114 -2995
rect 2046 -3059 2114 -3047
rect 2046 -3111 2054 -3059
rect 2106 -3111 2114 -3059
rect 2046 -3123 2114 -3111
rect 2046 -3175 2054 -3123
rect 2106 -3175 2114 -3123
rect 2046 -3472 2114 -3175
rect 2504 -563 2572 -264
rect 2504 -615 2512 -563
rect 2564 -615 2572 -563
rect 2504 -627 2572 -615
rect 2504 -679 2512 -627
rect 2564 -679 2572 -627
rect 2504 -691 2572 -679
rect 2504 -743 2512 -691
rect 2564 -743 2572 -691
rect 2504 -755 2572 -743
rect 2504 -807 2512 -755
rect 2564 -807 2572 -755
rect 2504 -819 2572 -807
rect 2504 -871 2512 -819
rect 2564 -871 2572 -819
rect 2504 -883 2572 -871
rect 2504 -935 2512 -883
rect 2564 -935 2572 -883
rect 2504 -947 2572 -935
rect 2504 -999 2512 -947
rect 2564 -999 2572 -947
rect 2504 -1011 2572 -999
rect 2504 -1063 2512 -1011
rect 2564 -1063 2572 -1011
rect 2504 -1075 2572 -1063
rect 2504 -1127 2512 -1075
rect 2564 -1127 2572 -1075
rect 2504 -1139 2572 -1127
rect 2504 -1191 2512 -1139
rect 2564 -1191 2572 -1139
rect 2504 -1203 2572 -1191
rect 2504 -1255 2512 -1203
rect 2564 -1255 2572 -1203
rect 2504 -1267 2572 -1255
rect 2504 -1319 2512 -1267
rect 2564 -1319 2572 -1267
rect 2504 -1331 2572 -1319
rect 2504 -1383 2512 -1331
rect 2564 -1383 2572 -1331
rect 2504 -1395 2572 -1383
rect 2504 -1447 2512 -1395
rect 2564 -1447 2572 -1395
rect 2504 -1459 2572 -1447
rect 2504 -1511 2512 -1459
rect 2564 -1511 2572 -1459
rect 2504 -1523 2572 -1511
rect 2504 -1575 2512 -1523
rect 2564 -1575 2572 -1523
rect 2504 -1587 2572 -1575
rect 2504 -1639 2512 -1587
rect 2564 -1639 2572 -1587
rect 2504 -1651 2572 -1639
rect 2504 -1703 2512 -1651
rect 2564 -1703 2572 -1651
rect 2504 -1715 2572 -1703
rect 2504 -1767 2512 -1715
rect 2564 -1767 2572 -1715
rect 2504 -1779 2572 -1767
rect 2504 -1831 2512 -1779
rect 2564 -1831 2572 -1779
rect 2504 -1843 2572 -1831
rect 2504 -1895 2512 -1843
rect 2564 -1895 2572 -1843
rect 2504 -1907 2572 -1895
rect 2504 -1959 2512 -1907
rect 2564 -1959 2572 -1907
rect 2504 -1971 2572 -1959
rect 2504 -2023 2512 -1971
rect 2564 -2023 2572 -1971
rect 2504 -2035 2572 -2023
rect 2504 -2087 2512 -2035
rect 2564 -2087 2572 -2035
rect 2504 -2099 2572 -2087
rect 2504 -2151 2512 -2099
rect 2564 -2151 2572 -2099
rect 2504 -2163 2572 -2151
rect 2504 -2215 2512 -2163
rect 2564 -2215 2572 -2163
rect 2504 -2227 2572 -2215
rect 2504 -2279 2512 -2227
rect 2564 -2279 2572 -2227
rect 2504 -2291 2572 -2279
rect 2504 -2343 2512 -2291
rect 2564 -2343 2572 -2291
rect 2504 -2355 2572 -2343
rect 2504 -2407 2512 -2355
rect 2564 -2407 2572 -2355
rect 2504 -2419 2572 -2407
rect 2504 -2471 2512 -2419
rect 2564 -2471 2572 -2419
rect 2504 -2483 2572 -2471
rect 2504 -2535 2512 -2483
rect 2564 -2535 2572 -2483
rect 2504 -2547 2572 -2535
rect 2504 -2599 2512 -2547
rect 2564 -2599 2572 -2547
rect 2504 -2611 2572 -2599
rect 2504 -2663 2512 -2611
rect 2564 -2663 2572 -2611
rect 2504 -2675 2572 -2663
rect 2504 -2727 2512 -2675
rect 2564 -2727 2572 -2675
rect 2504 -2739 2572 -2727
rect 2504 -2791 2512 -2739
rect 2564 -2791 2572 -2739
rect 2504 -2803 2572 -2791
rect 2504 -2855 2512 -2803
rect 2564 -2855 2572 -2803
rect 2504 -2867 2572 -2855
rect 2504 -2919 2512 -2867
rect 2564 -2919 2572 -2867
rect 2504 -2931 2572 -2919
rect 2504 -2983 2512 -2931
rect 2564 -2983 2572 -2931
rect 2504 -2995 2572 -2983
rect 2504 -3047 2512 -2995
rect 2564 -3047 2572 -2995
rect 2504 -3059 2572 -3047
rect 2504 -3111 2512 -3059
rect 2564 -3111 2572 -3059
rect 2504 -3123 2572 -3111
rect 2504 -3175 2512 -3123
rect 2564 -3175 2572 -3123
rect 2504 -3196 2572 -3175
rect 2962 -563 3030 -542
rect 2962 -615 2970 -563
rect 3022 -615 3030 -563
rect 2962 -627 3030 -615
rect 2962 -679 2970 -627
rect 3022 -679 3030 -627
rect 2962 -691 3030 -679
rect 2962 -743 2970 -691
rect 3022 -743 3030 -691
rect 2962 -755 3030 -743
rect 2962 -807 2970 -755
rect 3022 -807 3030 -755
rect 2962 -819 3030 -807
rect 2962 -871 2970 -819
rect 3022 -871 3030 -819
rect 2962 -883 3030 -871
rect 2962 -935 2970 -883
rect 3022 -935 3030 -883
rect 2962 -947 3030 -935
rect 2962 -999 2970 -947
rect 3022 -999 3030 -947
rect 2962 -1011 3030 -999
rect 2962 -1063 2970 -1011
rect 3022 -1063 3030 -1011
rect 2962 -1075 3030 -1063
rect 2962 -1127 2970 -1075
rect 3022 -1127 3030 -1075
rect 2962 -1139 3030 -1127
rect 2962 -1191 2970 -1139
rect 3022 -1191 3030 -1139
rect 2962 -1203 3030 -1191
rect 2962 -1255 2970 -1203
rect 3022 -1255 3030 -1203
rect 2962 -1267 3030 -1255
rect 2962 -1319 2970 -1267
rect 3022 -1319 3030 -1267
rect 2962 -1331 3030 -1319
rect 2962 -1383 2970 -1331
rect 3022 -1383 3030 -1331
rect 2962 -1395 3030 -1383
rect 2962 -1447 2970 -1395
rect 3022 -1447 3030 -1395
rect 2962 -1459 3030 -1447
rect 2962 -1511 2970 -1459
rect 3022 -1511 3030 -1459
rect 2962 -1523 3030 -1511
rect 2962 -1575 2970 -1523
rect 3022 -1575 3030 -1523
rect 2962 -1587 3030 -1575
rect 2962 -1639 2970 -1587
rect 3022 -1639 3030 -1587
rect 2962 -1651 3030 -1639
rect 2962 -1703 2970 -1651
rect 3022 -1703 3030 -1651
rect 2962 -1715 3030 -1703
rect 2962 -1767 2970 -1715
rect 3022 -1767 3030 -1715
rect 2962 -1779 3030 -1767
rect 2962 -1831 2970 -1779
rect 3022 -1831 3030 -1779
rect 2962 -1843 3030 -1831
rect 2962 -1895 2970 -1843
rect 3022 -1895 3030 -1843
rect 2962 -1907 3030 -1895
rect 2962 -1959 2970 -1907
rect 3022 -1959 3030 -1907
rect 2962 -1971 3030 -1959
rect 2962 -2023 2970 -1971
rect 3022 -2023 3030 -1971
rect 2962 -2035 3030 -2023
rect 2962 -2087 2970 -2035
rect 3022 -2087 3030 -2035
rect 2962 -2099 3030 -2087
rect 2962 -2151 2970 -2099
rect 3022 -2151 3030 -2099
rect 2962 -2163 3030 -2151
rect 2962 -2215 2970 -2163
rect 3022 -2215 3030 -2163
rect 2962 -2227 3030 -2215
rect 2962 -2279 2970 -2227
rect 3022 -2279 3030 -2227
rect 2962 -2291 3030 -2279
rect 2962 -2343 2970 -2291
rect 3022 -2343 3030 -2291
rect 2962 -2355 3030 -2343
rect 2962 -2407 2970 -2355
rect 3022 -2407 3030 -2355
rect 2962 -2419 3030 -2407
rect 2962 -2471 2970 -2419
rect 3022 -2471 3030 -2419
rect 2962 -2483 3030 -2471
rect 2962 -2535 2970 -2483
rect 3022 -2535 3030 -2483
rect 2962 -2547 3030 -2535
rect 2962 -2599 2970 -2547
rect 3022 -2599 3030 -2547
rect 2962 -2611 3030 -2599
rect 2962 -2663 2970 -2611
rect 3022 -2663 3030 -2611
rect 2962 -2675 3030 -2663
rect 2962 -2727 2970 -2675
rect 3022 -2727 3030 -2675
rect 2962 -2739 3030 -2727
rect 2962 -2791 2970 -2739
rect 3022 -2791 3030 -2739
rect 2962 -2803 3030 -2791
rect 2962 -2855 2970 -2803
rect 3022 -2855 3030 -2803
rect 2962 -2867 3030 -2855
rect 2962 -2919 2970 -2867
rect 3022 -2919 3030 -2867
rect 2962 -2931 3030 -2919
rect 2962 -2983 2970 -2931
rect 3022 -2983 3030 -2931
rect 2962 -2995 3030 -2983
rect 2962 -3047 2970 -2995
rect 3022 -3047 3030 -2995
rect 2962 -3059 3030 -3047
rect 2962 -3111 2970 -3059
rect 3022 -3111 3030 -3059
rect 2962 -3123 3030 -3111
rect 2962 -3175 2970 -3123
rect 3022 -3175 3030 -3123
rect 2962 -3472 3030 -3175
rect 3420 -563 3488 -264
rect 3420 -615 3428 -563
rect 3480 -615 3488 -563
rect 3420 -627 3488 -615
rect 3420 -679 3428 -627
rect 3480 -679 3488 -627
rect 3420 -691 3488 -679
rect 3420 -743 3428 -691
rect 3480 -743 3488 -691
rect 3420 -755 3488 -743
rect 3420 -807 3428 -755
rect 3480 -807 3488 -755
rect 3420 -819 3488 -807
rect 3420 -871 3428 -819
rect 3480 -871 3488 -819
rect 3420 -883 3488 -871
rect 3420 -935 3428 -883
rect 3480 -935 3488 -883
rect 3420 -947 3488 -935
rect 3420 -999 3428 -947
rect 3480 -999 3488 -947
rect 3420 -1011 3488 -999
rect 3420 -1063 3428 -1011
rect 3480 -1063 3488 -1011
rect 3420 -1075 3488 -1063
rect 3420 -1127 3428 -1075
rect 3480 -1127 3488 -1075
rect 3420 -1139 3488 -1127
rect 3420 -1191 3428 -1139
rect 3480 -1191 3488 -1139
rect 3420 -1203 3488 -1191
rect 3420 -1255 3428 -1203
rect 3480 -1255 3488 -1203
rect 3420 -1267 3488 -1255
rect 3420 -1319 3428 -1267
rect 3480 -1319 3488 -1267
rect 3420 -1331 3488 -1319
rect 3420 -1383 3428 -1331
rect 3480 -1383 3488 -1331
rect 3420 -1395 3488 -1383
rect 3420 -1447 3428 -1395
rect 3480 -1447 3488 -1395
rect 3420 -1459 3488 -1447
rect 3420 -1511 3428 -1459
rect 3480 -1511 3488 -1459
rect 3420 -1523 3488 -1511
rect 3420 -1575 3428 -1523
rect 3480 -1575 3488 -1523
rect 3420 -1587 3488 -1575
rect 3420 -1639 3428 -1587
rect 3480 -1639 3488 -1587
rect 3420 -1651 3488 -1639
rect 3420 -1703 3428 -1651
rect 3480 -1703 3488 -1651
rect 3420 -1715 3488 -1703
rect 3420 -1767 3428 -1715
rect 3480 -1767 3488 -1715
rect 3420 -1779 3488 -1767
rect 3420 -1831 3428 -1779
rect 3480 -1831 3488 -1779
rect 3420 -1843 3488 -1831
rect 3420 -1895 3428 -1843
rect 3480 -1895 3488 -1843
rect 3420 -1907 3488 -1895
rect 3420 -1959 3428 -1907
rect 3480 -1959 3488 -1907
rect 3420 -1971 3488 -1959
rect 3420 -2023 3428 -1971
rect 3480 -2023 3488 -1971
rect 3420 -2035 3488 -2023
rect 3420 -2087 3428 -2035
rect 3480 -2087 3488 -2035
rect 3420 -2099 3488 -2087
rect 3420 -2151 3428 -2099
rect 3480 -2151 3488 -2099
rect 3420 -2163 3488 -2151
rect 3420 -2215 3428 -2163
rect 3480 -2215 3488 -2163
rect 3420 -2227 3488 -2215
rect 3420 -2279 3428 -2227
rect 3480 -2279 3488 -2227
rect 3420 -2291 3488 -2279
rect 3420 -2343 3428 -2291
rect 3480 -2343 3488 -2291
rect 3420 -2355 3488 -2343
rect 3420 -2407 3428 -2355
rect 3480 -2407 3488 -2355
rect 3420 -2419 3488 -2407
rect 3420 -2471 3428 -2419
rect 3480 -2471 3488 -2419
rect 3420 -2483 3488 -2471
rect 3420 -2535 3428 -2483
rect 3480 -2535 3488 -2483
rect 3420 -2547 3488 -2535
rect 3420 -2599 3428 -2547
rect 3480 -2599 3488 -2547
rect 3420 -2611 3488 -2599
rect 3420 -2663 3428 -2611
rect 3480 -2663 3488 -2611
rect 3420 -2675 3488 -2663
rect 3420 -2727 3428 -2675
rect 3480 -2727 3488 -2675
rect 3420 -2739 3488 -2727
rect 3420 -2791 3428 -2739
rect 3480 -2791 3488 -2739
rect 3420 -2803 3488 -2791
rect 3420 -2855 3428 -2803
rect 3480 -2855 3488 -2803
rect 3420 -2867 3488 -2855
rect 3420 -2919 3428 -2867
rect 3480 -2919 3488 -2867
rect 3420 -2931 3488 -2919
rect 3420 -2983 3428 -2931
rect 3480 -2983 3488 -2931
rect 3420 -2995 3488 -2983
rect 3420 -3047 3428 -2995
rect 3480 -3047 3488 -2995
rect 3420 -3059 3488 -3047
rect 3420 -3111 3428 -3059
rect 3480 -3111 3488 -3059
rect 3420 -3123 3488 -3111
rect 3420 -3175 3428 -3123
rect 3480 -3175 3488 -3123
rect 3420 -3196 3488 -3175
rect -702 -3676 3030 -3472
<< via2 >>
rect 849 2712 905 2714
rect 849 2660 851 2712
rect 851 2660 903 2712
rect 903 2660 905 2712
rect 849 2658 905 2660
rect 1651 2712 1707 2714
rect 1651 2660 1653 2712
rect 1653 2660 1705 2712
rect 1705 2660 1707 2712
rect 1651 2658 1707 2660
rect 831 2083 887 2085
rect 831 2031 833 2083
rect 833 2031 885 2083
rect 885 2031 887 2083
rect 831 2029 887 2031
rect 1039 1869 1095 1925
rect 711 1243 767 1245
rect 711 1191 713 1243
rect 713 1191 765 1243
rect 765 1191 767 1243
rect 711 1189 767 1191
rect 715 1099 771 1101
rect 715 1047 717 1099
rect 717 1047 769 1099
rect 769 1047 771 1099
rect 715 1045 771 1047
rect 1553 1233 1609 1235
rect 1553 1181 1555 1233
rect 1555 1181 1607 1233
rect 1607 1181 1609 1233
rect 1553 1179 1609 1181
rect 1551 1103 1607 1105
rect 1551 1051 1553 1103
rect 1553 1051 1605 1103
rect 1605 1051 1607 1103
rect 1551 1049 1607 1051
rect 1043 297 1099 299
rect 1043 245 1045 297
rect 1045 245 1097 297
rect 1097 245 1099 297
rect 1043 243 1099 245
rect 1211 299 1267 301
rect 1211 247 1213 299
rect 1213 247 1265 299
rect 1265 247 1267 299
rect 1211 245 1267 247
rect -1104 -216 3432 0
<< metal3 >>
rect -1404 2714 3964 2730
rect -1404 2658 849 2714
rect 905 2658 1651 2714
rect 1707 2658 3964 2714
rect -1404 2644 3964 2658
rect 818 2085 898 2096
rect 818 2029 831 2085
rect 887 2082 898 2085
rect 887 2029 1256 2082
rect 818 2016 1256 2029
rect 1016 1925 1120 1950
rect 1016 1869 1039 1925
rect 1095 1869 1120 1925
rect 1016 1852 1120 1869
rect 650 1245 826 1298
rect 650 1189 711 1245
rect 767 1189 826 1245
rect 650 1174 826 1189
rect 650 1110 706 1174
rect 770 1110 826 1174
rect 650 1101 826 1110
rect 650 1045 715 1101
rect 771 1045 826 1101
rect 650 1002 826 1045
rect 1056 324 1120 1852
rect 1020 299 1120 324
rect 1020 243 1043 299
rect 1099 243 1120 299
rect 1020 226 1120 243
rect 1192 324 1256 2016
rect 1494 1235 1670 1298
rect 1494 1179 1553 1235
rect 1609 1179 1670 1235
rect 1494 1174 1670 1179
rect 1494 1110 1548 1174
rect 1612 1110 1670 1174
rect 1494 1105 1670 1110
rect 1494 1049 1551 1105
rect 1607 1049 1670 1105
rect 1494 1002 1670 1049
rect 1192 301 1292 324
rect 1192 245 1211 301
rect 1267 245 1292 301
rect 1192 226 1292 245
rect -1158 4 3486 36
rect -1158 -220 -1148 4
rect 3476 -220 3486 4
rect -1158 -252 3486 -220
<< via3 >>
rect 706 1110 770 1174
rect 1548 1110 1612 1174
rect -1148 0 3476 4
rect -1148 -216 -1104 0
rect -1104 -216 3432 0
rect 3432 -216 3476 0
rect -1148 -220 3476 -216
<< metal4 >>
rect 650 1266 1670 1298
rect 650 1174 1040 1266
rect 650 1110 706 1174
rect 770 1110 1040 1174
rect 650 1030 1040 1110
rect 1276 1174 1670 1266
rect 1276 1110 1548 1174
rect 1612 1110 1670 1174
rect 1276 1030 1670 1110
rect 650 1002 1670 1030
rect -1154 10 3482 42
rect -1154 4 -1034 10
rect -798 4 -714 10
rect -478 4 -394 10
rect -158 4 -74 10
rect 162 4 246 10
rect 482 4 566 10
rect 802 4 886 10
rect 1122 4 1206 10
rect 1442 4 1526 10
rect 1762 4 1846 10
rect 2082 4 2166 10
rect 2402 4 2486 10
rect 2722 4 2806 10
rect 3042 4 3126 10
rect 3362 4 3482 10
rect -1154 -220 -1148 4
rect 3476 -220 3482 4
rect -1154 -226 -1034 -220
rect -798 -226 -714 -220
rect -478 -226 -394 -220
rect -158 -226 -74 -220
rect 162 -226 246 -220
rect 482 -226 566 -220
rect 802 -226 886 -220
rect 1122 -226 1206 -220
rect 1442 -226 1526 -220
rect 1762 -226 1846 -220
rect 2082 -226 2166 -220
rect 2402 -226 2486 -220
rect 2722 -226 2806 -220
rect 3042 -226 3126 -220
rect 3362 -226 3482 -220
rect -1154 -258 3482 -226
<< via4 >>
rect 1040 1030 1276 1266
rect -1034 4 -798 10
rect -714 4 -478 10
rect -394 4 -158 10
rect -74 4 162 10
rect 246 4 482 10
rect 566 4 802 10
rect 886 4 1122 10
rect 1206 4 1442 10
rect 1526 4 1762 10
rect 1846 4 2082 10
rect 2166 4 2402 10
rect 2486 4 2722 10
rect 2806 4 3042 10
rect 3126 4 3362 10
rect -1034 -220 -798 4
rect -714 -220 -478 4
rect -394 -220 -158 4
rect -74 -220 162 4
rect 246 -220 482 4
rect 566 -220 802 4
rect 886 -220 1122 4
rect 1206 -220 1442 4
rect 1526 -220 1762 4
rect 1846 -220 2082 4
rect 2166 -220 2402 4
rect 2486 -220 2722 4
rect 2806 -220 3042 4
rect 3126 -220 3362 4
rect -1034 -226 -798 -220
rect -714 -226 -478 -220
rect -394 -226 -158 -220
rect -74 -226 162 -220
rect 246 -226 482 -220
rect 566 -226 802 -220
rect 886 -226 1122 -220
rect 1206 -226 1442 -220
rect 1526 -226 1762 -220
rect 1846 -226 2082 -220
rect 2166 -226 2402 -220
rect 2486 -226 2722 -220
rect 2806 -226 3042 -220
rect 3126 -226 3362 -220
<< metal5 >>
rect 990 1266 1330 1298
rect 990 1030 1040 1266
rect 1276 1030 1330 1266
rect 990 66 1330 1030
rect -1178 10 3506 66
rect -1178 -226 -1034 10
rect -798 -226 -714 10
rect -478 -226 -394 10
rect -158 -226 -74 10
rect 162 -226 246 10
rect 482 -226 566 10
rect 802 -226 886 10
rect 1122 -226 1206 10
rect 1442 -226 1526 10
rect 1762 -226 1846 10
rect 2082 -226 2166 10
rect 2402 -226 2486 10
rect 2722 -226 2806 10
rect 3042 -226 3126 10
rect 3362 -226 3506 10
rect -1178 -282 3506 -226
use sky130_fd_pr__nfet_01v8_lvt_MGW8MS  sky130_fd_pr__nfet_01v8_lvt_MGW8MS_0
timestamp 1611881054
transform 1 0 509 0 1 616
box -611 -224 611 224
use sky130_fd_pr__nfet_01v8_lvt_AV5GXG  sky130_fd_pr__nfet_01v8_lvt_AV5GXG_0
timestamp 1611881054
transform 1 0 1164 0 1 -1869
box -2421 -1500 2421 1494
use sky130_fd_pr__pfet_01v8_lvt_TGGFET  sky130_fd_pr__pfet_01v8_lvt_TGGFET_0
timestamp 1611881054
transform -1 0 -22 0 -1 5591
box -1312 -1019 1312 1019
use sky130_fd_pr__pfet_01v8_lvt_TGGFET  sky130_fd_pr__pfet_01v8_lvt_TGGFET_1
timestamp 1611881054
transform 1 0 2602 0 -1 5591
box -1312 -1019 1312 1019
use sky130_fd_pr__pfet_01v8_lvt_TGGFET  sky130_fd_pr__pfet_01v8_lvt_TGGFET_2
timestamp 1611881054
transform 1 0 2602 0 1 3553
box -1312 -1019 1312 1019
use sky130_fd_pr__pfet_01v8_lvt_TGGFET  sky130_fd_pr__pfet_01v8_lvt_TGGFET_3
timestamp 1611881054
transform -1 0 -22 0 1 3553
box -1312 -1019 1312 1019
<< end >>
