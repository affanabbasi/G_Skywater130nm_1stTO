magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect -296 -819 296 819
<< pmoslvt >>
rect -100 -600 100 600
<< pdiff >>
rect -158 561 -100 600
rect -158 527 -146 561
rect -112 527 -100 561
rect -158 493 -100 527
rect -158 459 -146 493
rect -112 459 -100 493
rect -158 425 -100 459
rect -158 391 -146 425
rect -112 391 -100 425
rect -158 357 -100 391
rect -158 323 -146 357
rect -112 323 -100 357
rect -158 289 -100 323
rect -158 255 -146 289
rect -112 255 -100 289
rect -158 221 -100 255
rect -158 187 -146 221
rect -112 187 -100 221
rect -158 153 -100 187
rect -158 119 -146 153
rect -112 119 -100 153
rect -158 85 -100 119
rect -158 51 -146 85
rect -112 51 -100 85
rect -158 17 -100 51
rect -158 -17 -146 17
rect -112 -17 -100 17
rect -158 -51 -100 -17
rect -158 -85 -146 -51
rect -112 -85 -100 -51
rect -158 -119 -100 -85
rect -158 -153 -146 -119
rect -112 -153 -100 -119
rect -158 -187 -100 -153
rect -158 -221 -146 -187
rect -112 -221 -100 -187
rect -158 -255 -100 -221
rect -158 -289 -146 -255
rect -112 -289 -100 -255
rect -158 -323 -100 -289
rect -158 -357 -146 -323
rect -112 -357 -100 -323
rect -158 -391 -100 -357
rect -158 -425 -146 -391
rect -112 -425 -100 -391
rect -158 -459 -100 -425
rect -158 -493 -146 -459
rect -112 -493 -100 -459
rect -158 -527 -100 -493
rect -158 -561 -146 -527
rect -112 -561 -100 -527
rect -158 -600 -100 -561
rect 100 561 158 600
rect 100 527 112 561
rect 146 527 158 561
rect 100 493 158 527
rect 100 459 112 493
rect 146 459 158 493
rect 100 425 158 459
rect 100 391 112 425
rect 146 391 158 425
rect 100 357 158 391
rect 100 323 112 357
rect 146 323 158 357
rect 100 289 158 323
rect 100 255 112 289
rect 146 255 158 289
rect 100 221 158 255
rect 100 187 112 221
rect 146 187 158 221
rect 100 153 158 187
rect 100 119 112 153
rect 146 119 158 153
rect 100 85 158 119
rect 100 51 112 85
rect 146 51 158 85
rect 100 17 158 51
rect 100 -17 112 17
rect 146 -17 158 17
rect 100 -51 158 -17
rect 100 -85 112 -51
rect 146 -85 158 -51
rect 100 -119 158 -85
rect 100 -153 112 -119
rect 146 -153 158 -119
rect 100 -187 158 -153
rect 100 -221 112 -187
rect 146 -221 158 -187
rect 100 -255 158 -221
rect 100 -289 112 -255
rect 146 -289 158 -255
rect 100 -323 158 -289
rect 100 -357 112 -323
rect 146 -357 158 -323
rect 100 -391 158 -357
rect 100 -425 112 -391
rect 146 -425 158 -391
rect 100 -459 158 -425
rect 100 -493 112 -459
rect 146 -493 158 -459
rect 100 -527 158 -493
rect 100 -561 112 -527
rect 146 -561 158 -527
rect 100 -600 158 -561
<< pdiffc >>
rect -146 527 -112 561
rect -146 459 -112 493
rect -146 391 -112 425
rect -146 323 -112 357
rect -146 255 -112 289
rect -146 187 -112 221
rect -146 119 -112 153
rect -146 51 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -51
rect -146 -153 -112 -119
rect -146 -221 -112 -187
rect -146 -289 -112 -255
rect -146 -357 -112 -323
rect -146 -425 -112 -391
rect -146 -493 -112 -459
rect -146 -561 -112 -527
rect 112 527 146 561
rect 112 459 146 493
rect 112 391 146 425
rect 112 323 146 357
rect 112 255 146 289
rect 112 187 146 221
rect 112 119 146 153
rect 112 51 146 85
rect 112 -17 146 17
rect 112 -85 146 -51
rect 112 -153 146 -119
rect 112 -221 146 -187
rect 112 -289 146 -255
rect 112 -357 146 -323
rect 112 -425 146 -391
rect 112 -493 146 -459
rect 112 -561 146 -527
<< nsubdiff >>
rect -260 749 -153 783
rect -119 749 -85 783
rect -51 749 -17 783
rect 17 749 51 783
rect 85 749 119 783
rect 153 749 260 783
rect -260 663 -226 749
rect -260 595 -226 629
rect 226 663 260 749
rect -260 527 -226 561
rect -260 459 -226 493
rect -260 391 -226 425
rect -260 323 -226 357
rect -260 255 -226 289
rect -260 187 -226 221
rect -260 119 -226 153
rect -260 51 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect -260 -153 -226 -119
rect -260 -221 -226 -187
rect -260 -289 -226 -255
rect -260 -357 -226 -323
rect -260 -425 -226 -391
rect -260 -493 -226 -459
rect -260 -561 -226 -527
rect -260 -629 -226 -595
rect 226 595 260 629
rect 226 527 260 561
rect 226 459 260 493
rect 226 391 260 425
rect 226 323 260 357
rect 226 255 260 289
rect 226 187 260 221
rect 226 119 260 153
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -153 260 -119
rect 226 -221 260 -187
rect 226 -289 260 -255
rect 226 -357 260 -323
rect 226 -425 260 -391
rect 226 -493 260 -459
rect 226 -561 260 -527
rect -260 -749 -226 -663
rect 226 -629 260 -595
rect 226 -749 260 -663
rect -260 -783 -153 -749
rect -119 -783 -85 -749
rect -51 -783 -17 -749
rect 17 -783 51 -749
rect 85 -783 119 -749
rect 153 -783 260 -749
<< nsubdiffcont >>
rect -153 749 -119 783
rect -85 749 -51 783
rect -17 749 17 783
rect 51 749 85 783
rect 119 749 153 783
rect -260 629 -226 663
rect 226 629 260 663
rect -260 561 -226 595
rect -260 493 -226 527
rect -260 425 -226 459
rect -260 357 -226 391
rect -260 289 -226 323
rect -260 221 -226 255
rect -260 153 -226 187
rect -260 85 -226 119
rect -260 17 -226 51
rect -260 -51 -226 -17
rect -260 -119 -226 -85
rect -260 -187 -226 -153
rect -260 -255 -226 -221
rect -260 -323 -226 -289
rect -260 -391 -226 -357
rect -260 -459 -226 -425
rect -260 -527 -226 -493
rect -260 -595 -226 -561
rect 226 561 260 595
rect 226 493 260 527
rect 226 425 260 459
rect 226 357 260 391
rect 226 289 260 323
rect 226 221 260 255
rect 226 153 260 187
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect 226 -119 260 -85
rect 226 -187 260 -153
rect 226 -255 260 -221
rect 226 -323 260 -289
rect 226 -391 260 -357
rect 226 -459 260 -425
rect 226 -527 260 -493
rect 226 -595 260 -561
rect -260 -663 -226 -629
rect 226 -663 260 -629
rect -153 -783 -119 -749
rect -85 -783 -51 -749
rect -17 -783 17 -749
rect 51 -783 85 -749
rect 119 -783 153 -749
<< poly >>
rect -100 681 100 697
rect -100 647 -51 681
rect -17 647 17 681
rect 51 647 100 681
rect -100 600 100 647
rect -100 -647 100 -600
rect -100 -681 -51 -647
rect -17 -681 17 -647
rect 51 -681 100 -647
rect -100 -697 100 -681
<< polycont >>
rect -51 647 -17 681
rect 17 647 51 681
rect -51 -681 -17 -647
rect 17 -681 51 -647
<< locali >>
rect -260 749 -153 783
rect -119 749 -85 783
rect -51 749 -17 783
rect 17 749 51 783
rect 85 749 119 783
rect 153 749 260 783
rect -260 663 -226 749
rect -100 647 -51 681
rect -17 647 17 681
rect 51 647 100 681
rect 226 663 260 749
rect -260 595 -226 629
rect -260 527 -226 561
rect -260 459 -226 493
rect -260 391 -226 425
rect -260 323 -226 357
rect -260 255 -226 289
rect -260 187 -226 221
rect -260 119 -226 153
rect -260 51 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect -260 -153 -226 -119
rect -260 -221 -226 -187
rect -260 -289 -226 -255
rect -260 -357 -226 -323
rect -260 -425 -226 -391
rect -260 -493 -226 -459
rect -260 -561 -226 -527
rect -260 -629 -226 -595
rect -146 561 -112 604
rect -146 493 -112 527
rect -146 425 -112 459
rect -146 357 -112 391
rect -146 289 -112 323
rect -146 221 -112 255
rect -146 153 -112 187
rect -146 85 -112 119
rect -146 17 -112 51
rect -146 -51 -112 -17
rect -146 -119 -112 -85
rect -146 -187 -112 -153
rect -146 -255 -112 -221
rect -146 -323 -112 -289
rect -146 -391 -112 -357
rect -146 -459 -112 -425
rect -146 -527 -112 -493
rect -146 -604 -112 -561
rect 112 561 146 604
rect 112 493 146 527
rect 112 425 146 459
rect 112 357 146 391
rect 112 289 146 323
rect 112 221 146 255
rect 112 153 146 187
rect 112 85 146 119
rect 112 17 146 51
rect 112 -51 146 -17
rect 112 -119 146 -85
rect 112 -187 146 -153
rect 112 -255 146 -221
rect 112 -323 146 -289
rect 112 -391 146 -357
rect 112 -459 146 -425
rect 112 -527 146 -493
rect 112 -604 146 -561
rect 226 595 260 629
rect 226 527 260 561
rect 226 459 260 493
rect 226 391 260 425
rect 226 323 260 357
rect 226 255 260 289
rect 226 187 260 221
rect 226 119 260 153
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -153 260 -119
rect 226 -221 260 -187
rect 226 -289 260 -255
rect 226 -357 260 -323
rect 226 -425 260 -391
rect 226 -493 260 -459
rect 226 -561 260 -527
rect 226 -629 260 -595
rect -260 -749 -226 -663
rect -100 -681 -51 -647
rect -17 -681 17 -647
rect 51 -681 100 -647
rect 226 -749 260 -663
rect -260 -783 -153 -749
rect -119 -783 -85 -749
rect -51 -783 -17 -749
rect 17 -783 51 -749
rect 85 -783 119 -749
rect 153 -783 260 -749
<< properties >>
string FIXED_BBOX -243 -766 243 766
<< end >>
