magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< error_s >>
rect -46 4706 1258 4758
rect -46 4658 6 4706
rect 26 4658 1186 4686
rect 54 4606 1186 4658
rect 54 3606 106 4606
rect 1106 3606 1186 4606
rect 54 3554 1186 3606
rect 1158 3526 1186 3554
rect 1206 3506 1258 4706
rect 1158 3454 1258 3506
rect 48 3040 1352 3092
rect 48 2992 100 3040
rect 120 2992 1280 3020
rect 148 2940 1280 2992
rect 148 1940 200 2940
rect 1200 1940 1280 2940
rect 148 1888 1280 1940
rect 1252 1860 1280 1888
rect 1300 1840 1352 3040
rect 1252 1788 1352 1840
<< nwell >>
rect 15068 3088 18654 3102
rect 15062 2808 18654 3088
rect 15062 2794 18648 2808
<< locali >>
rect 7244 2850 7320 2914
rect 7842 2864 7922 2914
rect 17426 2750 17466 2752
rect 16542 2729 16576 2730
rect 15740 2713 15774 2714
rect 15648 2711 15682 2712
rect 17426 2716 17429 2750
rect 17463 2716 17466 2750
rect 17426 2714 17466 2716
rect 16542 2694 16576 2695
rect 15740 2678 15774 2679
rect 15648 2676 15682 2677
rect 18546 2634 18584 2638
rect 16634 2632 16674 2634
rect 16634 2598 16637 2632
rect 16671 2598 16674 2632
rect 16634 2596 16674 2598
rect 17516 2632 17556 2634
rect 17516 2598 17519 2632
rect 17553 2598 17556 2632
rect 17516 2596 17556 2598
rect 18546 2600 18548 2634
rect 18582 2600 18584 2634
rect 18546 2596 18584 2600
rect 12064 2446 12098 2450
rect 12064 2433 12118 2446
rect 12064 2399 12072 2433
rect 12106 2399 12118 2433
rect 12064 2380 12118 2399
rect 12796 2398 12799 2432
rect 12833 2398 12836 2432
rect 12064 2376 12098 2380
rect 11148 1528 11184 1540
rect 11148 1494 11149 1528
rect 11183 1494 11184 1528
rect 11148 1482 11184 1494
rect 11234 1370 11241 1404
rect 11275 1370 11313 1404
rect 11347 1370 11385 1404
rect 11419 1370 11457 1404
rect 11491 1370 11529 1404
rect 11563 1370 11601 1404
rect 11635 1370 11673 1404
rect 11707 1370 11745 1404
rect 11779 1370 11817 1404
rect 11851 1370 11889 1404
rect 11923 1370 11961 1404
rect 11995 1370 12033 1404
rect 12067 1370 12105 1404
rect 12139 1370 12177 1404
rect 12211 1370 12249 1404
rect 12283 1370 12321 1404
rect 12355 1370 12393 1404
rect 12427 1370 12465 1404
rect 12499 1370 12537 1404
rect 12571 1370 12609 1404
rect 12643 1370 12681 1404
rect 12715 1370 12753 1404
rect 12787 1370 12825 1404
rect 12859 1370 12897 1404
rect 12931 1370 12969 1404
rect 13003 1370 13041 1404
rect 13075 1370 13113 1404
rect 13147 1370 13185 1404
rect 13219 1370 13257 1404
rect 13291 1370 13329 1404
rect 13363 1370 13401 1404
rect 13435 1370 13473 1404
rect 13507 1370 13545 1404
rect 13579 1370 13617 1404
rect 13651 1370 13689 1404
rect 13723 1370 13730 1404
rect 4798 90 4829 124
rect 4863 90 4901 124
rect 4935 90 4973 124
rect 5007 90 5045 124
rect 5079 90 5117 124
rect 5151 90 5189 124
rect 5223 90 5254 124
rect 1934 36 1965 70
rect 1999 36 2037 70
rect 2071 36 2109 70
rect 2143 36 2181 70
rect 2215 36 2253 70
rect 2287 36 2325 70
rect 2359 36 2390 70
<< viali >>
rect 15648 2677 15682 2711
rect 15740 2679 15774 2713
rect 16542 2695 16576 2729
rect 17429 2716 17463 2750
rect 18452 2726 18486 2760
rect 16637 2598 16671 2632
rect 17519 2598 17553 2632
rect 18548 2600 18582 2634
rect 12072 2399 12106 2433
rect 12799 2398 12833 2432
rect 11149 1494 11183 1528
rect 11241 1370 11275 1404
rect 11313 1370 11347 1404
rect 11385 1370 11419 1404
rect 11457 1370 11491 1404
rect 11529 1370 11563 1404
rect 11601 1370 11635 1404
rect 11673 1370 11707 1404
rect 11745 1370 11779 1404
rect 11817 1370 11851 1404
rect 11889 1370 11923 1404
rect 11961 1370 11995 1404
rect 12033 1370 12067 1404
rect 12105 1370 12139 1404
rect 12177 1370 12211 1404
rect 12249 1370 12283 1404
rect 12321 1370 12355 1404
rect 12393 1370 12427 1404
rect 12465 1370 12499 1404
rect 12537 1370 12571 1404
rect 12609 1370 12643 1404
rect 12681 1370 12715 1404
rect 12753 1370 12787 1404
rect 12825 1370 12859 1404
rect 12897 1370 12931 1404
rect 12969 1370 13003 1404
rect 13041 1370 13075 1404
rect 13113 1370 13147 1404
rect 13185 1370 13219 1404
rect 13257 1370 13291 1404
rect 13329 1370 13363 1404
rect 13401 1370 13435 1404
rect 13473 1370 13507 1404
rect 13545 1370 13579 1404
rect 13617 1370 13651 1404
rect 13689 1370 13723 1404
rect 4829 90 4863 124
rect 4901 90 4935 124
rect 4973 90 5007 124
rect 5045 90 5079 124
rect 5117 90 5151 124
rect 5189 90 5223 124
rect 1965 36 1999 70
rect 2037 36 2071 70
rect 2109 36 2143 70
rect 2181 36 2215 70
rect 2253 36 2287 70
rect 2325 36 2359 70
<< metal1 >>
rect -1515 5650 -424 5918
rect 2973 5672 18824 5872
rect -1515 5150 -1280 5650
rect -652 5150 -424 5650
rect 2962 5618 18824 5672
rect 4184 5528 18824 5618
rect 4184 5522 16971 5528
rect 5970 5426 16971 5522
rect 6051 5328 16971 5426
rect 6051 5280 9232 5328
rect 9136 5272 9232 5280
rect 9304 5280 16971 5328
rect 9304 5272 9802 5280
rect -1515 4860 -424 5150
rect 15558 5028 16971 5280
rect 17599 5028 18824 5528
rect 7930 4802 8014 4826
rect 7930 4750 7946 4802
rect 7998 4750 8014 4802
rect 7930 4726 8014 4750
rect 9448 4812 9558 4850
rect 9448 4760 9480 4812
rect 9532 4760 9558 4812
rect 7242 4676 7336 4680
rect 7242 4624 7263 4676
rect 7315 4624 7336 4676
rect 7242 4612 7336 4624
rect 7242 4560 7263 4612
rect 7315 4560 7336 4612
rect 7242 4556 7336 4560
rect -1515 4244 -424 4512
rect -1515 3744 -1280 4244
rect -652 3744 -424 4244
rect 9448 4264 9558 4760
rect 11498 4264 11596 4272
rect 9448 4180 11600 4264
rect 9454 4174 11600 4180
rect -1515 3454 -424 3744
rect 7746 3034 7806 3048
rect 7096 3023 7148 3028
rect 7096 2966 7148 2971
rect 7746 2982 7750 3034
rect 7802 2982 7806 3034
rect 7746 2968 7806 2982
rect 8110 3027 8162 3042
rect 8110 2960 8162 2975
rect 7254 2914 7316 2916
rect 7244 2906 7320 2914
rect 6920 2900 7324 2906
rect -1515 2585 -424 2853
rect 6920 2848 6935 2900
rect 6987 2848 7324 2900
rect 6920 2842 7324 2848
rect 7842 2904 7918 2912
rect 7842 2870 7866 2904
rect 7900 2870 7918 2904
rect 6886 2738 6980 2742
rect 6886 2686 6910 2738
rect 6962 2726 6980 2738
rect 7842 2726 7918 2870
rect 11498 2792 11596 4174
rect 15558 3029 18824 5028
rect 18996 3156 20087 3424
rect 15558 2952 15732 3029
rect 15828 2948 16478 3029
rect 16708 3008 18766 3029
rect 16708 3004 18672 3008
rect 6962 2686 7920 2726
rect 11498 2713 11634 2792
rect 17514 2762 18498 2774
rect 17452 2760 18498 2762
rect 16630 2750 18452 2760
rect 16630 2742 17429 2750
rect 15726 2729 17429 2742
rect 6886 2684 7920 2686
rect 6886 2668 6980 2684
rect 9228 2669 9378 2702
rect -1515 2085 -1280 2585
rect -652 2085 -424 2585
rect 9228 2617 9278 2669
rect 9330 2617 9378 2669
rect 11498 2661 11539 2713
rect 11591 2661 11634 2713
rect 11498 2652 11634 2661
rect 12608 2720 15200 2722
rect 12608 2711 15696 2720
rect 12608 2677 15648 2711
rect 15682 2677 15696 2711
rect 12608 2656 15696 2677
rect 15726 2713 16542 2729
rect 15726 2679 15740 2713
rect 15774 2695 16542 2713
rect 16576 2716 17429 2729
rect 17463 2726 18452 2750
rect 18486 2726 18498 2760
rect 17463 2716 18498 2726
rect 16576 2706 18498 2716
rect 16576 2695 17614 2706
rect 15774 2694 17614 2695
rect 15774 2688 17482 2694
rect 15774 2679 16844 2688
rect 15726 2678 16844 2679
rect 15726 2670 16598 2678
rect 18996 2658 19231 3156
rect 18712 2656 19231 2658
rect 19859 2656 20087 3156
rect 11504 2626 11634 2652
rect 18712 2650 20087 2656
rect 17510 2644 20087 2650
rect 16614 2634 20087 2644
rect 16614 2632 18548 2634
rect 9228 2448 9378 2617
rect 16614 2598 16637 2632
rect 16671 2613 17519 2632
rect 16671 2598 17280 2613
rect 16614 2582 17280 2598
rect 17354 2598 17519 2613
rect 17553 2617 18548 2632
rect 17553 2598 17629 2617
rect 17354 2586 17629 2598
rect 17703 2600 18548 2617
rect 18582 2625 20087 2634
rect 18582 2621 18824 2625
rect 18582 2600 18656 2621
rect 17703 2586 18656 2600
rect 18732 2586 18824 2621
rect 18898 2586 20087 2625
rect 17354 2582 17560 2586
rect 18644 2518 18754 2546
rect 15834 2485 16484 2518
rect 16696 2485 18754 2518
rect 11792 2448 12114 2452
rect 12980 2448 13090 2450
rect 9222 2433 12114 2448
rect 9222 2399 12072 2433
rect 12106 2399 12114 2433
rect 9222 2378 12114 2399
rect 12790 2432 13090 2448
rect 15658 2436 18824 2485
rect 12790 2398 12799 2432
rect 12833 2398 13090 2432
rect 12790 2378 13090 2398
rect 9222 2376 11806 2378
rect -1515 1795 -424 2085
rect 4478 1930 4582 2352
rect 7580 2146 7692 2176
rect 7580 2094 7610 2146
rect 7662 2094 7692 2146
rect 7580 2064 7692 2094
rect 12980 2125 13090 2378
rect 12980 2073 13004 2125
rect 13056 2073 13090 2125
rect 12980 2042 13090 2073
rect 5408 1930 7474 1958
rect 4478 1788 7474 1930
rect 9004 1883 9090 1896
rect 9004 1831 9021 1883
rect 9073 1831 9090 1883
rect 9004 1818 9090 1831
rect 5408 1253 7474 1788
rect 7562 1576 7714 1652
rect 7562 1524 7610 1576
rect 7662 1566 7714 1576
rect 7662 1528 11208 1566
rect 7662 1524 11149 1528
rect 7562 1494 11149 1524
rect 11183 1494 11208 1528
rect 7562 1474 11208 1494
rect 7562 1470 7714 1474
rect 11218 1404 13744 1416
rect 11218 1370 11241 1404
rect 11275 1370 11313 1404
rect 11347 1370 11385 1404
rect 11419 1370 11457 1404
rect 11491 1370 11529 1404
rect 11563 1370 11601 1404
rect 11635 1370 11673 1404
rect 11707 1370 11745 1404
rect 11779 1370 11817 1404
rect 11851 1370 11889 1404
rect 11923 1370 11961 1404
rect 11995 1370 12033 1404
rect 12067 1370 12105 1404
rect 12139 1370 12177 1404
rect 12211 1370 12249 1404
rect 12283 1370 12321 1404
rect 12355 1370 12393 1404
rect 12427 1370 12465 1404
rect 12499 1370 12537 1404
rect 12571 1370 12609 1404
rect 12643 1370 12681 1404
rect 12715 1370 12753 1404
rect 12787 1370 12825 1404
rect 12859 1370 12897 1404
rect 12931 1370 12969 1404
rect 13003 1370 13041 1404
rect 13075 1370 13113 1404
rect 13147 1370 13185 1404
rect 13219 1370 13257 1404
rect 13291 1370 13329 1404
rect 13363 1370 13401 1404
rect 13435 1370 13473 1404
rect 13507 1370 13545 1404
rect 13579 1370 13617 1404
rect 13651 1370 13689 1404
rect 13723 1370 13744 1404
rect 11218 1292 13744 1370
rect 15576 1322 18824 2436
rect 18996 2366 20087 2586
rect 4768 124 5294 135
rect 4768 90 4829 124
rect 4863 90 4901 124
rect 4935 90 4973 124
rect 5007 90 5045 124
rect 5079 90 5117 124
rect 5151 90 5189 124
rect 5223 90 5294 124
rect 1908 74 2403 89
rect 4768 74 5294 90
rect 5408 74 6519 1253
rect 10978 1251 11064 1264
rect 14068 1260 18824 1322
rect 10978 1199 10995 1251
rect 11047 1199 11064 1251
rect 10978 1186 11064 1199
rect 14057 1183 18824 1260
rect 1802 70 6519 74
rect 1802 36 1965 70
rect 1999 36 2037 70
rect 2071 36 2109 70
rect 2143 36 2181 70
rect 2215 36 2253 70
rect 2287 36 2325 70
rect 2359 36 6519 70
rect 1802 16 6519 36
rect 7196 806 8287 1074
rect 7196 306 7431 806
rect 8059 306 8287 806
rect 7196 16 8287 306
rect 8908 854 18824 1183
rect 8908 354 16899 854
rect 17527 354 18824 854
rect 8908 16 18824 354
<< via1 >>
rect -1280 5150 -652 5650
rect 16971 5028 17599 5528
rect 7946 4750 7998 4802
rect 9480 4760 9532 4812
rect 7263 4624 7315 4676
rect 7263 4560 7315 4612
rect -1280 3744 -652 4244
rect 7096 2971 7148 3023
rect 7750 2982 7802 3034
rect 8110 2975 8162 3027
rect 6935 2848 6987 2900
rect 6910 2686 6962 2738
rect -1280 2085 -652 2585
rect 9278 2617 9330 2669
rect 11539 2661 11591 2713
rect 19231 2656 19859 3156
rect 7610 2094 7662 2146
rect 13004 2073 13056 2125
rect 9021 1831 9073 1883
rect 7610 1524 7662 1576
rect 10995 1199 11047 1251
rect 7431 306 8059 806
rect 16899 354 17527 854
<< metal2 >>
rect -1515 5712 -424 5918
rect -1515 5096 -1318 5712
rect -622 5096 -424 5712
rect -1515 4860 -424 5096
rect 16736 5590 17827 5796
rect 7224 4676 7362 5002
rect 16736 4974 16933 5590
rect 17629 4974 17827 5590
rect 7888 4812 9560 4850
rect 7888 4802 9480 4812
rect 7888 4750 7946 4802
rect 7998 4760 9480 4802
rect 9532 4760 9560 4812
rect 7998 4750 9560 4760
rect 7888 4710 9560 4750
rect 16736 4738 17827 4974
rect 7224 4624 7263 4676
rect 7315 4624 7362 4676
rect 7224 4612 7362 4624
rect 7224 4560 7263 4612
rect 7315 4560 7362 4612
rect -1515 4306 -424 4512
rect -1515 3690 -1318 4306
rect -622 3690 -424 4306
rect -1515 3454 -424 3690
rect 5558 3582 5662 3584
rect 1942 3468 3596 3548
rect 1942 3414 3377 3468
rect 3302 3332 3377 3414
rect 3513 3436 3596 3468
rect 3513 3332 3598 3436
rect 5122 3434 5662 3582
rect 3302 3290 3598 3332
rect 5558 3170 5662 3434
rect 7224 3254 7362 4560
rect 6860 3170 6986 3172
rect 5558 3139 6986 3170
rect 5558 3083 6893 3139
rect 6949 3083 6986 3139
rect 5558 3060 6986 3083
rect 6860 3058 6986 3060
rect 7066 3026 7170 3064
rect 7066 2970 7096 3026
rect 7152 2970 7170 3026
rect 4154 2934 4284 2944
rect 7066 2940 7170 2970
rect 4154 2911 7010 2934
rect 4154 2855 4183 2911
rect 4239 2900 7010 2911
rect 4239 2855 6935 2900
rect -1515 2647 -424 2853
rect 4154 2848 6935 2855
rect 6987 2848 7010 2900
rect 4154 2824 7010 2848
rect 4158 2818 7010 2824
rect 6882 2738 6980 2748
rect 6882 2736 6910 2738
rect 6882 2680 6905 2736
rect 6962 2686 6980 2738
rect 6961 2680 6980 2686
rect 6882 2668 6980 2680
rect 7216 2702 7362 3254
rect 18996 3218 20087 3424
rect 8078 3060 8188 3066
rect 7704 3034 8192 3060
rect 7704 3032 7750 3034
rect 7704 2976 7744 3032
rect 7802 3027 8192 3034
rect 7802 2982 8110 3027
rect 7800 2976 8110 2982
rect 7704 2975 8110 2976
rect 8162 2975 8192 3027
rect 7704 2950 8192 2975
rect 11500 2713 11624 2754
rect 7216 2669 9386 2702
rect -1515 2031 -1318 2647
rect -622 2031 -424 2647
rect 7216 2617 9278 2669
rect 9330 2617 9386 2669
rect 7216 2578 9386 2617
rect 7322 2576 9386 2578
rect 11500 2661 11539 2713
rect 11591 2661 11624 2713
rect -1515 1795 -424 2031
rect 7562 2146 7716 2200
rect 7562 2094 7610 2146
rect 7662 2094 7716 2146
rect 7562 1576 7716 2094
rect 11500 2140 11624 2661
rect 18996 2602 19193 3218
rect 19889 2602 20087 3218
rect 18996 2366 20087 2602
rect 12594 2140 13090 2142
rect 11500 2125 13090 2140
rect 11500 2073 13004 2125
rect 13056 2073 13090 2125
rect 11500 2036 13090 2073
rect 7562 1524 7610 1576
rect 7662 1524 7716 1576
rect 7562 1074 7716 1524
rect 8958 1883 9124 1918
rect 8958 1831 9021 1883
rect 9073 1831 9124 1883
rect 8958 1292 9124 1831
rect 8958 1251 11118 1292
rect 8958 1199 10995 1251
rect 11047 1199 11118 1251
rect 8958 1144 11118 1199
rect 7196 868 8287 1074
rect 7196 252 7393 868
rect 8089 252 8287 868
rect 7196 16 8287 252
rect 16664 916 17755 1122
rect 16664 300 16861 916
rect 17557 300 17755 916
rect 16664 64 17755 300
<< via2 >>
rect -1318 5650 -622 5712
rect -1318 5150 -1280 5650
rect -1280 5150 -652 5650
rect -652 5150 -622 5650
rect -1318 5096 -622 5150
rect 16933 5528 17629 5590
rect 16933 5028 16971 5528
rect 16971 5028 17599 5528
rect 17599 5028 17629 5528
rect 16933 4974 17629 5028
rect -1318 4244 -622 4306
rect -1318 3744 -1280 4244
rect -1280 3744 -652 4244
rect -652 3744 -622 4244
rect -1318 3690 -622 3744
rect 3377 3332 3513 3468
rect 6893 3083 6949 3139
rect 7096 3023 7152 3026
rect 7096 2971 7148 3023
rect 7148 2971 7152 3023
rect 7096 2970 7152 2971
rect 4183 2855 4239 2911
rect 6905 2686 6910 2736
rect 6910 2686 6961 2736
rect 6905 2680 6961 2686
rect 7744 2982 7750 3032
rect 7750 2982 7800 3032
rect 7744 2976 7800 2982
rect -1318 2585 -622 2647
rect -1318 2085 -1280 2585
rect -1280 2085 -652 2585
rect -652 2085 -622 2585
rect -1318 2031 -622 2085
rect 19193 3156 19889 3218
rect 19193 2656 19231 3156
rect 19231 2656 19859 3156
rect 19859 2656 19889 3156
rect 19193 2602 19889 2656
rect 7393 806 8089 868
rect 7393 306 7431 806
rect 7431 306 8059 806
rect 8059 306 8089 806
rect 7393 252 8089 306
rect 16861 854 17557 916
rect 16861 354 16899 854
rect 16899 354 17527 854
rect 17527 354 17557 854
rect 16861 300 17557 354
<< metal3 >>
rect -1515 5788 -424 5918
rect -1515 5004 -1406 5788
rect -542 5556 -424 5788
rect 16736 5666 17827 5796
rect -542 5409 1768 5556
rect -542 5004 -424 5409
rect -1515 4860 -424 5004
rect 16736 4882 16845 5666
rect 17709 4882 17827 5666
rect 16736 4738 17827 4882
rect -1515 4382 -424 4512
rect -1515 3598 -1406 4382
rect -542 3598 -424 4382
rect -1515 3454 -424 3598
rect 3274 3472 3634 3554
rect 3274 3328 3373 3472
rect 3517 3328 3634 3472
rect 3274 3302 3634 3328
rect 18996 3294 20087 3424
rect 6866 3139 6988 3170
rect 6866 3083 6893 3139
rect 6949 3083 6988 3139
rect 4066 2915 4290 2960
rect -1515 2723 -424 2853
rect 4066 2851 4179 2915
rect 4243 2851 4290 2915
rect 4066 2806 4290 2851
rect -1515 1939 -1406 2723
rect -542 1939 -424 2723
rect 6866 2736 6988 3083
rect 7100 3066 7892 3068
rect 7064 3032 7892 3066
rect 7064 3026 7744 3032
rect 7064 2970 7096 3026
rect 7152 2976 7744 3026
rect 7800 2976 7892 3032
rect 7152 2970 7892 2976
rect 7064 2952 7892 2970
rect 7064 2938 7186 2952
rect 6866 2680 6905 2736
rect 6961 2680 6988 2736
rect 6866 2656 6988 2680
rect 18996 2510 19105 3294
rect 19969 2510 20087 3294
rect 18996 2366 20087 2510
rect -1515 1795 -424 1939
rect 7196 944 8287 1074
rect 7196 160 7305 944
rect 8169 160 8287 944
rect 7196 16 8287 160
rect 16664 992 17755 1122
rect 16664 208 16773 992
rect 17637 208 17755 992
rect 16664 64 17755 208
<< via3 >>
rect -1406 5712 -542 5788
rect -1406 5096 -1318 5712
rect -1318 5096 -622 5712
rect -622 5096 -542 5712
rect -1406 5004 -542 5096
rect 16845 5590 17709 5666
rect 16845 4974 16933 5590
rect 16933 4974 17629 5590
rect 17629 4974 17709 5590
rect 16845 4882 17709 4974
rect -1406 4306 -542 4382
rect -1406 3690 -1318 4306
rect -1318 3690 -622 4306
rect -622 3690 -542 4306
rect -1406 3598 -542 3690
rect 3373 3468 3517 3472
rect 3373 3332 3377 3468
rect 3377 3332 3513 3468
rect 3513 3332 3517 3468
rect 3373 3328 3517 3332
rect 4179 2911 4243 2915
rect 4179 2855 4183 2911
rect 4183 2855 4239 2911
rect 4239 2855 4243 2911
rect 4179 2851 4243 2855
rect -1406 2647 -542 2723
rect -1406 2031 -1318 2647
rect -1318 2031 -622 2647
rect -622 2031 -542 2647
rect -1406 1939 -542 2031
rect 19105 3218 19969 3294
rect 19105 2602 19193 3218
rect 19193 2602 19889 3218
rect 19889 2602 19969 3218
rect 19105 2510 19969 2602
rect 7305 868 8169 944
rect 7305 252 7393 868
rect 7393 252 8089 868
rect 8089 252 8169 868
rect 7305 160 8169 252
rect 16773 916 17637 992
rect 16773 300 16861 916
rect 16861 300 17557 916
rect 17557 300 17637 916
rect 16773 208 17637 300
<< metal4 >>
rect -1515 5833 -424 5918
rect -1515 4957 -1411 5833
rect -535 4957 -424 5833
rect -1515 4860 -424 4957
rect 16736 5711 17827 5796
rect 16736 4835 16840 5711
rect 17716 4835 17827 5711
rect 16736 4738 17827 4835
rect -1515 4427 -424 4512
rect -1515 3551 -1411 4427
rect -535 3551 -424 4427
rect -1515 3454 -424 3551
rect 3296 3484 3620 3548
rect 3296 3330 3338 3484
rect 3312 3248 3338 3330
rect 3574 3330 3620 3484
rect 18996 3339 20087 3424
rect 3574 3248 3600 3330
rect 3312 3242 3600 3248
rect 3990 3082 4278 3088
rect -1515 2768 -424 2853
rect 3990 2846 4016 3082
rect 4252 2962 4278 3082
rect 4252 2846 4288 2962
rect 3990 2840 4288 2846
rect 4066 2804 4288 2840
rect -1515 1892 -1411 2768
rect -535 2416 -424 2768
rect 18996 2463 19100 3339
rect 19976 2463 20087 3339
rect -535 2206 -104 2416
rect 18996 2366 20087 2463
rect -535 1892 -424 2206
rect -1515 1795 -424 1892
rect 7196 989 8287 1074
rect 7196 113 7300 989
rect 8176 113 8287 989
rect 7196 16 8287 113
rect 16664 1037 17755 1122
rect 16664 161 16768 1037
rect 17644 161 17755 1037
rect 16664 64 17755 161
<< via4 >>
rect -1411 5788 -535 5833
rect -1411 5004 -1406 5788
rect -1406 5004 -542 5788
rect -542 5004 -535 5788
rect -1411 4957 -535 5004
rect 16840 5666 17716 5711
rect 16840 4882 16845 5666
rect 16845 4882 17709 5666
rect 17709 4882 17716 5666
rect 16840 4835 17716 4882
rect -1411 4382 -535 4427
rect -1411 3598 -1406 4382
rect -1406 3598 -542 4382
rect -542 3598 -535 4382
rect -1411 3551 -535 3598
rect 3338 3472 3574 3484
rect 3338 3328 3373 3472
rect 3373 3328 3517 3472
rect 3517 3328 3574 3472
rect 3338 3248 3574 3328
rect 4016 2915 4252 3082
rect 4016 2851 4179 2915
rect 4179 2851 4243 2915
rect 4243 2851 4252 2915
rect 4016 2846 4252 2851
rect -1411 2723 -535 2768
rect -1411 1939 -1406 2723
rect -1406 1939 -542 2723
rect -542 1939 -535 2723
rect 19100 3294 19976 3339
rect 19100 2510 19105 3294
rect 19105 2510 19969 3294
rect 19969 2510 19976 3294
rect 19100 2463 19976 2510
rect -1411 1892 -535 1939
rect 7300 944 8176 989
rect 7300 160 7305 944
rect 7305 160 8169 944
rect 8169 160 8176 944
rect 7300 113 8176 160
rect 16768 992 17644 1037
rect 16768 208 16773 992
rect 16773 208 17637 992
rect 17637 208 17644 992
rect 16768 161 17644 208
<< metal5 >>
rect -1515 5833 -424 5918
rect -1515 4957 -1411 5833
rect -535 4957 -424 5833
rect -1515 4860 -424 4957
rect 16736 5711 17827 5796
rect 16736 4835 16840 5711
rect 17716 4835 17827 5711
rect 16736 4738 17827 4835
rect -1515 4427 -424 4512
rect -1515 3551 -1411 4427
rect -535 3551 -424 4427
rect -1515 3454 -424 3551
rect 3276 3484 3638 3552
rect 3276 3248 3338 3484
rect 3574 3248 3638 3484
rect 3276 3130 3638 3248
rect 18996 3339 20087 3424
rect 3276 3082 4302 3130
rect -1515 2768 -424 2853
rect 3276 2846 4016 3082
rect 4252 2846 4302 3082
rect 3276 2796 4302 2846
rect 3276 2792 3850 2796
rect -1515 1892 -1411 2768
rect -535 1892 -424 2768
rect 18996 2463 19100 3339
rect 19976 2463 20087 3339
rect 18996 2366 20087 2463
rect -1515 1795 -424 1892
rect 7196 989 8287 1074
rect 7196 113 7300 989
rect 8176 113 8287 989
rect 7196 16 8287 113
rect 16664 1037 17755 1122
rect 16664 161 16768 1037
rect 17644 161 17755 1037
rect 16664 64 17755 161
use LVDS2  LVDS2_0
timestamp 1611881054
transform 1 0 9778 0 1 2844
box -152 -1748 5398 2676
use LVDSBias  LVDSBias_0
timestamp 1611881054
transform 1 0 2998 0 1 5224
box -3498 -5188 2356 652
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1611881054
transform 1 0 18732 0 1 2508
box -38 -48 130 592
use LVDS1  LVDS1_0
timestamp 1611881054
transform 1 0 5879 0 1 3380
box -17 -1584 3470 2114
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1611881054
transform 1 0 15566 0 1 2458
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1611881054
transform 1 0 16464 0 1 2476
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1611881054
transform 1 0 17354 0 1 2492
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1611881054
transform 1 0 18380 0 1 2510
box -38 -48 314 592
<< labels >>
rlabel metal1 s 18748 2594 18786 2636 4 OUT
port 1 nsew
<< end >>
