magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -360 840 360 874
rect -360 -840 -326 840
rect 326 -840 360 840
rect -360 -874 360 -840
<< nmoslvt >>
rect -200 -700 200 700
<< ndiff >>
rect -258 663 -200 700
rect -258 629 -246 663
rect -212 629 -200 663
rect -258 595 -200 629
rect -258 561 -246 595
rect -212 561 -200 595
rect -258 527 -200 561
rect -258 493 -246 527
rect -212 493 -200 527
rect -258 459 -200 493
rect -258 425 -246 459
rect -212 425 -200 459
rect -258 391 -200 425
rect -258 357 -246 391
rect -212 357 -200 391
rect -258 323 -200 357
rect -258 289 -246 323
rect -212 289 -200 323
rect -258 255 -200 289
rect -258 221 -246 255
rect -212 221 -200 255
rect -258 187 -200 221
rect -258 153 -246 187
rect -212 153 -200 187
rect -258 119 -200 153
rect -258 85 -246 119
rect -212 85 -200 119
rect -258 51 -200 85
rect -258 17 -246 51
rect -212 17 -200 51
rect -258 -17 -200 17
rect -258 -51 -246 -17
rect -212 -51 -200 -17
rect -258 -85 -200 -51
rect -258 -119 -246 -85
rect -212 -119 -200 -85
rect -258 -153 -200 -119
rect -258 -187 -246 -153
rect -212 -187 -200 -153
rect -258 -221 -200 -187
rect -258 -255 -246 -221
rect -212 -255 -200 -221
rect -258 -289 -200 -255
rect -258 -323 -246 -289
rect -212 -323 -200 -289
rect -258 -357 -200 -323
rect -258 -391 -246 -357
rect -212 -391 -200 -357
rect -258 -425 -200 -391
rect -258 -459 -246 -425
rect -212 -459 -200 -425
rect -258 -493 -200 -459
rect -258 -527 -246 -493
rect -212 -527 -200 -493
rect -258 -561 -200 -527
rect -258 -595 -246 -561
rect -212 -595 -200 -561
rect -258 -629 -200 -595
rect -258 -663 -246 -629
rect -212 -663 -200 -629
rect -258 -700 -200 -663
rect 200 663 258 700
rect 200 629 212 663
rect 246 629 258 663
rect 200 595 258 629
rect 200 561 212 595
rect 246 561 258 595
rect 200 527 258 561
rect 200 493 212 527
rect 246 493 258 527
rect 200 459 258 493
rect 200 425 212 459
rect 246 425 258 459
rect 200 391 258 425
rect 200 357 212 391
rect 246 357 258 391
rect 200 323 258 357
rect 200 289 212 323
rect 246 289 258 323
rect 200 255 258 289
rect 200 221 212 255
rect 246 221 258 255
rect 200 187 258 221
rect 200 153 212 187
rect 246 153 258 187
rect 200 119 258 153
rect 200 85 212 119
rect 246 85 258 119
rect 200 51 258 85
rect 200 17 212 51
rect 246 17 258 51
rect 200 -17 258 17
rect 200 -51 212 -17
rect 246 -51 258 -17
rect 200 -85 258 -51
rect 200 -119 212 -85
rect 246 -119 258 -85
rect 200 -153 258 -119
rect 200 -187 212 -153
rect 246 -187 258 -153
rect 200 -221 258 -187
rect 200 -255 212 -221
rect 246 -255 258 -221
rect 200 -289 258 -255
rect 200 -323 212 -289
rect 246 -323 258 -289
rect 200 -357 258 -323
rect 200 -391 212 -357
rect 246 -391 258 -357
rect 200 -425 258 -391
rect 200 -459 212 -425
rect 246 -459 258 -425
rect 200 -493 258 -459
rect 200 -527 212 -493
rect 246 -527 258 -493
rect 200 -561 258 -527
rect 200 -595 212 -561
rect 246 -595 258 -561
rect 200 -629 258 -595
rect 200 -663 212 -629
rect 246 -663 258 -629
rect 200 -700 258 -663
<< ndiffc >>
rect -246 629 -212 663
rect -246 561 -212 595
rect -246 493 -212 527
rect -246 425 -212 459
rect -246 357 -212 391
rect -246 289 -212 323
rect -246 221 -212 255
rect -246 153 -212 187
rect -246 85 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -85
rect -246 -187 -212 -153
rect -246 -255 -212 -221
rect -246 -323 -212 -289
rect -246 -391 -212 -357
rect -246 -459 -212 -425
rect -246 -527 -212 -493
rect -246 -595 -212 -561
rect -246 -663 -212 -629
rect 212 629 246 663
rect 212 561 246 595
rect 212 493 246 527
rect 212 425 246 459
rect 212 357 246 391
rect 212 289 246 323
rect 212 221 246 255
rect 212 153 246 187
rect 212 85 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -85
rect 212 -187 246 -153
rect 212 -255 246 -221
rect 212 -323 246 -289
rect 212 -391 246 -357
rect 212 -459 246 -425
rect 212 -527 246 -493
rect 212 -595 246 -561
rect 212 -663 246 -629
<< psubdiff >>
rect -360 840 -255 874
rect -221 840 -187 874
rect -153 840 -119 874
rect -85 840 -51 874
rect -17 840 17 874
rect 51 840 85 874
rect 119 840 153 874
rect 187 840 221 874
rect 255 840 360 874
rect -360 765 -326 840
rect -360 697 -326 731
rect 326 765 360 840
rect -360 629 -326 663
rect -360 561 -326 595
rect -360 493 -326 527
rect -360 425 -326 459
rect -360 357 -326 391
rect -360 289 -326 323
rect -360 221 -326 255
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect -360 -255 -326 -221
rect -360 -323 -326 -289
rect -360 -391 -326 -357
rect -360 -459 -326 -425
rect -360 -527 -326 -493
rect -360 -595 -326 -561
rect -360 -663 -326 -629
rect -360 -731 -326 -697
rect 326 697 360 731
rect 326 629 360 663
rect 326 561 360 595
rect 326 493 360 527
rect 326 425 360 459
rect 326 357 360 391
rect 326 289 360 323
rect 326 221 360 255
rect 326 153 360 187
rect 326 85 360 119
rect 326 17 360 51
rect 326 -51 360 -17
rect 326 -119 360 -85
rect 326 -187 360 -153
rect 326 -255 360 -221
rect 326 -323 360 -289
rect 326 -391 360 -357
rect 326 -459 360 -425
rect 326 -527 360 -493
rect 326 -595 360 -561
rect 326 -663 360 -629
rect -360 -840 -326 -765
rect 326 -731 360 -697
rect 326 -840 360 -765
rect -360 -874 -255 -840
rect -221 -874 -187 -840
rect -153 -874 -119 -840
rect -85 -874 -51 -840
rect -17 -874 17 -840
rect 51 -874 85 -840
rect 119 -874 153 -840
rect 187 -874 221 -840
rect 255 -874 360 -840
<< psubdiffcont >>
rect -255 840 -221 874
rect -187 840 -153 874
rect -119 840 -85 874
rect -51 840 -17 874
rect 17 840 51 874
rect 85 840 119 874
rect 153 840 187 874
rect 221 840 255 874
rect -360 731 -326 765
rect 326 731 360 765
rect -360 663 -326 697
rect -360 595 -326 629
rect -360 527 -326 561
rect -360 459 -326 493
rect -360 391 -326 425
rect -360 323 -326 357
rect -360 255 -326 289
rect -360 187 -326 221
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
rect -360 -289 -326 -255
rect -360 -357 -326 -323
rect -360 -425 -326 -391
rect -360 -493 -326 -459
rect -360 -561 -326 -527
rect -360 -629 -326 -595
rect -360 -697 -326 -663
rect 326 663 360 697
rect 326 595 360 629
rect 326 527 360 561
rect 326 459 360 493
rect 326 391 360 425
rect 326 323 360 357
rect 326 255 360 289
rect 326 187 360 221
rect 326 119 360 153
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect 326 -153 360 -119
rect 326 -221 360 -187
rect 326 -289 360 -255
rect 326 -357 360 -323
rect 326 -425 360 -391
rect 326 -493 360 -459
rect 326 -561 360 -527
rect 326 -629 360 -595
rect 326 -697 360 -663
rect -360 -765 -326 -731
rect 326 -765 360 -731
rect -255 -874 -221 -840
rect -187 -874 -153 -840
rect -119 -874 -85 -840
rect -51 -874 -17 -840
rect 17 -874 51 -840
rect 85 -874 119 -840
rect 153 -874 187 -840
rect 221 -874 255 -840
<< poly >>
rect -200 772 200 788
rect -200 738 -153 772
rect -119 738 -85 772
rect -51 738 -17 772
rect 17 738 51 772
rect 85 738 119 772
rect 153 738 200 772
rect -200 700 200 738
rect -200 -738 200 -700
rect -200 -772 -153 -738
rect -119 -772 -85 -738
rect -51 -772 -17 -738
rect 17 -772 51 -738
rect 85 -772 119 -738
rect 153 -772 200 -738
rect -200 -788 200 -772
<< polycont >>
rect -153 738 -119 772
rect -85 738 -51 772
rect -17 738 17 772
rect 51 738 85 772
rect 119 738 153 772
rect -153 -772 -119 -738
rect -85 -772 -51 -738
rect -17 -772 17 -738
rect 51 -772 85 -738
rect 119 -772 153 -738
<< locali >>
rect -360 840 -255 874
rect -221 840 -187 874
rect -153 840 -119 874
rect -85 840 -51 874
rect -17 840 17 874
rect 51 840 85 874
rect 119 840 153 874
rect 187 840 221 874
rect 255 840 360 874
rect -360 765 -326 840
rect -200 738 -153 772
rect -119 738 -85 772
rect -51 738 -17 772
rect 17 738 51 772
rect 85 738 119 772
rect 153 738 200 772
rect 326 765 360 840
rect -360 697 -326 731
rect -360 629 -326 663
rect -360 561 -326 595
rect -360 493 -326 527
rect -360 425 -326 459
rect -360 357 -326 391
rect -360 289 -326 323
rect -360 221 -326 255
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect -360 -255 -326 -221
rect -360 -323 -326 -289
rect -360 -391 -326 -357
rect -360 -459 -326 -425
rect -360 -527 -326 -493
rect -360 -595 -326 -561
rect -360 -663 -326 -629
rect -360 -731 -326 -697
rect -246 663 -212 704
rect -246 595 -212 629
rect -246 527 -212 561
rect -246 459 -212 493
rect -246 391 -212 425
rect -246 323 -212 357
rect -246 255 -212 289
rect -246 187 -212 221
rect -246 119 -212 153
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect -246 -153 -212 -119
rect -246 -221 -212 -187
rect -246 -289 -212 -255
rect -246 -357 -212 -323
rect -246 -425 -212 -391
rect -246 -493 -212 -459
rect -246 -561 -212 -527
rect -246 -629 -212 -595
rect -246 -704 -212 -663
rect 212 663 246 704
rect 212 595 246 629
rect 212 527 246 561
rect 212 459 246 493
rect 212 391 246 425
rect 212 323 246 357
rect 212 255 246 289
rect 212 187 246 221
rect 212 119 246 153
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
rect 212 -153 246 -119
rect 212 -221 246 -187
rect 212 -289 246 -255
rect 212 -357 246 -323
rect 212 -425 246 -391
rect 212 -493 246 -459
rect 212 -561 246 -527
rect 212 -629 246 -595
rect 212 -704 246 -663
rect 326 697 360 731
rect 326 629 360 663
rect 326 561 360 595
rect 326 493 360 527
rect 326 425 360 459
rect 326 357 360 391
rect 326 289 360 323
rect 326 221 360 255
rect 326 153 360 187
rect 326 85 360 119
rect 326 17 360 51
rect 326 -51 360 -17
rect 326 -119 360 -85
rect 326 -187 360 -153
rect 326 -255 360 -221
rect 326 -323 360 -289
rect 326 -391 360 -357
rect 326 -459 360 -425
rect 326 -527 360 -493
rect 326 -595 360 -561
rect 326 -663 360 -629
rect 326 -731 360 -697
rect -360 -840 -326 -765
rect -200 -772 -153 -738
rect -119 -772 -85 -738
rect -51 -772 -17 -738
rect 17 -772 51 -738
rect 85 -772 119 -738
rect 153 -772 200 -738
rect 326 -840 360 -765
rect -360 -874 -255 -840
rect -221 -874 -187 -840
rect -153 -874 -119 -840
rect -85 -874 -51 -840
rect -17 -874 17 -840
rect 51 -874 85 -840
rect 119 -874 153 -840
rect 187 -874 221 -840
rect 255 -874 360 -840
<< properties >>
string FIXED_BBOX -342 -856 342 856
<< end >>
