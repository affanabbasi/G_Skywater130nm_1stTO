magic
tech sky130A
timestamp 1607293554
<< nwell >>
rect 5043 3888 10735 3916
rect 14736 3912 21141 3916
rect 25305 3912 31710 3916
rect 14684 3911 21141 3912
rect 25253 3911 31710 3912
rect 14483 3908 21141 3911
rect 25052 3908 31710 3911
rect 13075 3906 21141 3908
rect 23644 3906 31710 3908
rect 11804 3888 21141 3906
rect 22373 3888 31710 3906
rect 5043 2496 31710 3888
rect 5043 2485 10735 2496
rect 11653 2493 21445 2496
rect 11653 2492 12054 2493
rect 13042 2485 21445 2493
rect 22222 2493 31710 2496
rect 22222 2492 22623 2493
rect 23611 2485 31710 2493
rect 8090 2480 9173 2485
rect 13394 2480 14477 2485
rect 18658 2480 19741 2485
rect 23963 2480 25046 2485
rect 29227 2480 30310 2485
<< pwell >>
rect 7134 2141 8682 2143
rect 12438 2141 13986 2143
rect 17702 2141 19250 2143
rect 23007 2141 24555 2143
rect 28271 2141 29819 2143
rect 7134 2136 9870 2141
rect 12438 2136 15174 2141
rect 17702 2136 20438 2141
rect 23007 2136 25743 2141
rect 28271 2136 31007 2141
rect 5935 1930 9870 2136
rect 11239 1930 15174 2136
rect 16503 1930 20438 2136
rect 21808 1930 25743 2136
rect 27072 1930 31007 2136
rect 5935 1925 8682 1930
rect 11239 1925 13986 1930
rect 16503 1925 19250 1930
rect 21808 1925 24555 1930
rect 27072 1925 29819 1930
rect 7134 1923 8682 1925
rect 12438 1923 13986 1925
rect 17702 1923 19250 1925
rect 23007 1923 24555 1925
rect 28271 1923 29819 1925
rect 7139 221 9825 1631
rect 12443 221 15129 1631
rect 17707 221 20393 1631
rect 23012 221 25698 1631
rect 28276 221 30962 1631
<< pmos >>
rect 6780 2602 6980 3602
rect 7009 2602 7209 3602
rect 7238 2602 7438 3602
rect 7467 2602 7667 3602
rect 12084 2602 12284 3602
rect 12313 2602 12513 3602
rect 12542 2602 12742 3602
rect 12771 2602 12971 3602
rect 17348 2602 17548 3602
rect 17577 2602 17777 3602
rect 17806 2602 18006 3602
rect 18035 2602 18235 3602
rect 22653 2602 22853 3602
rect 22882 2602 23082 3602
rect 23111 2602 23311 3602
rect 23340 2602 23540 3602
rect 27917 2602 28117 3602
rect 28146 2602 28346 3602
rect 28375 2602 28575 3602
rect 28604 2602 28804 3602
<< pmoslvt >>
rect 5403 2605 5603 3605
rect 5632 2605 5832 3605
rect 5861 2605 6061 3605
rect 6090 2605 6290 3605
rect 8188 2589 8388 3589
rect 8417 2589 8617 3589
rect 8646 2589 8846 3589
rect 8875 2589 9075 3589
rect 9450 2600 9650 3600
rect 9679 2600 9879 3600
rect 9908 2600 10108 3600
rect 10137 2600 10337 3600
rect 10707 2605 10907 3605
rect 10936 2605 11136 3605
rect 11165 2605 11365 3605
rect 11394 2605 11594 3605
rect 13492 2589 13692 3589
rect 13721 2589 13921 3589
rect 13950 2589 14150 3589
rect 14179 2589 14379 3589
rect 14754 2600 14954 3600
rect 14983 2600 15183 3600
rect 15212 2600 15412 3600
rect 15441 2600 15641 3600
rect 15971 2605 16171 3605
rect 16200 2605 16400 3605
rect 16429 2605 16629 3605
rect 16658 2605 16858 3605
rect 18756 2589 18956 3589
rect 18985 2589 19185 3589
rect 19214 2589 19414 3589
rect 19443 2589 19643 3589
rect 20018 2600 20218 3600
rect 20247 2600 20447 3600
rect 20476 2600 20676 3600
rect 20705 2600 20905 3600
rect 21276 2605 21476 3605
rect 21505 2605 21705 3605
rect 21734 2605 21934 3605
rect 21963 2605 22163 3605
rect 24061 2589 24261 3589
rect 24290 2589 24490 3589
rect 24519 2589 24719 3589
rect 24748 2589 24948 3589
rect 25323 2600 25523 3600
rect 25552 2600 25752 3600
rect 25781 2600 25981 3600
rect 26010 2600 26210 3600
rect 26540 2605 26740 3605
rect 26769 2605 26969 3605
rect 26998 2605 27198 3605
rect 27227 2605 27427 3605
rect 29325 2589 29525 3589
rect 29554 2589 29754 3589
rect 29783 2589 29983 3589
rect 30012 2589 30212 3589
rect 30587 2600 30787 3600
rect 30816 2600 31016 3600
rect 31045 2600 31245 3600
rect 31274 2600 31474 3600
<< nmoslvt >>
rect 6040 2023 7040 2038
rect 8765 2028 9765 2043
rect 11344 2023 12344 2038
rect 14069 2028 15069 2043
rect 16608 2023 17608 2038
rect 19333 2028 20333 2043
rect 21913 2023 22913 2038
rect 24638 2028 25638 2043
rect 27177 2023 28177 2038
rect 29902 2028 30902 2043
rect 7237 326 7437 1526
rect 7466 326 7666 1526
rect 7695 326 7895 1526
rect 7924 326 8124 1526
rect 8153 326 8353 1526
rect 8382 326 8582 1526
rect 8611 326 8811 1526
rect 8840 326 9040 1526
rect 9069 326 9269 1526
rect 9298 326 9498 1526
rect 9527 326 9727 1526
rect 12541 326 12741 1526
rect 12770 326 12970 1526
rect 12999 326 13199 1526
rect 13228 326 13428 1526
rect 13457 326 13657 1526
rect 13686 326 13886 1526
rect 13915 326 14115 1526
rect 14144 326 14344 1526
rect 14373 326 14573 1526
rect 14602 326 14802 1526
rect 14831 326 15031 1526
rect 17805 326 18005 1526
rect 18034 326 18234 1526
rect 18263 326 18463 1526
rect 18492 326 18692 1526
rect 18721 326 18921 1526
rect 18950 326 19150 1526
rect 19179 326 19379 1526
rect 19408 326 19608 1526
rect 19637 326 19837 1526
rect 19866 326 20066 1526
rect 20095 326 20295 1526
rect 23110 326 23310 1526
rect 23339 326 23539 1526
rect 23568 326 23768 1526
rect 23797 326 23997 1526
rect 24026 326 24226 1526
rect 24255 326 24455 1526
rect 24484 326 24684 1526
rect 24713 326 24913 1526
rect 24942 326 25142 1526
rect 25171 326 25371 1526
rect 25400 326 25600 1526
rect 28374 326 28574 1526
rect 28603 326 28803 1526
rect 28832 326 29032 1526
rect 29061 326 29261 1526
rect 29290 326 29490 1526
rect 29519 326 29719 1526
rect 29748 326 29948 1526
rect 29977 326 30177 1526
rect 30206 326 30406 1526
rect 30435 326 30635 1526
rect 30664 326 30864 1526
<< ndiff >>
rect 6040 2061 7040 2067
rect 6040 2044 6046 2061
rect 7034 2044 7040 2061
rect 6040 2038 7040 2044
rect 6040 2017 7040 2023
rect 6040 2000 6046 2017
rect 7034 2000 7040 2017
rect 6040 1994 7040 2000
rect 8765 2066 9765 2072
rect 8765 2049 8771 2066
rect 9759 2049 9765 2066
rect 8765 2043 9765 2049
rect 8765 2022 9765 2028
rect 8765 2005 8771 2022
rect 9759 2005 9765 2022
rect 8765 1999 9765 2005
rect 11344 2061 12344 2067
rect 11344 2044 11350 2061
rect 12338 2044 12344 2061
rect 11344 2038 12344 2044
rect 11344 2017 12344 2023
rect 11344 2000 11350 2017
rect 12338 2000 12344 2017
rect 11344 1994 12344 2000
rect 14069 2066 15069 2072
rect 14069 2049 14075 2066
rect 15063 2049 15069 2066
rect 14069 2043 15069 2049
rect 14069 2022 15069 2028
rect 14069 2005 14075 2022
rect 15063 2005 15069 2022
rect 14069 1999 15069 2005
rect 16608 2061 17608 2067
rect 16608 2044 16614 2061
rect 17602 2044 17608 2061
rect 16608 2038 17608 2044
rect 16608 2017 17608 2023
rect 16608 2000 16614 2017
rect 17602 2000 17608 2017
rect 16608 1994 17608 2000
rect 19333 2066 20333 2072
rect 19333 2049 19339 2066
rect 20327 2049 20333 2066
rect 19333 2043 20333 2049
rect 19333 2022 20333 2028
rect 19333 2005 19339 2022
rect 20327 2005 20333 2022
rect 19333 1999 20333 2005
rect 21913 2061 22913 2067
rect 21913 2044 21919 2061
rect 22907 2044 22913 2061
rect 21913 2038 22913 2044
rect 21913 2017 22913 2023
rect 21913 2000 21919 2017
rect 22907 2000 22913 2017
rect 21913 1994 22913 2000
rect 24638 2066 25638 2072
rect 24638 2049 24644 2066
rect 25632 2049 25638 2066
rect 24638 2043 25638 2049
rect 24638 2022 25638 2028
rect 24638 2005 24644 2022
rect 25632 2005 25638 2022
rect 24638 1999 25638 2005
rect 27177 2061 28177 2067
rect 27177 2044 27183 2061
rect 28171 2044 28177 2061
rect 27177 2038 28177 2044
rect 27177 2017 28177 2023
rect 27177 2000 27183 2017
rect 28171 2000 28177 2017
rect 27177 1994 28177 2000
rect 29902 2066 30902 2072
rect 29902 2049 29908 2066
rect 30896 2049 30902 2066
rect 29902 2043 30902 2049
rect 29902 2022 30902 2028
rect 29902 2005 29908 2022
rect 30896 2005 30902 2022
rect 29902 1999 30902 2005
rect 7208 1520 7237 1526
rect 7208 332 7214 1520
rect 7231 332 7237 1520
rect 7208 326 7237 332
rect 7437 1520 7466 1526
rect 7437 332 7443 1520
rect 7460 332 7466 1520
rect 7437 326 7466 332
rect 7666 1520 7695 1526
rect 7666 332 7672 1520
rect 7689 332 7695 1520
rect 7666 326 7695 332
rect 7895 1520 7924 1526
rect 7895 332 7901 1520
rect 7918 332 7924 1520
rect 7895 326 7924 332
rect 8124 1520 8153 1526
rect 8124 332 8130 1520
rect 8147 332 8153 1520
rect 8124 326 8153 332
rect 8353 1520 8382 1526
rect 8353 332 8359 1520
rect 8376 332 8382 1520
rect 8353 326 8382 332
rect 8582 1520 8611 1526
rect 8582 332 8588 1520
rect 8605 332 8611 1520
rect 8582 326 8611 332
rect 8811 1520 8840 1526
rect 8811 332 8817 1520
rect 8834 332 8840 1520
rect 8811 326 8840 332
rect 9040 1520 9069 1526
rect 9040 332 9046 1520
rect 9063 332 9069 1520
rect 9040 326 9069 332
rect 9269 1520 9298 1526
rect 9269 332 9275 1520
rect 9292 332 9298 1520
rect 9269 326 9298 332
rect 9498 1520 9527 1526
rect 9498 332 9504 1520
rect 9521 332 9527 1520
rect 9498 326 9527 332
rect 9727 1520 9756 1526
rect 9727 332 9733 1520
rect 9750 332 9756 1520
rect 9727 326 9756 332
rect 12512 1520 12541 1526
rect 12512 332 12518 1520
rect 12535 332 12541 1520
rect 12512 326 12541 332
rect 12741 1520 12770 1526
rect 12741 332 12747 1520
rect 12764 332 12770 1520
rect 12741 326 12770 332
rect 12970 1520 12999 1526
rect 12970 332 12976 1520
rect 12993 332 12999 1520
rect 12970 326 12999 332
rect 13199 1520 13228 1526
rect 13199 332 13205 1520
rect 13222 332 13228 1520
rect 13199 326 13228 332
rect 13428 1520 13457 1526
rect 13428 332 13434 1520
rect 13451 332 13457 1520
rect 13428 326 13457 332
rect 13657 1520 13686 1526
rect 13657 332 13663 1520
rect 13680 332 13686 1520
rect 13657 326 13686 332
rect 13886 1520 13915 1526
rect 13886 332 13892 1520
rect 13909 332 13915 1520
rect 13886 326 13915 332
rect 14115 1520 14144 1526
rect 14115 332 14121 1520
rect 14138 332 14144 1520
rect 14115 326 14144 332
rect 14344 1520 14373 1526
rect 14344 332 14350 1520
rect 14367 332 14373 1520
rect 14344 326 14373 332
rect 14573 1520 14602 1526
rect 14573 332 14579 1520
rect 14596 332 14602 1520
rect 14573 326 14602 332
rect 14802 1520 14831 1526
rect 14802 332 14808 1520
rect 14825 332 14831 1520
rect 14802 326 14831 332
rect 15031 1520 15060 1526
rect 15031 332 15037 1520
rect 15054 332 15060 1520
rect 15031 326 15060 332
rect 17776 1520 17805 1526
rect 17776 332 17782 1520
rect 17799 332 17805 1520
rect 17776 326 17805 332
rect 18005 1520 18034 1526
rect 18005 332 18011 1520
rect 18028 332 18034 1520
rect 18005 326 18034 332
rect 18234 1520 18263 1526
rect 18234 332 18240 1520
rect 18257 332 18263 1520
rect 18234 326 18263 332
rect 18463 1520 18492 1526
rect 18463 332 18469 1520
rect 18486 332 18492 1520
rect 18463 326 18492 332
rect 18692 1520 18721 1526
rect 18692 332 18698 1520
rect 18715 332 18721 1520
rect 18692 326 18721 332
rect 18921 1520 18950 1526
rect 18921 332 18927 1520
rect 18944 332 18950 1520
rect 18921 326 18950 332
rect 19150 1520 19179 1526
rect 19150 332 19156 1520
rect 19173 332 19179 1520
rect 19150 326 19179 332
rect 19379 1520 19408 1526
rect 19379 332 19385 1520
rect 19402 332 19408 1520
rect 19379 326 19408 332
rect 19608 1520 19637 1526
rect 19608 332 19614 1520
rect 19631 332 19637 1520
rect 19608 326 19637 332
rect 19837 1520 19866 1526
rect 19837 332 19843 1520
rect 19860 332 19866 1520
rect 19837 326 19866 332
rect 20066 1520 20095 1526
rect 20066 332 20072 1520
rect 20089 332 20095 1520
rect 20066 326 20095 332
rect 20295 1520 20324 1526
rect 20295 332 20301 1520
rect 20318 332 20324 1520
rect 20295 326 20324 332
rect 23081 1520 23110 1526
rect 23081 332 23087 1520
rect 23104 332 23110 1520
rect 23081 326 23110 332
rect 23310 1520 23339 1526
rect 23310 332 23316 1520
rect 23333 332 23339 1520
rect 23310 326 23339 332
rect 23539 1520 23568 1526
rect 23539 332 23545 1520
rect 23562 332 23568 1520
rect 23539 326 23568 332
rect 23768 1520 23797 1526
rect 23768 332 23774 1520
rect 23791 332 23797 1520
rect 23768 326 23797 332
rect 23997 1520 24026 1526
rect 23997 332 24003 1520
rect 24020 332 24026 1520
rect 23997 326 24026 332
rect 24226 1520 24255 1526
rect 24226 332 24232 1520
rect 24249 332 24255 1520
rect 24226 326 24255 332
rect 24455 1520 24484 1526
rect 24455 332 24461 1520
rect 24478 332 24484 1520
rect 24455 326 24484 332
rect 24684 1520 24713 1526
rect 24684 332 24690 1520
rect 24707 332 24713 1520
rect 24684 326 24713 332
rect 24913 1520 24942 1526
rect 24913 332 24919 1520
rect 24936 332 24942 1520
rect 24913 326 24942 332
rect 25142 1520 25171 1526
rect 25142 332 25148 1520
rect 25165 332 25171 1520
rect 25142 326 25171 332
rect 25371 1520 25400 1526
rect 25371 332 25377 1520
rect 25394 332 25400 1520
rect 25371 326 25400 332
rect 25600 1520 25629 1526
rect 25600 332 25606 1520
rect 25623 332 25629 1520
rect 25600 326 25629 332
rect 28345 1520 28374 1526
rect 28345 332 28351 1520
rect 28368 332 28374 1520
rect 28345 326 28374 332
rect 28574 1520 28603 1526
rect 28574 332 28580 1520
rect 28597 332 28603 1520
rect 28574 326 28603 332
rect 28803 1520 28832 1526
rect 28803 332 28809 1520
rect 28826 332 28832 1520
rect 28803 326 28832 332
rect 29032 1520 29061 1526
rect 29032 332 29038 1520
rect 29055 332 29061 1520
rect 29032 326 29061 332
rect 29261 1520 29290 1526
rect 29261 332 29267 1520
rect 29284 332 29290 1520
rect 29261 326 29290 332
rect 29490 1520 29519 1526
rect 29490 332 29496 1520
rect 29513 332 29519 1520
rect 29490 326 29519 332
rect 29719 1520 29748 1526
rect 29719 332 29725 1520
rect 29742 332 29748 1520
rect 29719 326 29748 332
rect 29948 1520 29977 1526
rect 29948 332 29954 1520
rect 29971 332 29977 1520
rect 29948 326 29977 332
rect 30177 1520 30206 1526
rect 30177 332 30183 1520
rect 30200 332 30206 1520
rect 30177 326 30206 332
rect 30406 1520 30435 1526
rect 30406 332 30412 1520
rect 30429 332 30435 1520
rect 30406 326 30435 332
rect 30635 1520 30664 1526
rect 30635 332 30641 1520
rect 30658 332 30664 1520
rect 30635 326 30664 332
rect 30864 1520 30893 1526
rect 30864 332 30870 1520
rect 30887 332 30893 1520
rect 30864 326 30893 332
<< pdiff >>
rect 5374 3599 5403 3605
rect 5374 2611 5380 3599
rect 5397 2611 5403 3599
rect 5374 2605 5403 2611
rect 5603 3599 5632 3605
rect 5603 2611 5609 3599
rect 5626 2611 5632 3599
rect 5603 2605 5632 2611
rect 5832 3599 5861 3605
rect 5832 2611 5838 3599
rect 5855 2611 5861 3599
rect 5832 2605 5861 2611
rect 6061 3599 6090 3605
rect 6061 2611 6067 3599
rect 6084 2611 6090 3599
rect 6061 2605 6090 2611
rect 6290 3599 6319 3605
rect 6290 2611 6296 3599
rect 6313 2611 6319 3599
rect 6290 2605 6319 2611
rect 6751 3596 6780 3602
rect 6751 2608 6757 3596
rect 6774 2608 6780 3596
rect 6751 2602 6780 2608
rect 6980 3596 7009 3602
rect 6980 2608 6986 3596
rect 7003 2608 7009 3596
rect 6980 2602 7009 2608
rect 7209 3596 7238 3602
rect 7209 2608 7215 3596
rect 7232 2608 7238 3596
rect 7209 2602 7238 2608
rect 7438 3596 7467 3602
rect 7438 2608 7444 3596
rect 7461 2608 7467 3596
rect 7438 2602 7467 2608
rect 7667 3596 7696 3602
rect 7667 2608 7673 3596
rect 7690 2608 7696 3596
rect 7667 2602 7696 2608
rect 8159 3583 8188 3589
rect 8159 2595 8165 3583
rect 8182 2595 8188 3583
rect 8159 2589 8188 2595
rect 8388 3583 8417 3589
rect 8388 2595 8394 3583
rect 8411 2595 8417 3583
rect 8388 2589 8417 2595
rect 8617 3583 8646 3589
rect 8617 2595 8623 3583
rect 8640 2595 8646 3583
rect 8617 2589 8646 2595
rect 8846 3583 8875 3589
rect 8846 2595 8852 3583
rect 8869 2595 8875 3583
rect 8846 2589 8875 2595
rect 9075 3583 9104 3589
rect 9075 2595 9081 3583
rect 9098 2595 9104 3583
rect 9075 2589 9104 2595
rect 9421 3594 9450 3600
rect 9421 2606 9427 3594
rect 9444 2606 9450 3594
rect 9421 2600 9450 2606
rect 9650 3594 9679 3600
rect 9650 2606 9656 3594
rect 9673 2606 9679 3594
rect 9650 2600 9679 2606
rect 9879 3594 9908 3600
rect 9879 2606 9885 3594
rect 9902 2606 9908 3594
rect 9879 2600 9908 2606
rect 10108 3594 10137 3600
rect 10108 2606 10114 3594
rect 10131 2606 10137 3594
rect 10108 2600 10137 2606
rect 10337 3594 10366 3600
rect 10337 2606 10343 3594
rect 10360 2606 10366 3594
rect 10337 2600 10366 2606
rect 10678 3599 10707 3605
rect 10678 2611 10684 3599
rect 10701 2611 10707 3599
rect 10678 2605 10707 2611
rect 10907 3599 10936 3605
rect 10907 2611 10913 3599
rect 10930 2611 10936 3599
rect 10907 2605 10936 2611
rect 11136 3599 11165 3605
rect 11136 2611 11142 3599
rect 11159 2611 11165 3599
rect 11136 2605 11165 2611
rect 11365 3599 11394 3605
rect 11365 2611 11371 3599
rect 11388 2611 11394 3599
rect 11365 2605 11394 2611
rect 11594 3599 11623 3605
rect 11594 2611 11600 3599
rect 11617 2611 11623 3599
rect 11594 2605 11623 2611
rect 12055 3596 12084 3602
rect 12055 2608 12061 3596
rect 12078 2608 12084 3596
rect 12055 2602 12084 2608
rect 12284 3596 12313 3602
rect 12284 2608 12290 3596
rect 12307 2608 12313 3596
rect 12284 2602 12313 2608
rect 12513 3596 12542 3602
rect 12513 2608 12519 3596
rect 12536 2608 12542 3596
rect 12513 2602 12542 2608
rect 12742 3596 12771 3602
rect 12742 2608 12748 3596
rect 12765 2608 12771 3596
rect 12742 2602 12771 2608
rect 12971 3596 13000 3602
rect 12971 2608 12977 3596
rect 12994 2608 13000 3596
rect 12971 2602 13000 2608
rect 13463 3583 13492 3589
rect 13463 2595 13469 3583
rect 13486 2595 13492 3583
rect 13463 2589 13492 2595
rect 13692 3583 13721 3589
rect 13692 2595 13698 3583
rect 13715 2595 13721 3583
rect 13692 2589 13721 2595
rect 13921 3583 13950 3589
rect 13921 2595 13927 3583
rect 13944 2595 13950 3583
rect 13921 2589 13950 2595
rect 14150 3583 14179 3589
rect 14150 2595 14156 3583
rect 14173 2595 14179 3583
rect 14150 2589 14179 2595
rect 14379 3583 14408 3589
rect 14379 2595 14385 3583
rect 14402 2595 14408 3583
rect 14379 2589 14408 2595
rect 14725 3594 14754 3600
rect 14725 2606 14731 3594
rect 14748 2606 14754 3594
rect 14725 2600 14754 2606
rect 14954 3594 14983 3600
rect 14954 2606 14960 3594
rect 14977 2606 14983 3594
rect 14954 2600 14983 2606
rect 15183 3594 15212 3600
rect 15183 2606 15189 3594
rect 15206 2606 15212 3594
rect 15183 2600 15212 2606
rect 15412 3594 15441 3600
rect 15412 2606 15418 3594
rect 15435 2606 15441 3594
rect 15412 2600 15441 2606
rect 15641 3594 15670 3600
rect 15641 2606 15647 3594
rect 15664 2606 15670 3594
rect 15641 2600 15670 2606
rect 15942 3599 15971 3605
rect 15942 2611 15948 3599
rect 15965 2611 15971 3599
rect 15942 2605 15971 2611
rect 16171 3599 16200 3605
rect 16171 2611 16177 3599
rect 16194 2611 16200 3599
rect 16171 2605 16200 2611
rect 16400 3599 16429 3605
rect 16400 2611 16406 3599
rect 16423 2611 16429 3599
rect 16400 2605 16429 2611
rect 16629 3599 16658 3605
rect 16629 2611 16635 3599
rect 16652 2611 16658 3599
rect 16629 2605 16658 2611
rect 16858 3599 16887 3605
rect 16858 2611 16864 3599
rect 16881 2611 16887 3599
rect 16858 2605 16887 2611
rect 17319 3596 17348 3602
rect 17319 2608 17325 3596
rect 17342 2608 17348 3596
rect 17319 2602 17348 2608
rect 17548 3596 17577 3602
rect 17548 2608 17554 3596
rect 17571 2608 17577 3596
rect 17548 2602 17577 2608
rect 17777 3596 17806 3602
rect 17777 2608 17783 3596
rect 17800 2608 17806 3596
rect 17777 2602 17806 2608
rect 18006 3596 18035 3602
rect 18006 2608 18012 3596
rect 18029 2608 18035 3596
rect 18006 2602 18035 2608
rect 18235 3596 18264 3602
rect 18235 2608 18241 3596
rect 18258 2608 18264 3596
rect 18235 2602 18264 2608
rect 18727 3583 18756 3589
rect 18727 2595 18733 3583
rect 18750 2595 18756 3583
rect 18727 2589 18756 2595
rect 18956 3583 18985 3589
rect 18956 2595 18962 3583
rect 18979 2595 18985 3583
rect 18956 2589 18985 2595
rect 19185 3583 19214 3589
rect 19185 2595 19191 3583
rect 19208 2595 19214 3583
rect 19185 2589 19214 2595
rect 19414 3583 19443 3589
rect 19414 2595 19420 3583
rect 19437 2595 19443 3583
rect 19414 2589 19443 2595
rect 19643 3583 19672 3589
rect 19643 2595 19649 3583
rect 19666 2595 19672 3583
rect 19643 2589 19672 2595
rect 19989 3594 20018 3600
rect 19989 2606 19995 3594
rect 20012 2606 20018 3594
rect 19989 2600 20018 2606
rect 20218 3594 20247 3600
rect 20218 2606 20224 3594
rect 20241 2606 20247 3594
rect 20218 2600 20247 2606
rect 20447 3594 20476 3600
rect 20447 2606 20453 3594
rect 20470 2606 20476 3594
rect 20447 2600 20476 2606
rect 20676 3594 20705 3600
rect 20676 2606 20682 3594
rect 20699 2606 20705 3594
rect 20676 2600 20705 2606
rect 20905 3594 20934 3600
rect 20905 2606 20911 3594
rect 20928 2606 20934 3594
rect 20905 2600 20934 2606
rect 21247 3599 21276 3605
rect 21247 2611 21253 3599
rect 21270 2611 21276 3599
rect 21247 2605 21276 2611
rect 21476 3599 21505 3605
rect 21476 2611 21482 3599
rect 21499 2611 21505 3599
rect 21476 2605 21505 2611
rect 21705 3599 21734 3605
rect 21705 2611 21711 3599
rect 21728 2611 21734 3599
rect 21705 2605 21734 2611
rect 21934 3599 21963 3605
rect 21934 2611 21940 3599
rect 21957 2611 21963 3599
rect 21934 2605 21963 2611
rect 22163 3599 22192 3605
rect 22163 2611 22169 3599
rect 22186 2611 22192 3599
rect 22163 2605 22192 2611
rect 22624 3596 22653 3602
rect 22624 2608 22630 3596
rect 22647 2608 22653 3596
rect 22624 2602 22653 2608
rect 22853 3596 22882 3602
rect 22853 2608 22859 3596
rect 22876 2608 22882 3596
rect 22853 2602 22882 2608
rect 23082 3596 23111 3602
rect 23082 2608 23088 3596
rect 23105 2608 23111 3596
rect 23082 2602 23111 2608
rect 23311 3596 23340 3602
rect 23311 2608 23317 3596
rect 23334 2608 23340 3596
rect 23311 2602 23340 2608
rect 23540 3596 23569 3602
rect 23540 2608 23546 3596
rect 23563 2608 23569 3596
rect 23540 2602 23569 2608
rect 24032 3583 24061 3589
rect 24032 2595 24038 3583
rect 24055 2595 24061 3583
rect 24032 2589 24061 2595
rect 24261 3583 24290 3589
rect 24261 2595 24267 3583
rect 24284 2595 24290 3583
rect 24261 2589 24290 2595
rect 24490 3583 24519 3589
rect 24490 2595 24496 3583
rect 24513 2595 24519 3583
rect 24490 2589 24519 2595
rect 24719 3583 24748 3589
rect 24719 2595 24725 3583
rect 24742 2595 24748 3583
rect 24719 2589 24748 2595
rect 24948 3583 24977 3589
rect 24948 2595 24954 3583
rect 24971 2595 24977 3583
rect 24948 2589 24977 2595
rect 25294 3594 25323 3600
rect 25294 2606 25300 3594
rect 25317 2606 25323 3594
rect 25294 2600 25323 2606
rect 25523 3594 25552 3600
rect 25523 2606 25529 3594
rect 25546 2606 25552 3594
rect 25523 2600 25552 2606
rect 25752 3594 25781 3600
rect 25752 2606 25758 3594
rect 25775 2606 25781 3594
rect 25752 2600 25781 2606
rect 25981 3594 26010 3600
rect 25981 2606 25987 3594
rect 26004 2606 26010 3594
rect 25981 2600 26010 2606
rect 26210 3594 26239 3600
rect 26210 2606 26216 3594
rect 26233 2606 26239 3594
rect 26210 2600 26239 2606
rect 26511 3599 26540 3605
rect 26511 2611 26517 3599
rect 26534 2611 26540 3599
rect 26511 2605 26540 2611
rect 26740 3599 26769 3605
rect 26740 2611 26746 3599
rect 26763 2611 26769 3599
rect 26740 2605 26769 2611
rect 26969 3599 26998 3605
rect 26969 2611 26975 3599
rect 26992 2611 26998 3599
rect 26969 2605 26998 2611
rect 27198 3599 27227 3605
rect 27198 2611 27204 3599
rect 27221 2611 27227 3599
rect 27198 2605 27227 2611
rect 27427 3599 27456 3605
rect 27427 2611 27433 3599
rect 27450 2611 27456 3599
rect 27427 2605 27456 2611
rect 27888 3596 27917 3602
rect 27888 2608 27894 3596
rect 27911 2608 27917 3596
rect 27888 2602 27917 2608
rect 28117 3596 28146 3602
rect 28117 2608 28123 3596
rect 28140 2608 28146 3596
rect 28117 2602 28146 2608
rect 28346 3596 28375 3602
rect 28346 2608 28352 3596
rect 28369 2608 28375 3596
rect 28346 2602 28375 2608
rect 28575 3596 28604 3602
rect 28575 2608 28581 3596
rect 28598 2608 28604 3596
rect 28575 2602 28604 2608
rect 28804 3596 28833 3602
rect 28804 2608 28810 3596
rect 28827 2608 28833 3596
rect 28804 2602 28833 2608
rect 29296 3583 29325 3589
rect 29296 2595 29302 3583
rect 29319 2595 29325 3583
rect 29296 2589 29325 2595
rect 29525 3583 29554 3589
rect 29525 2595 29531 3583
rect 29548 2595 29554 3583
rect 29525 2589 29554 2595
rect 29754 3583 29783 3589
rect 29754 2595 29760 3583
rect 29777 2595 29783 3583
rect 29754 2589 29783 2595
rect 29983 3583 30012 3589
rect 29983 2595 29989 3583
rect 30006 2595 30012 3583
rect 29983 2589 30012 2595
rect 30212 3583 30241 3589
rect 30212 2595 30218 3583
rect 30235 2595 30241 3583
rect 30212 2589 30241 2595
rect 30558 3594 30587 3600
rect 30558 2606 30564 3594
rect 30581 2606 30587 3594
rect 30558 2600 30587 2606
rect 30787 3594 30816 3600
rect 30787 2606 30793 3594
rect 30810 2606 30816 3594
rect 30787 2600 30816 2606
rect 31016 3594 31045 3600
rect 31016 2606 31022 3594
rect 31039 2606 31045 3594
rect 31016 2600 31045 2606
rect 31245 3594 31274 3600
rect 31245 2606 31251 3594
rect 31268 2606 31274 3594
rect 31245 2600 31274 2606
rect 31474 3594 31503 3600
rect 31474 2606 31480 3594
rect 31497 2606 31503 3594
rect 31474 2600 31503 2606
<< ndiffc >>
rect 6046 2044 7034 2061
rect 6046 2000 7034 2017
rect 8771 2049 9759 2066
rect 8771 2005 9759 2022
rect 11350 2044 12338 2061
rect 11350 2000 12338 2017
rect 14075 2049 15063 2066
rect 14075 2005 15063 2022
rect 16614 2044 17602 2061
rect 16614 2000 17602 2017
rect 19339 2049 20327 2066
rect 19339 2005 20327 2022
rect 21919 2044 22907 2061
rect 21919 2000 22907 2017
rect 24644 2049 25632 2066
rect 24644 2005 25632 2022
rect 27183 2044 28171 2061
rect 27183 2000 28171 2017
rect 29908 2049 30896 2066
rect 29908 2005 30896 2022
rect 7214 332 7231 1520
rect 7443 332 7460 1520
rect 7672 332 7689 1520
rect 7901 332 7918 1520
rect 8130 332 8147 1520
rect 8359 332 8376 1520
rect 8588 332 8605 1520
rect 8817 332 8834 1520
rect 9046 332 9063 1520
rect 9275 332 9292 1520
rect 9504 332 9521 1520
rect 9733 332 9750 1520
rect 12518 332 12535 1520
rect 12747 332 12764 1520
rect 12976 332 12993 1520
rect 13205 332 13222 1520
rect 13434 332 13451 1520
rect 13663 332 13680 1520
rect 13892 332 13909 1520
rect 14121 332 14138 1520
rect 14350 332 14367 1520
rect 14579 332 14596 1520
rect 14808 332 14825 1520
rect 15037 332 15054 1520
rect 17782 332 17799 1520
rect 18011 332 18028 1520
rect 18240 332 18257 1520
rect 18469 332 18486 1520
rect 18698 332 18715 1520
rect 18927 332 18944 1520
rect 19156 332 19173 1520
rect 19385 332 19402 1520
rect 19614 332 19631 1520
rect 19843 332 19860 1520
rect 20072 332 20089 1520
rect 20301 332 20318 1520
rect 23087 332 23104 1520
rect 23316 332 23333 1520
rect 23545 332 23562 1520
rect 23774 332 23791 1520
rect 24003 332 24020 1520
rect 24232 332 24249 1520
rect 24461 332 24478 1520
rect 24690 332 24707 1520
rect 24919 332 24936 1520
rect 25148 332 25165 1520
rect 25377 332 25394 1520
rect 25606 332 25623 1520
rect 28351 332 28368 1520
rect 28580 332 28597 1520
rect 28809 332 28826 1520
rect 29038 332 29055 1520
rect 29267 332 29284 1520
rect 29496 332 29513 1520
rect 29725 332 29742 1520
rect 29954 332 29971 1520
rect 30183 332 30200 1520
rect 30412 332 30429 1520
rect 30641 332 30658 1520
rect 30870 332 30887 1520
<< pdiffc >>
rect 5380 2611 5397 3599
rect 5609 2611 5626 3599
rect 5838 2611 5855 3599
rect 6067 2611 6084 3599
rect 6296 2611 6313 3599
rect 6757 2608 6774 3596
rect 6986 2608 7003 3596
rect 7215 2608 7232 3596
rect 7444 2608 7461 3596
rect 7673 2608 7690 3596
rect 8165 2595 8182 3583
rect 8394 2595 8411 3583
rect 8623 2595 8640 3583
rect 8852 2595 8869 3583
rect 9081 2595 9098 3583
rect 9427 2606 9444 3594
rect 9656 2606 9673 3594
rect 9885 2606 9902 3594
rect 10114 2606 10131 3594
rect 10343 2606 10360 3594
rect 10684 2611 10701 3599
rect 10913 2611 10930 3599
rect 11142 2611 11159 3599
rect 11371 2611 11388 3599
rect 11600 2611 11617 3599
rect 12061 2608 12078 3596
rect 12290 2608 12307 3596
rect 12519 2608 12536 3596
rect 12748 2608 12765 3596
rect 12977 2608 12994 3596
rect 13469 2595 13486 3583
rect 13698 2595 13715 3583
rect 13927 2595 13944 3583
rect 14156 2595 14173 3583
rect 14385 2595 14402 3583
rect 14731 2606 14748 3594
rect 14960 2606 14977 3594
rect 15189 2606 15206 3594
rect 15418 2606 15435 3594
rect 15647 2606 15664 3594
rect 15948 2611 15965 3599
rect 16177 2611 16194 3599
rect 16406 2611 16423 3599
rect 16635 2611 16652 3599
rect 16864 2611 16881 3599
rect 17325 2608 17342 3596
rect 17554 2608 17571 3596
rect 17783 2608 17800 3596
rect 18012 2608 18029 3596
rect 18241 2608 18258 3596
rect 18733 2595 18750 3583
rect 18962 2595 18979 3583
rect 19191 2595 19208 3583
rect 19420 2595 19437 3583
rect 19649 2595 19666 3583
rect 19995 2606 20012 3594
rect 20224 2606 20241 3594
rect 20453 2606 20470 3594
rect 20682 2606 20699 3594
rect 20911 2606 20928 3594
rect 21253 2611 21270 3599
rect 21482 2611 21499 3599
rect 21711 2611 21728 3599
rect 21940 2611 21957 3599
rect 22169 2611 22186 3599
rect 22630 2608 22647 3596
rect 22859 2608 22876 3596
rect 23088 2608 23105 3596
rect 23317 2608 23334 3596
rect 23546 2608 23563 3596
rect 24038 2595 24055 3583
rect 24267 2595 24284 3583
rect 24496 2595 24513 3583
rect 24725 2595 24742 3583
rect 24954 2595 24971 3583
rect 25300 2606 25317 3594
rect 25529 2606 25546 3594
rect 25758 2606 25775 3594
rect 25987 2606 26004 3594
rect 26216 2606 26233 3594
rect 26517 2611 26534 3599
rect 26746 2611 26763 3599
rect 26975 2611 26992 3599
rect 27204 2611 27221 3599
rect 27433 2611 27450 3599
rect 27894 2608 27911 3596
rect 28123 2608 28140 3596
rect 28352 2608 28369 3596
rect 28581 2608 28598 3596
rect 28810 2608 28827 3596
rect 29302 2595 29319 3583
rect 29531 2595 29548 3583
rect 29760 2595 29777 3583
rect 29989 2595 30006 3583
rect 30218 2595 30235 3583
rect 30564 2606 30581 3594
rect 30793 2606 30810 3594
rect 31022 2606 31039 3594
rect 31251 2606 31268 3594
rect 31480 2606 31497 3594
<< psubdiff >>
rect 5953 2101 6001 2118
rect 7079 2101 7127 2118
rect 5953 2070 5970 2101
rect 7110 2070 7127 2101
rect 5953 1960 5970 1991
rect 7110 1960 7127 1991
rect 5953 1943 6001 1960
rect 7079 1943 7127 1960
rect 8678 2106 8726 2123
rect 9804 2106 9852 2123
rect 8678 2075 8695 2106
rect 9835 2075 9852 2106
rect 8678 1965 8695 1996
rect 9835 1965 9852 1996
rect 8678 1948 8726 1965
rect 9804 1948 9852 1965
rect 11257 2101 11305 2118
rect 12383 2101 12431 2118
rect 11257 2070 11274 2101
rect 12414 2070 12431 2101
rect 11257 1960 11274 1991
rect 12414 1960 12431 1991
rect 11257 1943 11305 1960
rect 12383 1943 12431 1960
rect 13982 2106 14030 2123
rect 15108 2106 15156 2123
rect 13982 2075 13999 2106
rect 15139 2075 15156 2106
rect 13982 1965 13999 1996
rect 15139 1965 15156 1996
rect 13982 1948 14030 1965
rect 15108 1948 15156 1965
rect 16521 2101 16569 2118
rect 17647 2101 17695 2118
rect 16521 2070 16538 2101
rect 17678 2070 17695 2101
rect 16521 1960 16538 1991
rect 17678 1960 17695 1991
rect 16521 1943 16569 1960
rect 17647 1943 17695 1960
rect 19246 2106 19294 2123
rect 20372 2106 20420 2123
rect 19246 2075 19263 2106
rect 20403 2075 20420 2106
rect 19246 1965 19263 1996
rect 20403 1965 20420 1996
rect 19246 1948 19294 1965
rect 20372 1948 20420 1965
rect 21826 2101 21874 2118
rect 22952 2101 23000 2118
rect 21826 2070 21843 2101
rect 22983 2070 23000 2101
rect 21826 1960 21843 1991
rect 22983 1960 23000 1991
rect 21826 1943 21874 1960
rect 22952 1943 23000 1960
rect 24551 2106 24599 2123
rect 25677 2106 25725 2123
rect 24551 2075 24568 2106
rect 25708 2075 25725 2106
rect 24551 1965 24568 1996
rect 25708 1965 25725 1996
rect 24551 1948 24599 1965
rect 25677 1948 25725 1965
rect 27090 2101 27138 2118
rect 28216 2101 28264 2118
rect 27090 2070 27107 2101
rect 28247 2070 28264 2101
rect 27090 1960 27107 1991
rect 28247 1960 28264 1991
rect 27090 1943 27138 1960
rect 28216 1943 28264 1960
rect 29815 2106 29863 2123
rect 30941 2106 30989 2123
rect 29815 2075 29832 2106
rect 30972 2075 30989 2106
rect 29815 1965 29832 1996
rect 30972 1965 30989 1996
rect 29815 1948 29863 1965
rect 30941 1948 30989 1965
rect 7157 1596 7205 1613
rect 9759 1596 9807 1613
rect 7157 1565 7174 1596
rect 9790 1565 9807 1596
rect 7157 256 7174 287
rect 9790 256 9807 287
rect 7157 239 7205 256
rect 9759 239 9807 256
rect 12461 1596 12509 1613
rect 15063 1596 15111 1613
rect 12461 1565 12478 1596
rect 15094 1565 15111 1596
rect 12461 256 12478 287
rect 15094 256 15111 287
rect 12461 239 12509 256
rect 15063 239 15111 256
rect 17725 1596 17773 1613
rect 20327 1596 20375 1613
rect 17725 1565 17742 1596
rect 20358 1565 20375 1596
rect 17725 256 17742 287
rect 20358 256 20375 287
rect 17725 239 17773 256
rect 20327 239 20375 256
rect 23030 1596 23078 1613
rect 25632 1596 25680 1613
rect 23030 1565 23047 1596
rect 25663 1565 25680 1596
rect 23030 256 23047 287
rect 25663 256 25680 287
rect 23030 239 23078 256
rect 25632 239 25680 256
rect 28294 1596 28342 1613
rect 30896 1596 30944 1613
rect 28294 1565 28311 1596
rect 30927 1565 30944 1596
rect 28294 256 28311 287
rect 30927 256 30944 287
rect 28294 239 28342 256
rect 30896 239 30944 256
rect 7122 134 9888 161
rect 7122 132 9295 134
rect 7122 129 7861 132
rect 7122 71 7414 129
rect 7493 74 7861 129
rect 7940 74 8746 132
rect 8825 76 9295 132
rect 9374 76 9888 134
rect 8825 74 9888 76
rect 7493 71 9888 74
rect 7122 47 9888 71
rect 12426 134 15192 161
rect 12426 132 14599 134
rect 12426 129 13165 132
rect 12426 71 12718 129
rect 12797 74 13165 129
rect 13244 74 14050 132
rect 14129 76 14599 132
rect 14678 76 15192 134
rect 14129 74 15192 76
rect 12797 71 15192 74
rect 12426 47 15192 71
rect 17690 134 20456 161
rect 17690 132 19863 134
rect 17690 129 18429 132
rect 17690 71 17982 129
rect 18061 74 18429 129
rect 18508 74 19314 132
rect 19393 76 19863 132
rect 19942 76 20456 134
rect 19393 74 20456 76
rect 18061 71 20456 74
rect 17690 47 20456 71
rect 22995 134 25761 161
rect 22995 132 25168 134
rect 22995 129 23734 132
rect 22995 71 23287 129
rect 23366 74 23734 129
rect 23813 74 24619 132
rect 24698 76 25168 132
rect 25247 76 25761 134
rect 24698 74 25761 76
rect 23366 71 25761 74
rect 22995 47 25761 71
rect 28259 134 31025 161
rect 28259 132 30432 134
rect 28259 129 28998 132
rect 28259 71 28551 129
rect 28630 74 28998 129
rect 29077 74 29883 132
rect 29962 76 30432 132
rect 30511 76 31025 134
rect 29962 74 31025 76
rect 28630 71 31025 74
rect 28259 47 31025 71
<< nsubdiff >>
rect 9208 3855 10443 3865
rect 14512 3855 15747 3865
rect 19776 3855 21011 3865
rect 25081 3855 26316 3865
rect 30345 3855 31580 3865
rect 7711 3854 10443 3855
rect 13015 3854 15747 3855
rect 18279 3854 21011 3855
rect 23584 3854 26316 3855
rect 28848 3854 31580 3855
rect 5329 3848 10443 3854
rect 5329 3839 8354 3848
rect 5329 3834 6958 3839
rect 5329 3829 6037 3834
rect 5329 3782 5570 3829
rect 5638 3787 6037 3829
rect 6105 3794 6958 3834
rect 7014 3835 8354 3839
rect 7014 3794 7417 3835
rect 6105 3790 7417 3794
rect 7473 3797 8354 3835
rect 8407 3845 10443 3848
rect 8407 3797 8835 3845
rect 7473 3794 8835 3797
rect 8888 3842 10443 3845
rect 8888 3841 10097 3842
rect 8888 3795 9624 3841
rect 9669 3796 10097 3841
rect 10142 3796 10443 3842
rect 9669 3795 10443 3796
rect 8888 3794 10443 3795
rect 7473 3790 10443 3794
rect 6105 3787 10443 3790
rect 5638 3782 10443 3787
rect 5329 3778 10443 3782
rect 5329 3774 6390 3778
rect 7711 3776 10443 3778
rect 9208 3774 10443 3776
rect 10633 3848 15747 3854
rect 10633 3839 13658 3848
rect 10633 3834 12262 3839
rect 10633 3829 11341 3834
rect 10633 3782 10874 3829
rect 10942 3787 11341 3829
rect 11409 3794 12262 3834
rect 12318 3835 13658 3839
rect 12318 3794 12721 3835
rect 11409 3790 12721 3794
rect 12777 3797 13658 3835
rect 13711 3845 15747 3848
rect 13711 3797 14139 3845
rect 12777 3794 14139 3797
rect 14192 3842 15747 3845
rect 14192 3841 15401 3842
rect 14192 3795 14928 3841
rect 14973 3796 15401 3841
rect 15446 3796 15747 3842
rect 14973 3795 15747 3796
rect 14192 3794 15747 3795
rect 12777 3790 15747 3794
rect 11409 3787 15747 3790
rect 10942 3782 15747 3787
rect 10633 3778 15747 3782
rect 10633 3774 11694 3778
rect 13015 3776 15747 3778
rect 14512 3774 15747 3776
rect 15897 3848 21011 3854
rect 15897 3839 18922 3848
rect 15897 3834 17526 3839
rect 15897 3829 16605 3834
rect 15897 3782 16138 3829
rect 16206 3787 16605 3829
rect 16673 3794 17526 3834
rect 17582 3835 18922 3839
rect 17582 3794 17985 3835
rect 16673 3790 17985 3794
rect 18041 3797 18922 3835
rect 18975 3845 21011 3848
rect 18975 3797 19403 3845
rect 18041 3794 19403 3797
rect 19456 3842 21011 3845
rect 19456 3841 20665 3842
rect 19456 3795 20192 3841
rect 20237 3796 20665 3841
rect 20710 3796 21011 3842
rect 20237 3795 21011 3796
rect 19456 3794 21011 3795
rect 18041 3790 21011 3794
rect 16673 3787 21011 3790
rect 16206 3782 21011 3787
rect 15897 3778 21011 3782
rect 15897 3774 16958 3778
rect 18279 3776 21011 3778
rect 19776 3774 21011 3776
rect 21202 3848 26316 3854
rect 21202 3839 24227 3848
rect 21202 3834 22831 3839
rect 21202 3829 21910 3834
rect 21202 3782 21443 3829
rect 21511 3787 21910 3829
rect 21978 3794 22831 3834
rect 22887 3835 24227 3839
rect 22887 3794 23290 3835
rect 21978 3790 23290 3794
rect 23346 3797 24227 3835
rect 24280 3845 26316 3848
rect 24280 3797 24708 3845
rect 23346 3794 24708 3797
rect 24761 3842 26316 3845
rect 24761 3841 25970 3842
rect 24761 3795 25497 3841
rect 25542 3796 25970 3841
rect 26015 3796 26316 3842
rect 25542 3795 26316 3796
rect 24761 3794 26316 3795
rect 23346 3790 26316 3794
rect 21978 3787 26316 3790
rect 21511 3782 26316 3787
rect 21202 3778 26316 3782
rect 21202 3774 22263 3778
rect 23584 3776 26316 3778
rect 25081 3774 26316 3776
rect 26466 3848 31580 3854
rect 26466 3839 29491 3848
rect 26466 3834 28095 3839
rect 26466 3829 27174 3834
rect 26466 3782 26707 3829
rect 26775 3787 27174 3829
rect 27242 3794 28095 3834
rect 28151 3835 29491 3839
rect 28151 3794 28554 3835
rect 27242 3790 28554 3794
rect 28610 3797 29491 3835
rect 29544 3845 31580 3848
rect 29544 3797 29972 3845
rect 28610 3794 29972 3797
rect 30025 3842 31580 3845
rect 30025 3841 31234 3842
rect 30025 3795 30761 3841
rect 30806 3796 31234 3841
rect 31279 3796 31580 3842
rect 30806 3795 31580 3796
rect 30025 3794 31580 3795
rect 28610 3790 31580 3794
rect 27242 3787 31580 3790
rect 26775 3782 31580 3787
rect 26466 3778 31580 3782
rect 26466 3774 27527 3778
rect 28848 3776 31580 3778
rect 30345 3774 31580 3776
rect 5323 3680 5371 3697
rect 6322 3680 6370 3697
rect 5323 3649 5340 3680
rect 6353 3649 6370 3680
rect 5323 2531 5340 2562
rect 6353 2531 6370 2562
rect 5323 2514 5371 2531
rect 6322 2514 6370 2531
rect 6700 3677 6748 3694
rect 7699 3677 7747 3694
rect 6700 3646 6717 3677
rect 7730 3646 7747 3677
rect 6700 2528 6717 2559
rect 7730 2528 7747 2559
rect 6700 2511 6748 2528
rect 7699 2511 7747 2528
rect 8108 3664 8156 3681
rect 9107 3664 9155 3681
rect 8108 3633 8125 3664
rect 9138 3633 9155 3664
rect 8108 2515 8125 2546
rect 9138 2515 9155 2546
rect 8108 2498 8156 2515
rect 9107 2498 9155 2515
rect 9370 3675 9418 3692
rect 10369 3675 10417 3692
rect 9370 3644 9387 3675
rect 10400 3644 10417 3675
rect 9370 2526 9387 2557
rect 10400 2526 10417 2557
rect 9370 2509 9418 2526
rect 10369 2509 10417 2526
rect 10627 3680 10675 3697
rect 11626 3680 11674 3697
rect 10627 3649 10644 3680
rect 11657 3649 11674 3680
rect 10627 2531 10644 2562
rect 11657 2531 11674 2562
rect 10627 2514 10675 2531
rect 11626 2514 11674 2531
rect 12004 3677 12052 3694
rect 13003 3677 13051 3694
rect 12004 3646 12021 3677
rect 13034 3646 13051 3677
rect 12004 2528 12021 2559
rect 13034 2528 13051 2559
rect 12004 2511 12052 2528
rect 13003 2511 13051 2528
rect 13412 3664 13460 3681
rect 14411 3664 14459 3681
rect 13412 3633 13429 3664
rect 14442 3633 14459 3664
rect 13412 2515 13429 2546
rect 14442 2515 14459 2546
rect 13412 2498 13460 2515
rect 14411 2498 14459 2515
rect 14674 3675 14722 3692
rect 15673 3675 15721 3692
rect 14674 3644 14691 3675
rect 15704 3644 15721 3675
rect 14674 2526 14691 2557
rect 15704 2526 15721 2557
rect 14674 2509 14722 2526
rect 15673 2509 15721 2526
rect 15891 3680 15939 3697
rect 16890 3680 16938 3697
rect 15891 3649 15908 3680
rect 16921 3649 16938 3680
rect 15891 2531 15908 2562
rect 16921 2531 16938 2562
rect 15891 2514 15939 2531
rect 16890 2514 16938 2531
rect 17268 3677 17316 3694
rect 18267 3677 18315 3694
rect 17268 3646 17285 3677
rect 18298 3646 18315 3677
rect 17268 2528 17285 2559
rect 18298 2528 18315 2559
rect 17268 2511 17316 2528
rect 18267 2511 18315 2528
rect 18676 3664 18724 3681
rect 19675 3664 19723 3681
rect 18676 3633 18693 3664
rect 19706 3633 19723 3664
rect 18676 2515 18693 2546
rect 19706 2515 19723 2546
rect 18676 2498 18724 2515
rect 19675 2498 19723 2515
rect 19938 3675 19986 3692
rect 20937 3675 20985 3692
rect 19938 3644 19955 3675
rect 20968 3644 20985 3675
rect 19938 2526 19955 2557
rect 20968 2526 20985 2557
rect 19938 2509 19986 2526
rect 20937 2509 20985 2526
rect 21196 3680 21244 3697
rect 22195 3680 22243 3697
rect 21196 3649 21213 3680
rect 22226 3649 22243 3680
rect 21196 2531 21213 2562
rect 22226 2531 22243 2562
rect 21196 2514 21244 2531
rect 22195 2514 22243 2531
rect 22573 3677 22621 3694
rect 23572 3677 23620 3694
rect 22573 3646 22590 3677
rect 23603 3646 23620 3677
rect 22573 2528 22590 2559
rect 23603 2528 23620 2559
rect 22573 2511 22621 2528
rect 23572 2511 23620 2528
rect 23981 3664 24029 3681
rect 24980 3664 25028 3681
rect 23981 3633 23998 3664
rect 25011 3633 25028 3664
rect 23981 2515 23998 2546
rect 25011 2515 25028 2546
rect 23981 2498 24029 2515
rect 24980 2498 25028 2515
rect 25243 3675 25291 3692
rect 26242 3675 26290 3692
rect 25243 3644 25260 3675
rect 26273 3644 26290 3675
rect 25243 2526 25260 2557
rect 26273 2526 26290 2557
rect 25243 2509 25291 2526
rect 26242 2509 26290 2526
rect 26460 3680 26508 3697
rect 27459 3680 27507 3697
rect 26460 3649 26477 3680
rect 27490 3649 27507 3680
rect 26460 2531 26477 2562
rect 27490 2531 27507 2562
rect 26460 2514 26508 2531
rect 27459 2514 27507 2531
rect 27837 3677 27885 3694
rect 28836 3677 28884 3694
rect 27837 3646 27854 3677
rect 28867 3646 28884 3677
rect 27837 2528 27854 2559
rect 28867 2528 28884 2559
rect 27837 2511 27885 2528
rect 28836 2511 28884 2528
rect 29245 3664 29293 3681
rect 30244 3664 30292 3681
rect 29245 3633 29262 3664
rect 30275 3633 30292 3664
rect 29245 2515 29262 2546
rect 30275 2515 30292 2546
rect 29245 2498 29293 2515
rect 30244 2498 30292 2515
rect 30507 3675 30555 3692
rect 31506 3675 31554 3692
rect 30507 3644 30524 3675
rect 31537 3644 31554 3675
rect 30507 2526 30524 2557
rect 31537 2526 31554 2557
rect 30507 2509 30555 2526
rect 31506 2509 31554 2526
<< psubdiffcont >>
rect 6001 2101 7079 2118
rect 5953 1991 5970 2070
rect 7110 1991 7127 2070
rect 6001 1943 7079 1960
rect 8726 2106 9804 2123
rect 8678 1996 8695 2075
rect 9835 1996 9852 2075
rect 8726 1948 9804 1965
rect 11305 2101 12383 2118
rect 11257 1991 11274 2070
rect 12414 1991 12431 2070
rect 11305 1943 12383 1960
rect 14030 2106 15108 2123
rect 13982 1996 13999 2075
rect 15139 1996 15156 2075
rect 14030 1948 15108 1965
rect 16569 2101 17647 2118
rect 16521 1991 16538 2070
rect 17678 1991 17695 2070
rect 16569 1943 17647 1960
rect 19294 2106 20372 2123
rect 19246 1996 19263 2075
rect 20403 1996 20420 2075
rect 19294 1948 20372 1965
rect 21874 2101 22952 2118
rect 21826 1991 21843 2070
rect 22983 1991 23000 2070
rect 21874 1943 22952 1960
rect 24599 2106 25677 2123
rect 24551 1996 24568 2075
rect 25708 1996 25725 2075
rect 24599 1948 25677 1965
rect 27138 2101 28216 2118
rect 27090 1991 27107 2070
rect 28247 1991 28264 2070
rect 27138 1943 28216 1960
rect 29863 2106 30941 2123
rect 29815 1996 29832 2075
rect 30972 1996 30989 2075
rect 29863 1948 30941 1965
rect 7205 1596 9759 1613
rect 7157 287 7174 1565
rect 9790 287 9807 1565
rect 7205 239 9759 256
rect 12509 1596 15063 1613
rect 12461 287 12478 1565
rect 15094 287 15111 1565
rect 12509 239 15063 256
rect 17773 1596 20327 1613
rect 17725 287 17742 1565
rect 20358 287 20375 1565
rect 17773 239 20327 256
rect 23078 1596 25632 1613
rect 23030 287 23047 1565
rect 25663 287 25680 1565
rect 23078 239 25632 256
rect 28342 1596 30896 1613
rect 28294 287 28311 1565
rect 30927 287 30944 1565
rect 28342 239 30896 256
rect 7414 71 7493 129
rect 7861 74 7940 132
rect 8746 74 8825 132
rect 9295 76 9374 134
rect 12718 71 12797 129
rect 13165 74 13244 132
rect 14050 74 14129 132
rect 14599 76 14678 134
rect 17982 71 18061 129
rect 18429 74 18508 132
rect 19314 74 19393 132
rect 19863 76 19942 134
rect 23287 71 23366 129
rect 23734 74 23813 132
rect 24619 74 24698 132
rect 25168 76 25247 134
rect 28551 71 28630 129
rect 28998 74 29077 132
rect 29883 74 29962 132
rect 30432 76 30511 134
<< nsubdiffcont >>
rect 5570 3782 5638 3829
rect 6037 3787 6105 3834
rect 6958 3794 7014 3839
rect 7417 3790 7473 3835
rect 8354 3797 8407 3848
rect 8835 3794 8888 3845
rect 9624 3795 9669 3841
rect 10097 3796 10142 3842
rect 10874 3782 10942 3829
rect 11341 3787 11409 3834
rect 12262 3794 12318 3839
rect 12721 3790 12777 3835
rect 13658 3797 13711 3848
rect 14139 3794 14192 3845
rect 14928 3795 14973 3841
rect 15401 3796 15446 3842
rect 16138 3782 16206 3829
rect 16605 3787 16673 3834
rect 17526 3794 17582 3839
rect 17985 3790 18041 3835
rect 18922 3797 18975 3848
rect 19403 3794 19456 3845
rect 20192 3795 20237 3841
rect 20665 3796 20710 3842
rect 21443 3782 21511 3829
rect 21910 3787 21978 3834
rect 22831 3794 22887 3839
rect 23290 3790 23346 3835
rect 24227 3797 24280 3848
rect 24708 3794 24761 3845
rect 25497 3795 25542 3841
rect 25970 3796 26015 3842
rect 26707 3782 26775 3829
rect 27174 3787 27242 3834
rect 28095 3794 28151 3839
rect 28554 3790 28610 3835
rect 29491 3797 29544 3848
rect 29972 3794 30025 3845
rect 30761 3795 30806 3841
rect 31234 3796 31279 3842
rect 5371 3680 6322 3697
rect 5323 2562 5340 3649
rect 6353 2562 6370 3649
rect 5371 2514 6322 2531
rect 6748 3677 7699 3694
rect 6700 2559 6717 3646
rect 7730 2559 7747 3646
rect 6748 2511 7699 2528
rect 8156 3664 9107 3681
rect 8108 2546 8125 3633
rect 9138 2546 9155 3633
rect 8156 2498 9107 2515
rect 9418 3675 10369 3692
rect 9370 2557 9387 3644
rect 10400 2557 10417 3644
rect 9418 2509 10369 2526
rect 10675 3680 11626 3697
rect 10627 2562 10644 3649
rect 11657 2562 11674 3649
rect 10675 2514 11626 2531
rect 12052 3677 13003 3694
rect 12004 2559 12021 3646
rect 13034 2559 13051 3646
rect 12052 2511 13003 2528
rect 13460 3664 14411 3681
rect 13412 2546 13429 3633
rect 14442 2546 14459 3633
rect 13460 2498 14411 2515
rect 14722 3675 15673 3692
rect 14674 2557 14691 3644
rect 15704 2557 15721 3644
rect 14722 2509 15673 2526
rect 15939 3680 16890 3697
rect 15891 2562 15908 3649
rect 16921 2562 16938 3649
rect 15939 2514 16890 2531
rect 17316 3677 18267 3694
rect 17268 2559 17285 3646
rect 18298 2559 18315 3646
rect 17316 2511 18267 2528
rect 18724 3664 19675 3681
rect 18676 2546 18693 3633
rect 19706 2546 19723 3633
rect 18724 2498 19675 2515
rect 19986 3675 20937 3692
rect 19938 2557 19955 3644
rect 20968 2557 20985 3644
rect 19986 2509 20937 2526
rect 21244 3680 22195 3697
rect 21196 2562 21213 3649
rect 22226 2562 22243 3649
rect 21244 2514 22195 2531
rect 22621 3677 23572 3694
rect 22573 2559 22590 3646
rect 23603 2559 23620 3646
rect 22621 2511 23572 2528
rect 24029 3664 24980 3681
rect 23981 2546 23998 3633
rect 25011 2546 25028 3633
rect 24029 2498 24980 2515
rect 25291 3675 26242 3692
rect 25243 2557 25260 3644
rect 26273 2557 26290 3644
rect 25291 2509 26242 2526
rect 26508 3680 27459 3697
rect 26460 2562 26477 3649
rect 27490 2562 27507 3649
rect 26508 2514 27459 2531
rect 27885 3677 28836 3694
rect 27837 2559 27854 3646
rect 28867 2559 28884 3646
rect 27885 2511 28836 2528
rect 29293 3664 30244 3681
rect 29245 2546 29262 3633
rect 30275 2546 30292 3633
rect 29293 2498 30244 2515
rect 30555 3675 31506 3692
rect 30507 2557 30524 3644
rect 31537 2557 31554 3644
rect 30555 2509 31506 2526
<< poly >>
rect 5403 3646 5603 3654
rect 5403 3629 5411 3646
rect 5595 3629 5603 3646
rect 5403 3605 5603 3629
rect 5632 3646 5832 3654
rect 5632 3629 5640 3646
rect 5824 3629 5832 3646
rect 5632 3605 5832 3629
rect 5861 3646 6061 3654
rect 5861 3629 5869 3646
rect 6053 3629 6061 3646
rect 5861 3605 6061 3629
rect 6090 3646 6290 3654
rect 6090 3629 6098 3646
rect 6282 3629 6290 3646
rect 6090 3605 6290 3629
rect 5403 2582 5603 2605
rect 5403 2565 5411 2582
rect 5595 2565 5603 2582
rect 5403 2557 5603 2565
rect 5632 2582 5832 2605
rect 5632 2565 5640 2582
rect 5824 2565 5832 2582
rect 5632 2557 5832 2565
rect 5861 2582 6061 2605
rect 5861 2565 5869 2582
rect 6053 2565 6061 2582
rect 5861 2557 6061 2565
rect 6090 2582 6290 2605
rect 6090 2565 6098 2582
rect 6282 2565 6290 2582
rect 6090 2557 6290 2565
rect 6780 3643 6980 3651
rect 6780 3626 6788 3643
rect 6972 3626 6980 3643
rect 6780 3602 6980 3626
rect 7009 3643 7209 3651
rect 7009 3626 7017 3643
rect 7201 3626 7209 3643
rect 7009 3602 7209 3626
rect 7238 3643 7438 3651
rect 7238 3626 7246 3643
rect 7430 3626 7438 3643
rect 7238 3602 7438 3626
rect 7467 3643 7667 3651
rect 7467 3626 7475 3643
rect 7659 3626 7667 3643
rect 7467 3602 7667 3626
rect 6780 2579 6980 2602
rect 6780 2562 6788 2579
rect 6972 2562 6980 2579
rect 6780 2554 6980 2562
rect 7009 2579 7209 2602
rect 7009 2562 7017 2579
rect 7201 2562 7209 2579
rect 7009 2554 7209 2562
rect 7238 2579 7438 2602
rect 7238 2562 7246 2579
rect 7430 2562 7438 2579
rect 7238 2554 7438 2562
rect 7467 2579 7667 2602
rect 7467 2562 7475 2579
rect 7659 2562 7667 2579
rect 7467 2554 7667 2562
rect 8188 3630 8388 3638
rect 8188 3613 8196 3630
rect 8380 3613 8388 3630
rect 8188 3589 8388 3613
rect 8417 3630 8617 3638
rect 8417 3613 8425 3630
rect 8609 3613 8617 3630
rect 8417 3589 8617 3613
rect 8646 3630 8846 3638
rect 8646 3613 8654 3630
rect 8838 3613 8846 3630
rect 8646 3589 8846 3613
rect 8875 3630 9075 3638
rect 8875 3613 8883 3630
rect 9067 3613 9075 3630
rect 8875 3589 9075 3613
rect 8188 2566 8388 2589
rect 8188 2549 8196 2566
rect 8380 2549 8388 2566
rect 8188 2541 8388 2549
rect 8417 2566 8617 2589
rect 8417 2549 8425 2566
rect 8609 2549 8617 2566
rect 8417 2541 8617 2549
rect 8646 2566 8846 2589
rect 8646 2549 8654 2566
rect 8838 2549 8846 2566
rect 8646 2541 8846 2549
rect 8875 2566 9075 2589
rect 8875 2549 8883 2566
rect 9067 2549 9075 2566
rect 8875 2541 9075 2549
rect 9450 3641 9650 3649
rect 9450 3624 9458 3641
rect 9642 3624 9650 3641
rect 9450 3600 9650 3624
rect 9679 3641 9879 3649
rect 9679 3624 9687 3641
rect 9871 3624 9879 3641
rect 9679 3600 9879 3624
rect 9908 3641 10108 3649
rect 9908 3624 9916 3641
rect 10100 3624 10108 3641
rect 9908 3600 10108 3624
rect 10137 3641 10337 3649
rect 10137 3624 10145 3641
rect 10329 3624 10337 3641
rect 10137 3600 10337 3624
rect 9450 2577 9650 2600
rect 9450 2560 9458 2577
rect 9642 2560 9650 2577
rect 9450 2552 9650 2560
rect 9679 2577 9879 2600
rect 9679 2560 9687 2577
rect 9871 2560 9879 2577
rect 9679 2552 9879 2560
rect 9908 2577 10108 2600
rect 9908 2560 9916 2577
rect 10100 2560 10108 2577
rect 9908 2552 10108 2560
rect 10137 2577 10337 2600
rect 10137 2560 10145 2577
rect 10329 2560 10337 2577
rect 10137 2552 10337 2560
rect 10707 3646 10907 3654
rect 10707 3629 10715 3646
rect 10899 3629 10907 3646
rect 10707 3605 10907 3629
rect 10936 3646 11136 3654
rect 10936 3629 10944 3646
rect 11128 3629 11136 3646
rect 10936 3605 11136 3629
rect 11165 3646 11365 3654
rect 11165 3629 11173 3646
rect 11357 3629 11365 3646
rect 11165 3605 11365 3629
rect 11394 3646 11594 3654
rect 11394 3629 11402 3646
rect 11586 3629 11594 3646
rect 11394 3605 11594 3629
rect 10707 2582 10907 2605
rect 10707 2565 10715 2582
rect 10899 2565 10907 2582
rect 10707 2557 10907 2565
rect 10936 2582 11136 2605
rect 10936 2565 10944 2582
rect 11128 2565 11136 2582
rect 10936 2557 11136 2565
rect 11165 2582 11365 2605
rect 11165 2565 11173 2582
rect 11357 2565 11365 2582
rect 11165 2557 11365 2565
rect 11394 2582 11594 2605
rect 11394 2565 11402 2582
rect 11586 2565 11594 2582
rect 11394 2557 11594 2565
rect 12084 3643 12284 3651
rect 12084 3626 12092 3643
rect 12276 3626 12284 3643
rect 12084 3602 12284 3626
rect 12313 3643 12513 3651
rect 12313 3626 12321 3643
rect 12505 3626 12513 3643
rect 12313 3602 12513 3626
rect 12542 3643 12742 3651
rect 12542 3626 12550 3643
rect 12734 3626 12742 3643
rect 12542 3602 12742 3626
rect 12771 3643 12971 3651
rect 12771 3626 12779 3643
rect 12963 3626 12971 3643
rect 12771 3602 12971 3626
rect 12084 2579 12284 2602
rect 12084 2562 12092 2579
rect 12276 2562 12284 2579
rect 12084 2554 12284 2562
rect 12313 2579 12513 2602
rect 12313 2562 12321 2579
rect 12505 2562 12513 2579
rect 12313 2554 12513 2562
rect 12542 2579 12742 2602
rect 12542 2562 12550 2579
rect 12734 2562 12742 2579
rect 12542 2554 12742 2562
rect 12771 2579 12971 2602
rect 12771 2562 12779 2579
rect 12963 2562 12971 2579
rect 12771 2554 12971 2562
rect 13492 3630 13692 3638
rect 13492 3613 13500 3630
rect 13684 3613 13692 3630
rect 13492 3589 13692 3613
rect 13721 3630 13921 3638
rect 13721 3613 13729 3630
rect 13913 3613 13921 3630
rect 13721 3589 13921 3613
rect 13950 3630 14150 3638
rect 13950 3613 13958 3630
rect 14142 3613 14150 3630
rect 13950 3589 14150 3613
rect 14179 3630 14379 3638
rect 14179 3613 14187 3630
rect 14371 3613 14379 3630
rect 14179 3589 14379 3613
rect 13492 2566 13692 2589
rect 13492 2549 13500 2566
rect 13684 2549 13692 2566
rect 13492 2541 13692 2549
rect 13721 2566 13921 2589
rect 13721 2549 13729 2566
rect 13913 2549 13921 2566
rect 13721 2541 13921 2549
rect 13950 2566 14150 2589
rect 13950 2549 13958 2566
rect 14142 2549 14150 2566
rect 13950 2541 14150 2549
rect 14179 2566 14379 2589
rect 14179 2549 14187 2566
rect 14371 2549 14379 2566
rect 14179 2541 14379 2549
rect 14754 3641 14954 3649
rect 14754 3624 14762 3641
rect 14946 3624 14954 3641
rect 14754 3600 14954 3624
rect 14983 3641 15183 3649
rect 14983 3624 14991 3641
rect 15175 3624 15183 3641
rect 14983 3600 15183 3624
rect 15212 3641 15412 3649
rect 15212 3624 15220 3641
rect 15404 3624 15412 3641
rect 15212 3600 15412 3624
rect 15441 3641 15641 3649
rect 15441 3624 15449 3641
rect 15633 3624 15641 3641
rect 15441 3600 15641 3624
rect 14754 2577 14954 2600
rect 14754 2560 14762 2577
rect 14946 2560 14954 2577
rect 14754 2552 14954 2560
rect 14983 2577 15183 2600
rect 14983 2560 14991 2577
rect 15175 2560 15183 2577
rect 14983 2552 15183 2560
rect 15212 2577 15412 2600
rect 15212 2560 15220 2577
rect 15404 2560 15412 2577
rect 15212 2552 15412 2560
rect 15441 2577 15641 2600
rect 15441 2560 15449 2577
rect 15633 2560 15641 2577
rect 15441 2552 15641 2560
rect 15971 3646 16171 3654
rect 15971 3629 15979 3646
rect 16163 3629 16171 3646
rect 15971 3605 16171 3629
rect 16200 3646 16400 3654
rect 16200 3629 16208 3646
rect 16392 3629 16400 3646
rect 16200 3605 16400 3629
rect 16429 3646 16629 3654
rect 16429 3629 16437 3646
rect 16621 3629 16629 3646
rect 16429 3605 16629 3629
rect 16658 3646 16858 3654
rect 16658 3629 16666 3646
rect 16850 3629 16858 3646
rect 16658 3605 16858 3629
rect 15971 2582 16171 2605
rect 15971 2565 15979 2582
rect 16163 2565 16171 2582
rect 15971 2557 16171 2565
rect 16200 2582 16400 2605
rect 16200 2565 16208 2582
rect 16392 2565 16400 2582
rect 16200 2557 16400 2565
rect 16429 2582 16629 2605
rect 16429 2565 16437 2582
rect 16621 2565 16629 2582
rect 16429 2557 16629 2565
rect 16658 2582 16858 2605
rect 16658 2565 16666 2582
rect 16850 2565 16858 2582
rect 16658 2557 16858 2565
rect 17348 3643 17548 3651
rect 17348 3626 17356 3643
rect 17540 3626 17548 3643
rect 17348 3602 17548 3626
rect 17577 3643 17777 3651
rect 17577 3626 17585 3643
rect 17769 3626 17777 3643
rect 17577 3602 17777 3626
rect 17806 3643 18006 3651
rect 17806 3626 17814 3643
rect 17998 3626 18006 3643
rect 17806 3602 18006 3626
rect 18035 3643 18235 3651
rect 18035 3626 18043 3643
rect 18227 3626 18235 3643
rect 18035 3602 18235 3626
rect 17348 2579 17548 2602
rect 17348 2562 17356 2579
rect 17540 2562 17548 2579
rect 17348 2554 17548 2562
rect 17577 2579 17777 2602
rect 17577 2562 17585 2579
rect 17769 2562 17777 2579
rect 17577 2554 17777 2562
rect 17806 2579 18006 2602
rect 17806 2562 17814 2579
rect 17998 2562 18006 2579
rect 17806 2554 18006 2562
rect 18035 2579 18235 2602
rect 18035 2562 18043 2579
rect 18227 2562 18235 2579
rect 18035 2554 18235 2562
rect 18756 3630 18956 3638
rect 18756 3613 18764 3630
rect 18948 3613 18956 3630
rect 18756 3589 18956 3613
rect 18985 3630 19185 3638
rect 18985 3613 18993 3630
rect 19177 3613 19185 3630
rect 18985 3589 19185 3613
rect 19214 3630 19414 3638
rect 19214 3613 19222 3630
rect 19406 3613 19414 3630
rect 19214 3589 19414 3613
rect 19443 3630 19643 3638
rect 19443 3613 19451 3630
rect 19635 3613 19643 3630
rect 19443 3589 19643 3613
rect 18756 2566 18956 2589
rect 18756 2549 18764 2566
rect 18948 2549 18956 2566
rect 18756 2541 18956 2549
rect 18985 2566 19185 2589
rect 18985 2549 18993 2566
rect 19177 2549 19185 2566
rect 18985 2541 19185 2549
rect 19214 2566 19414 2589
rect 19214 2549 19222 2566
rect 19406 2549 19414 2566
rect 19214 2541 19414 2549
rect 19443 2566 19643 2589
rect 19443 2549 19451 2566
rect 19635 2549 19643 2566
rect 19443 2541 19643 2549
rect 20018 3641 20218 3649
rect 20018 3624 20026 3641
rect 20210 3624 20218 3641
rect 20018 3600 20218 3624
rect 20247 3641 20447 3649
rect 20247 3624 20255 3641
rect 20439 3624 20447 3641
rect 20247 3600 20447 3624
rect 20476 3641 20676 3649
rect 20476 3624 20484 3641
rect 20668 3624 20676 3641
rect 20476 3600 20676 3624
rect 20705 3641 20905 3649
rect 20705 3624 20713 3641
rect 20897 3624 20905 3641
rect 20705 3600 20905 3624
rect 20018 2577 20218 2600
rect 20018 2560 20026 2577
rect 20210 2560 20218 2577
rect 20018 2552 20218 2560
rect 20247 2577 20447 2600
rect 20247 2560 20255 2577
rect 20439 2560 20447 2577
rect 20247 2552 20447 2560
rect 20476 2577 20676 2600
rect 20476 2560 20484 2577
rect 20668 2560 20676 2577
rect 20476 2552 20676 2560
rect 20705 2577 20905 2600
rect 20705 2560 20713 2577
rect 20897 2560 20905 2577
rect 20705 2552 20905 2560
rect 21276 3646 21476 3654
rect 21276 3629 21284 3646
rect 21468 3629 21476 3646
rect 21276 3605 21476 3629
rect 21505 3646 21705 3654
rect 21505 3629 21513 3646
rect 21697 3629 21705 3646
rect 21505 3605 21705 3629
rect 21734 3646 21934 3654
rect 21734 3629 21742 3646
rect 21926 3629 21934 3646
rect 21734 3605 21934 3629
rect 21963 3646 22163 3654
rect 21963 3629 21971 3646
rect 22155 3629 22163 3646
rect 21963 3605 22163 3629
rect 21276 2582 21476 2605
rect 21276 2565 21284 2582
rect 21468 2565 21476 2582
rect 21276 2557 21476 2565
rect 21505 2582 21705 2605
rect 21505 2565 21513 2582
rect 21697 2565 21705 2582
rect 21505 2557 21705 2565
rect 21734 2582 21934 2605
rect 21734 2565 21742 2582
rect 21926 2565 21934 2582
rect 21734 2557 21934 2565
rect 21963 2582 22163 2605
rect 21963 2565 21971 2582
rect 22155 2565 22163 2582
rect 21963 2557 22163 2565
rect 22653 3643 22853 3651
rect 22653 3626 22661 3643
rect 22845 3626 22853 3643
rect 22653 3602 22853 3626
rect 22882 3643 23082 3651
rect 22882 3626 22890 3643
rect 23074 3626 23082 3643
rect 22882 3602 23082 3626
rect 23111 3643 23311 3651
rect 23111 3626 23119 3643
rect 23303 3626 23311 3643
rect 23111 3602 23311 3626
rect 23340 3643 23540 3651
rect 23340 3626 23348 3643
rect 23532 3626 23540 3643
rect 23340 3602 23540 3626
rect 22653 2579 22853 2602
rect 22653 2562 22661 2579
rect 22845 2562 22853 2579
rect 22653 2554 22853 2562
rect 22882 2579 23082 2602
rect 22882 2562 22890 2579
rect 23074 2562 23082 2579
rect 22882 2554 23082 2562
rect 23111 2579 23311 2602
rect 23111 2562 23119 2579
rect 23303 2562 23311 2579
rect 23111 2554 23311 2562
rect 23340 2579 23540 2602
rect 23340 2562 23348 2579
rect 23532 2562 23540 2579
rect 23340 2554 23540 2562
rect 24061 3630 24261 3638
rect 24061 3613 24069 3630
rect 24253 3613 24261 3630
rect 24061 3589 24261 3613
rect 24290 3630 24490 3638
rect 24290 3613 24298 3630
rect 24482 3613 24490 3630
rect 24290 3589 24490 3613
rect 24519 3630 24719 3638
rect 24519 3613 24527 3630
rect 24711 3613 24719 3630
rect 24519 3589 24719 3613
rect 24748 3630 24948 3638
rect 24748 3613 24756 3630
rect 24940 3613 24948 3630
rect 24748 3589 24948 3613
rect 24061 2566 24261 2589
rect 24061 2549 24069 2566
rect 24253 2549 24261 2566
rect 24061 2541 24261 2549
rect 24290 2566 24490 2589
rect 24290 2549 24298 2566
rect 24482 2549 24490 2566
rect 24290 2541 24490 2549
rect 24519 2566 24719 2589
rect 24519 2549 24527 2566
rect 24711 2549 24719 2566
rect 24519 2541 24719 2549
rect 24748 2566 24948 2589
rect 24748 2549 24756 2566
rect 24940 2549 24948 2566
rect 24748 2541 24948 2549
rect 25323 3641 25523 3649
rect 25323 3624 25331 3641
rect 25515 3624 25523 3641
rect 25323 3600 25523 3624
rect 25552 3641 25752 3649
rect 25552 3624 25560 3641
rect 25744 3624 25752 3641
rect 25552 3600 25752 3624
rect 25781 3641 25981 3649
rect 25781 3624 25789 3641
rect 25973 3624 25981 3641
rect 25781 3600 25981 3624
rect 26010 3641 26210 3649
rect 26010 3624 26018 3641
rect 26202 3624 26210 3641
rect 26010 3600 26210 3624
rect 25323 2577 25523 2600
rect 25323 2560 25331 2577
rect 25515 2560 25523 2577
rect 25323 2552 25523 2560
rect 25552 2577 25752 2600
rect 25552 2560 25560 2577
rect 25744 2560 25752 2577
rect 25552 2552 25752 2560
rect 25781 2577 25981 2600
rect 25781 2560 25789 2577
rect 25973 2560 25981 2577
rect 25781 2552 25981 2560
rect 26010 2577 26210 2600
rect 26010 2560 26018 2577
rect 26202 2560 26210 2577
rect 26010 2552 26210 2560
rect 26540 3646 26740 3654
rect 26540 3629 26548 3646
rect 26732 3629 26740 3646
rect 26540 3605 26740 3629
rect 26769 3646 26969 3654
rect 26769 3629 26777 3646
rect 26961 3629 26969 3646
rect 26769 3605 26969 3629
rect 26998 3646 27198 3654
rect 26998 3629 27006 3646
rect 27190 3629 27198 3646
rect 26998 3605 27198 3629
rect 27227 3646 27427 3654
rect 27227 3629 27235 3646
rect 27419 3629 27427 3646
rect 27227 3605 27427 3629
rect 26540 2582 26740 2605
rect 26540 2565 26548 2582
rect 26732 2565 26740 2582
rect 26540 2557 26740 2565
rect 26769 2582 26969 2605
rect 26769 2565 26777 2582
rect 26961 2565 26969 2582
rect 26769 2557 26969 2565
rect 26998 2582 27198 2605
rect 26998 2565 27006 2582
rect 27190 2565 27198 2582
rect 26998 2557 27198 2565
rect 27227 2582 27427 2605
rect 27227 2565 27235 2582
rect 27419 2565 27427 2582
rect 27227 2557 27427 2565
rect 27917 3643 28117 3651
rect 27917 3626 27925 3643
rect 28109 3626 28117 3643
rect 27917 3602 28117 3626
rect 28146 3643 28346 3651
rect 28146 3626 28154 3643
rect 28338 3626 28346 3643
rect 28146 3602 28346 3626
rect 28375 3643 28575 3651
rect 28375 3626 28383 3643
rect 28567 3626 28575 3643
rect 28375 3602 28575 3626
rect 28604 3643 28804 3651
rect 28604 3626 28612 3643
rect 28796 3626 28804 3643
rect 28604 3602 28804 3626
rect 27917 2579 28117 2602
rect 27917 2562 27925 2579
rect 28109 2562 28117 2579
rect 27917 2554 28117 2562
rect 28146 2579 28346 2602
rect 28146 2562 28154 2579
rect 28338 2562 28346 2579
rect 28146 2554 28346 2562
rect 28375 2579 28575 2602
rect 28375 2562 28383 2579
rect 28567 2562 28575 2579
rect 28375 2554 28575 2562
rect 28604 2579 28804 2602
rect 28604 2562 28612 2579
rect 28796 2562 28804 2579
rect 28604 2554 28804 2562
rect 29325 3630 29525 3638
rect 29325 3613 29333 3630
rect 29517 3613 29525 3630
rect 29325 3589 29525 3613
rect 29554 3630 29754 3638
rect 29554 3613 29562 3630
rect 29746 3613 29754 3630
rect 29554 3589 29754 3613
rect 29783 3630 29983 3638
rect 29783 3613 29791 3630
rect 29975 3613 29983 3630
rect 29783 3589 29983 3613
rect 30012 3630 30212 3638
rect 30012 3613 30020 3630
rect 30204 3613 30212 3630
rect 30012 3589 30212 3613
rect 29325 2566 29525 2589
rect 29325 2549 29333 2566
rect 29517 2549 29525 2566
rect 29325 2541 29525 2549
rect 29554 2566 29754 2589
rect 29554 2549 29562 2566
rect 29746 2549 29754 2566
rect 29554 2541 29754 2549
rect 29783 2566 29983 2589
rect 29783 2549 29791 2566
rect 29975 2549 29983 2566
rect 29783 2541 29983 2549
rect 30012 2566 30212 2589
rect 30012 2549 30020 2566
rect 30204 2549 30212 2566
rect 30012 2541 30212 2549
rect 30587 3641 30787 3649
rect 30587 3624 30595 3641
rect 30779 3624 30787 3641
rect 30587 3600 30787 3624
rect 30816 3641 31016 3649
rect 30816 3624 30824 3641
rect 31008 3624 31016 3641
rect 30816 3600 31016 3624
rect 31045 3641 31245 3649
rect 31045 3624 31053 3641
rect 31237 3624 31245 3641
rect 31045 3600 31245 3624
rect 31274 3641 31474 3649
rect 31274 3624 31282 3641
rect 31466 3624 31474 3641
rect 31274 3600 31474 3624
rect 30587 2577 30787 2600
rect 30587 2560 30595 2577
rect 30779 2560 30787 2577
rect 30587 2552 30787 2560
rect 30816 2577 31016 2600
rect 30816 2560 30824 2577
rect 31008 2560 31016 2577
rect 30816 2552 31016 2560
rect 31045 2577 31245 2600
rect 31045 2560 31053 2577
rect 31237 2560 31245 2577
rect 31045 2552 31245 2560
rect 31274 2577 31474 2600
rect 31274 2560 31282 2577
rect 31466 2560 31474 2577
rect 31274 2552 31474 2560
rect 5996 2039 6029 2047
rect 5996 2022 6004 2039
rect 6021 2038 6029 2039
rect 7051 2039 7084 2047
rect 7051 2038 7059 2039
rect 6021 2023 6040 2038
rect 7040 2023 7059 2038
rect 6021 2022 6029 2023
rect 5996 2014 6029 2022
rect 7051 2022 7059 2023
rect 7076 2022 7084 2039
rect 7051 2014 7084 2022
rect 8721 2044 8754 2052
rect 8721 2027 8729 2044
rect 8746 2043 8754 2044
rect 9776 2044 9809 2052
rect 9776 2043 9784 2044
rect 8746 2028 8765 2043
rect 9765 2028 9784 2043
rect 8746 2027 8754 2028
rect 8721 2019 8754 2027
rect 9776 2027 9784 2028
rect 9801 2027 9809 2044
rect 9776 2019 9809 2027
rect 11300 2039 11333 2047
rect 11300 2022 11308 2039
rect 11325 2038 11333 2039
rect 12355 2039 12388 2047
rect 12355 2038 12363 2039
rect 11325 2023 11344 2038
rect 12344 2023 12363 2038
rect 11325 2022 11333 2023
rect 11300 2014 11333 2022
rect 12355 2022 12363 2023
rect 12380 2022 12388 2039
rect 12355 2014 12388 2022
rect 14025 2044 14058 2052
rect 14025 2027 14033 2044
rect 14050 2043 14058 2044
rect 15080 2044 15113 2052
rect 15080 2043 15088 2044
rect 14050 2028 14069 2043
rect 15069 2028 15088 2043
rect 14050 2027 14058 2028
rect 14025 2019 14058 2027
rect 15080 2027 15088 2028
rect 15105 2027 15113 2044
rect 15080 2019 15113 2027
rect 16564 2039 16597 2047
rect 16564 2022 16572 2039
rect 16589 2038 16597 2039
rect 17619 2039 17652 2047
rect 17619 2038 17627 2039
rect 16589 2023 16608 2038
rect 17608 2023 17627 2038
rect 16589 2022 16597 2023
rect 16564 2014 16597 2022
rect 17619 2022 17627 2023
rect 17644 2022 17652 2039
rect 17619 2014 17652 2022
rect 19289 2044 19322 2052
rect 19289 2027 19297 2044
rect 19314 2043 19322 2044
rect 20344 2044 20377 2052
rect 20344 2043 20352 2044
rect 19314 2028 19333 2043
rect 20333 2028 20352 2043
rect 19314 2027 19322 2028
rect 19289 2019 19322 2027
rect 20344 2027 20352 2028
rect 20369 2027 20377 2044
rect 20344 2019 20377 2027
rect 21869 2039 21902 2047
rect 21869 2022 21877 2039
rect 21894 2038 21902 2039
rect 22924 2039 22957 2047
rect 22924 2038 22932 2039
rect 21894 2023 21913 2038
rect 22913 2023 22932 2038
rect 21894 2022 21902 2023
rect 21869 2014 21902 2022
rect 22924 2022 22932 2023
rect 22949 2022 22957 2039
rect 22924 2014 22957 2022
rect 24594 2044 24627 2052
rect 24594 2027 24602 2044
rect 24619 2043 24627 2044
rect 25649 2044 25682 2052
rect 25649 2043 25657 2044
rect 24619 2028 24638 2043
rect 25638 2028 25657 2043
rect 24619 2027 24627 2028
rect 24594 2019 24627 2027
rect 25649 2027 25657 2028
rect 25674 2027 25682 2044
rect 25649 2019 25682 2027
rect 27133 2039 27166 2047
rect 27133 2022 27141 2039
rect 27158 2038 27166 2039
rect 28188 2039 28221 2047
rect 28188 2038 28196 2039
rect 27158 2023 27177 2038
rect 28177 2023 28196 2038
rect 27158 2022 27166 2023
rect 27133 2014 27166 2022
rect 28188 2022 28196 2023
rect 28213 2022 28221 2039
rect 28188 2014 28221 2022
rect 29858 2044 29891 2052
rect 29858 2027 29866 2044
rect 29883 2043 29891 2044
rect 30913 2044 30946 2052
rect 30913 2043 30921 2044
rect 29883 2028 29902 2043
rect 30902 2028 30921 2043
rect 29883 2027 29891 2028
rect 29858 2019 29891 2027
rect 30913 2027 30921 2028
rect 30938 2027 30946 2044
rect 30913 2019 30946 2027
rect 7237 1562 7437 1570
rect 7237 1545 7245 1562
rect 7429 1545 7437 1562
rect 7237 1526 7437 1545
rect 7466 1562 7666 1570
rect 7466 1545 7474 1562
rect 7658 1545 7666 1562
rect 7466 1526 7666 1545
rect 7695 1562 7895 1570
rect 7695 1545 7703 1562
rect 7887 1545 7895 1562
rect 7695 1526 7895 1545
rect 7924 1562 8124 1570
rect 7924 1545 7932 1562
rect 8116 1545 8124 1562
rect 7924 1526 8124 1545
rect 8153 1562 8353 1570
rect 8153 1545 8161 1562
rect 8345 1545 8353 1562
rect 8153 1526 8353 1545
rect 8382 1562 8582 1570
rect 8382 1545 8390 1562
rect 8574 1545 8582 1562
rect 8382 1526 8582 1545
rect 8611 1562 8811 1570
rect 8611 1545 8619 1562
rect 8803 1545 8811 1562
rect 8611 1526 8811 1545
rect 8840 1562 9040 1570
rect 8840 1545 8848 1562
rect 9032 1545 9040 1562
rect 8840 1526 9040 1545
rect 9069 1562 9269 1570
rect 9069 1545 9077 1562
rect 9261 1545 9269 1562
rect 9069 1526 9269 1545
rect 9298 1562 9498 1570
rect 9298 1545 9306 1562
rect 9490 1545 9498 1562
rect 9298 1526 9498 1545
rect 9527 1562 9727 1570
rect 9527 1545 9535 1562
rect 9719 1545 9727 1562
rect 9527 1526 9727 1545
rect 7237 307 7437 326
rect 7237 290 7245 307
rect 7429 290 7437 307
rect 7237 282 7437 290
rect 7466 307 7666 326
rect 7466 290 7474 307
rect 7658 290 7666 307
rect 7466 282 7666 290
rect 7695 307 7895 326
rect 7695 290 7703 307
rect 7887 290 7895 307
rect 7695 282 7895 290
rect 7924 307 8124 326
rect 7924 290 7932 307
rect 8116 290 8124 307
rect 7924 282 8124 290
rect 8153 307 8353 326
rect 8153 290 8161 307
rect 8345 290 8353 307
rect 8153 282 8353 290
rect 8382 307 8582 326
rect 8382 290 8390 307
rect 8574 290 8582 307
rect 8382 282 8582 290
rect 8611 307 8811 326
rect 8611 290 8619 307
rect 8803 290 8811 307
rect 8611 282 8811 290
rect 8840 307 9040 326
rect 8840 290 8848 307
rect 9032 290 9040 307
rect 8840 282 9040 290
rect 9069 307 9269 326
rect 9069 290 9077 307
rect 9261 290 9269 307
rect 9069 282 9269 290
rect 9298 307 9498 326
rect 9298 290 9306 307
rect 9490 290 9498 307
rect 9298 282 9498 290
rect 9527 307 9727 326
rect 9527 290 9535 307
rect 9719 290 9727 307
rect 9527 282 9727 290
rect 12541 1562 12741 1570
rect 12541 1545 12549 1562
rect 12733 1545 12741 1562
rect 12541 1526 12741 1545
rect 12770 1562 12970 1570
rect 12770 1545 12778 1562
rect 12962 1545 12970 1562
rect 12770 1526 12970 1545
rect 12999 1562 13199 1570
rect 12999 1545 13007 1562
rect 13191 1545 13199 1562
rect 12999 1526 13199 1545
rect 13228 1562 13428 1570
rect 13228 1545 13236 1562
rect 13420 1545 13428 1562
rect 13228 1526 13428 1545
rect 13457 1562 13657 1570
rect 13457 1545 13465 1562
rect 13649 1545 13657 1562
rect 13457 1526 13657 1545
rect 13686 1562 13886 1570
rect 13686 1545 13694 1562
rect 13878 1545 13886 1562
rect 13686 1526 13886 1545
rect 13915 1562 14115 1570
rect 13915 1545 13923 1562
rect 14107 1545 14115 1562
rect 13915 1526 14115 1545
rect 14144 1562 14344 1570
rect 14144 1545 14152 1562
rect 14336 1545 14344 1562
rect 14144 1526 14344 1545
rect 14373 1562 14573 1570
rect 14373 1545 14381 1562
rect 14565 1545 14573 1562
rect 14373 1526 14573 1545
rect 14602 1562 14802 1570
rect 14602 1545 14610 1562
rect 14794 1545 14802 1562
rect 14602 1526 14802 1545
rect 14831 1562 15031 1570
rect 14831 1545 14839 1562
rect 15023 1545 15031 1562
rect 14831 1526 15031 1545
rect 12541 307 12741 326
rect 12541 290 12549 307
rect 12733 290 12741 307
rect 12541 282 12741 290
rect 12770 307 12970 326
rect 12770 290 12778 307
rect 12962 290 12970 307
rect 12770 282 12970 290
rect 12999 307 13199 326
rect 12999 290 13007 307
rect 13191 290 13199 307
rect 12999 282 13199 290
rect 13228 307 13428 326
rect 13228 290 13236 307
rect 13420 290 13428 307
rect 13228 282 13428 290
rect 13457 307 13657 326
rect 13457 290 13465 307
rect 13649 290 13657 307
rect 13457 282 13657 290
rect 13686 307 13886 326
rect 13686 290 13694 307
rect 13878 290 13886 307
rect 13686 282 13886 290
rect 13915 307 14115 326
rect 13915 290 13923 307
rect 14107 290 14115 307
rect 13915 282 14115 290
rect 14144 307 14344 326
rect 14144 290 14152 307
rect 14336 290 14344 307
rect 14144 282 14344 290
rect 14373 307 14573 326
rect 14373 290 14381 307
rect 14565 290 14573 307
rect 14373 282 14573 290
rect 14602 307 14802 326
rect 14602 290 14610 307
rect 14794 290 14802 307
rect 14602 282 14802 290
rect 14831 307 15031 326
rect 14831 290 14839 307
rect 15023 290 15031 307
rect 14831 282 15031 290
rect 17805 1562 18005 1570
rect 17805 1545 17813 1562
rect 17997 1545 18005 1562
rect 17805 1526 18005 1545
rect 18034 1562 18234 1570
rect 18034 1545 18042 1562
rect 18226 1545 18234 1562
rect 18034 1526 18234 1545
rect 18263 1562 18463 1570
rect 18263 1545 18271 1562
rect 18455 1545 18463 1562
rect 18263 1526 18463 1545
rect 18492 1562 18692 1570
rect 18492 1545 18500 1562
rect 18684 1545 18692 1562
rect 18492 1526 18692 1545
rect 18721 1562 18921 1570
rect 18721 1545 18729 1562
rect 18913 1545 18921 1562
rect 18721 1526 18921 1545
rect 18950 1562 19150 1570
rect 18950 1545 18958 1562
rect 19142 1545 19150 1562
rect 18950 1526 19150 1545
rect 19179 1562 19379 1570
rect 19179 1545 19187 1562
rect 19371 1545 19379 1562
rect 19179 1526 19379 1545
rect 19408 1562 19608 1570
rect 19408 1545 19416 1562
rect 19600 1545 19608 1562
rect 19408 1526 19608 1545
rect 19637 1562 19837 1570
rect 19637 1545 19645 1562
rect 19829 1545 19837 1562
rect 19637 1526 19837 1545
rect 19866 1562 20066 1570
rect 19866 1545 19874 1562
rect 20058 1545 20066 1562
rect 19866 1526 20066 1545
rect 20095 1562 20295 1570
rect 20095 1545 20103 1562
rect 20287 1545 20295 1562
rect 20095 1526 20295 1545
rect 17805 307 18005 326
rect 17805 290 17813 307
rect 17997 290 18005 307
rect 17805 282 18005 290
rect 18034 307 18234 326
rect 18034 290 18042 307
rect 18226 290 18234 307
rect 18034 282 18234 290
rect 18263 307 18463 326
rect 18263 290 18271 307
rect 18455 290 18463 307
rect 18263 282 18463 290
rect 18492 307 18692 326
rect 18492 290 18500 307
rect 18684 290 18692 307
rect 18492 282 18692 290
rect 18721 307 18921 326
rect 18721 290 18729 307
rect 18913 290 18921 307
rect 18721 282 18921 290
rect 18950 307 19150 326
rect 18950 290 18958 307
rect 19142 290 19150 307
rect 18950 282 19150 290
rect 19179 307 19379 326
rect 19179 290 19187 307
rect 19371 290 19379 307
rect 19179 282 19379 290
rect 19408 307 19608 326
rect 19408 290 19416 307
rect 19600 290 19608 307
rect 19408 282 19608 290
rect 19637 307 19837 326
rect 19637 290 19645 307
rect 19829 290 19837 307
rect 19637 282 19837 290
rect 19866 307 20066 326
rect 19866 290 19874 307
rect 20058 290 20066 307
rect 19866 282 20066 290
rect 20095 307 20295 326
rect 20095 290 20103 307
rect 20287 290 20295 307
rect 20095 282 20295 290
rect 23110 1562 23310 1570
rect 23110 1545 23118 1562
rect 23302 1545 23310 1562
rect 23110 1526 23310 1545
rect 23339 1562 23539 1570
rect 23339 1545 23347 1562
rect 23531 1545 23539 1562
rect 23339 1526 23539 1545
rect 23568 1562 23768 1570
rect 23568 1545 23576 1562
rect 23760 1545 23768 1562
rect 23568 1526 23768 1545
rect 23797 1562 23997 1570
rect 23797 1545 23805 1562
rect 23989 1545 23997 1562
rect 23797 1526 23997 1545
rect 24026 1562 24226 1570
rect 24026 1545 24034 1562
rect 24218 1545 24226 1562
rect 24026 1526 24226 1545
rect 24255 1562 24455 1570
rect 24255 1545 24263 1562
rect 24447 1545 24455 1562
rect 24255 1526 24455 1545
rect 24484 1562 24684 1570
rect 24484 1545 24492 1562
rect 24676 1545 24684 1562
rect 24484 1526 24684 1545
rect 24713 1562 24913 1570
rect 24713 1545 24721 1562
rect 24905 1545 24913 1562
rect 24713 1526 24913 1545
rect 24942 1562 25142 1570
rect 24942 1545 24950 1562
rect 25134 1545 25142 1562
rect 24942 1526 25142 1545
rect 25171 1562 25371 1570
rect 25171 1545 25179 1562
rect 25363 1545 25371 1562
rect 25171 1526 25371 1545
rect 25400 1562 25600 1570
rect 25400 1545 25408 1562
rect 25592 1545 25600 1562
rect 25400 1526 25600 1545
rect 23110 307 23310 326
rect 23110 290 23118 307
rect 23302 290 23310 307
rect 23110 282 23310 290
rect 23339 307 23539 326
rect 23339 290 23347 307
rect 23531 290 23539 307
rect 23339 282 23539 290
rect 23568 307 23768 326
rect 23568 290 23576 307
rect 23760 290 23768 307
rect 23568 282 23768 290
rect 23797 307 23997 326
rect 23797 290 23805 307
rect 23989 290 23997 307
rect 23797 282 23997 290
rect 24026 307 24226 326
rect 24026 290 24034 307
rect 24218 290 24226 307
rect 24026 282 24226 290
rect 24255 307 24455 326
rect 24255 290 24263 307
rect 24447 290 24455 307
rect 24255 282 24455 290
rect 24484 307 24684 326
rect 24484 290 24492 307
rect 24676 290 24684 307
rect 24484 282 24684 290
rect 24713 307 24913 326
rect 24713 290 24721 307
rect 24905 290 24913 307
rect 24713 282 24913 290
rect 24942 307 25142 326
rect 24942 290 24950 307
rect 25134 290 25142 307
rect 24942 282 25142 290
rect 25171 307 25371 326
rect 25171 290 25179 307
rect 25363 290 25371 307
rect 25171 282 25371 290
rect 25400 307 25600 326
rect 25400 290 25408 307
rect 25592 290 25600 307
rect 25400 282 25600 290
rect 28374 1562 28574 1570
rect 28374 1545 28382 1562
rect 28566 1545 28574 1562
rect 28374 1526 28574 1545
rect 28603 1562 28803 1570
rect 28603 1545 28611 1562
rect 28795 1545 28803 1562
rect 28603 1526 28803 1545
rect 28832 1562 29032 1570
rect 28832 1545 28840 1562
rect 29024 1545 29032 1562
rect 28832 1526 29032 1545
rect 29061 1562 29261 1570
rect 29061 1545 29069 1562
rect 29253 1545 29261 1562
rect 29061 1526 29261 1545
rect 29290 1562 29490 1570
rect 29290 1545 29298 1562
rect 29482 1545 29490 1562
rect 29290 1526 29490 1545
rect 29519 1562 29719 1570
rect 29519 1545 29527 1562
rect 29711 1545 29719 1562
rect 29519 1526 29719 1545
rect 29748 1562 29948 1570
rect 29748 1545 29756 1562
rect 29940 1545 29948 1562
rect 29748 1526 29948 1545
rect 29977 1562 30177 1570
rect 29977 1545 29985 1562
rect 30169 1545 30177 1562
rect 29977 1526 30177 1545
rect 30206 1562 30406 1570
rect 30206 1545 30214 1562
rect 30398 1545 30406 1562
rect 30206 1526 30406 1545
rect 30435 1562 30635 1570
rect 30435 1545 30443 1562
rect 30627 1545 30635 1562
rect 30435 1526 30635 1545
rect 30664 1562 30864 1570
rect 30664 1545 30672 1562
rect 30856 1545 30864 1562
rect 30664 1526 30864 1545
rect 28374 307 28574 326
rect 28374 290 28382 307
rect 28566 290 28574 307
rect 28374 282 28574 290
rect 28603 307 28803 326
rect 28603 290 28611 307
rect 28795 290 28803 307
rect 28603 282 28803 290
rect 28832 307 29032 326
rect 28832 290 28840 307
rect 29024 290 29032 307
rect 28832 282 29032 290
rect 29061 307 29261 326
rect 29061 290 29069 307
rect 29253 290 29261 307
rect 29061 282 29261 290
rect 29290 307 29490 326
rect 29290 290 29298 307
rect 29482 290 29490 307
rect 29290 282 29490 290
rect 29519 307 29719 326
rect 29519 290 29527 307
rect 29711 290 29719 307
rect 29519 282 29719 290
rect 29748 307 29948 326
rect 29748 290 29756 307
rect 29940 290 29948 307
rect 29748 282 29948 290
rect 29977 307 30177 326
rect 29977 290 29985 307
rect 30169 290 30177 307
rect 29977 282 30177 290
rect 30206 307 30406 326
rect 30206 290 30214 307
rect 30398 290 30406 307
rect 30206 282 30406 290
rect 30435 307 30635 326
rect 30435 290 30443 307
rect 30627 290 30635 307
rect 30435 282 30635 290
rect 30664 307 30864 326
rect 30664 290 30672 307
rect 30856 290 30864 307
rect 30664 282 30864 290
<< polycont >>
rect 5411 3629 5595 3646
rect 5640 3629 5824 3646
rect 5869 3629 6053 3646
rect 6098 3629 6282 3646
rect 5411 2565 5595 2582
rect 5640 2565 5824 2582
rect 5869 2565 6053 2582
rect 6098 2565 6282 2582
rect 6788 3626 6972 3643
rect 7017 3626 7201 3643
rect 7246 3626 7430 3643
rect 7475 3626 7659 3643
rect 6788 2562 6972 2579
rect 7017 2562 7201 2579
rect 7246 2562 7430 2579
rect 7475 2562 7659 2579
rect 8196 3613 8380 3630
rect 8425 3613 8609 3630
rect 8654 3613 8838 3630
rect 8883 3613 9067 3630
rect 8196 2549 8380 2566
rect 8425 2549 8609 2566
rect 8654 2549 8838 2566
rect 8883 2549 9067 2566
rect 9458 3624 9642 3641
rect 9687 3624 9871 3641
rect 9916 3624 10100 3641
rect 10145 3624 10329 3641
rect 9458 2560 9642 2577
rect 9687 2560 9871 2577
rect 9916 2560 10100 2577
rect 10145 2560 10329 2577
rect 10715 3629 10899 3646
rect 10944 3629 11128 3646
rect 11173 3629 11357 3646
rect 11402 3629 11586 3646
rect 10715 2565 10899 2582
rect 10944 2565 11128 2582
rect 11173 2565 11357 2582
rect 11402 2565 11586 2582
rect 12092 3626 12276 3643
rect 12321 3626 12505 3643
rect 12550 3626 12734 3643
rect 12779 3626 12963 3643
rect 12092 2562 12276 2579
rect 12321 2562 12505 2579
rect 12550 2562 12734 2579
rect 12779 2562 12963 2579
rect 13500 3613 13684 3630
rect 13729 3613 13913 3630
rect 13958 3613 14142 3630
rect 14187 3613 14371 3630
rect 13500 2549 13684 2566
rect 13729 2549 13913 2566
rect 13958 2549 14142 2566
rect 14187 2549 14371 2566
rect 14762 3624 14946 3641
rect 14991 3624 15175 3641
rect 15220 3624 15404 3641
rect 15449 3624 15633 3641
rect 14762 2560 14946 2577
rect 14991 2560 15175 2577
rect 15220 2560 15404 2577
rect 15449 2560 15633 2577
rect 15979 3629 16163 3646
rect 16208 3629 16392 3646
rect 16437 3629 16621 3646
rect 16666 3629 16850 3646
rect 15979 2565 16163 2582
rect 16208 2565 16392 2582
rect 16437 2565 16621 2582
rect 16666 2565 16850 2582
rect 17356 3626 17540 3643
rect 17585 3626 17769 3643
rect 17814 3626 17998 3643
rect 18043 3626 18227 3643
rect 17356 2562 17540 2579
rect 17585 2562 17769 2579
rect 17814 2562 17998 2579
rect 18043 2562 18227 2579
rect 18764 3613 18948 3630
rect 18993 3613 19177 3630
rect 19222 3613 19406 3630
rect 19451 3613 19635 3630
rect 18764 2549 18948 2566
rect 18993 2549 19177 2566
rect 19222 2549 19406 2566
rect 19451 2549 19635 2566
rect 20026 3624 20210 3641
rect 20255 3624 20439 3641
rect 20484 3624 20668 3641
rect 20713 3624 20897 3641
rect 20026 2560 20210 2577
rect 20255 2560 20439 2577
rect 20484 2560 20668 2577
rect 20713 2560 20897 2577
rect 21284 3629 21468 3646
rect 21513 3629 21697 3646
rect 21742 3629 21926 3646
rect 21971 3629 22155 3646
rect 21284 2565 21468 2582
rect 21513 2565 21697 2582
rect 21742 2565 21926 2582
rect 21971 2565 22155 2582
rect 22661 3626 22845 3643
rect 22890 3626 23074 3643
rect 23119 3626 23303 3643
rect 23348 3626 23532 3643
rect 22661 2562 22845 2579
rect 22890 2562 23074 2579
rect 23119 2562 23303 2579
rect 23348 2562 23532 2579
rect 24069 3613 24253 3630
rect 24298 3613 24482 3630
rect 24527 3613 24711 3630
rect 24756 3613 24940 3630
rect 24069 2549 24253 2566
rect 24298 2549 24482 2566
rect 24527 2549 24711 2566
rect 24756 2549 24940 2566
rect 25331 3624 25515 3641
rect 25560 3624 25744 3641
rect 25789 3624 25973 3641
rect 26018 3624 26202 3641
rect 25331 2560 25515 2577
rect 25560 2560 25744 2577
rect 25789 2560 25973 2577
rect 26018 2560 26202 2577
rect 26548 3629 26732 3646
rect 26777 3629 26961 3646
rect 27006 3629 27190 3646
rect 27235 3629 27419 3646
rect 26548 2565 26732 2582
rect 26777 2565 26961 2582
rect 27006 2565 27190 2582
rect 27235 2565 27419 2582
rect 27925 3626 28109 3643
rect 28154 3626 28338 3643
rect 28383 3626 28567 3643
rect 28612 3626 28796 3643
rect 27925 2562 28109 2579
rect 28154 2562 28338 2579
rect 28383 2562 28567 2579
rect 28612 2562 28796 2579
rect 29333 3613 29517 3630
rect 29562 3613 29746 3630
rect 29791 3613 29975 3630
rect 30020 3613 30204 3630
rect 29333 2549 29517 2566
rect 29562 2549 29746 2566
rect 29791 2549 29975 2566
rect 30020 2549 30204 2566
rect 30595 3624 30779 3641
rect 30824 3624 31008 3641
rect 31053 3624 31237 3641
rect 31282 3624 31466 3641
rect 30595 2560 30779 2577
rect 30824 2560 31008 2577
rect 31053 2560 31237 2577
rect 31282 2560 31466 2577
rect 6004 2022 6021 2039
rect 7059 2022 7076 2039
rect 8729 2027 8746 2044
rect 9784 2027 9801 2044
rect 11308 2022 11325 2039
rect 12363 2022 12380 2039
rect 14033 2027 14050 2044
rect 15088 2027 15105 2044
rect 16572 2022 16589 2039
rect 17627 2022 17644 2039
rect 19297 2027 19314 2044
rect 20352 2027 20369 2044
rect 21877 2022 21894 2039
rect 22932 2022 22949 2039
rect 24602 2027 24619 2044
rect 25657 2027 25674 2044
rect 27141 2022 27158 2039
rect 28196 2022 28213 2039
rect 29866 2027 29883 2044
rect 30921 2027 30938 2044
rect 7245 1545 7429 1562
rect 7474 1545 7658 1562
rect 7703 1545 7887 1562
rect 7932 1545 8116 1562
rect 8161 1545 8345 1562
rect 8390 1545 8574 1562
rect 8619 1545 8803 1562
rect 8848 1545 9032 1562
rect 9077 1545 9261 1562
rect 9306 1545 9490 1562
rect 9535 1545 9719 1562
rect 7245 290 7429 307
rect 7474 290 7658 307
rect 7703 290 7887 307
rect 7932 290 8116 307
rect 8161 290 8345 307
rect 8390 290 8574 307
rect 8619 290 8803 307
rect 8848 290 9032 307
rect 9077 290 9261 307
rect 9306 290 9490 307
rect 9535 290 9719 307
rect 12549 1545 12733 1562
rect 12778 1545 12962 1562
rect 13007 1545 13191 1562
rect 13236 1545 13420 1562
rect 13465 1545 13649 1562
rect 13694 1545 13878 1562
rect 13923 1545 14107 1562
rect 14152 1545 14336 1562
rect 14381 1545 14565 1562
rect 14610 1545 14794 1562
rect 14839 1545 15023 1562
rect 12549 290 12733 307
rect 12778 290 12962 307
rect 13007 290 13191 307
rect 13236 290 13420 307
rect 13465 290 13649 307
rect 13694 290 13878 307
rect 13923 290 14107 307
rect 14152 290 14336 307
rect 14381 290 14565 307
rect 14610 290 14794 307
rect 14839 290 15023 307
rect 17813 1545 17997 1562
rect 18042 1545 18226 1562
rect 18271 1545 18455 1562
rect 18500 1545 18684 1562
rect 18729 1545 18913 1562
rect 18958 1545 19142 1562
rect 19187 1545 19371 1562
rect 19416 1545 19600 1562
rect 19645 1545 19829 1562
rect 19874 1545 20058 1562
rect 20103 1545 20287 1562
rect 17813 290 17997 307
rect 18042 290 18226 307
rect 18271 290 18455 307
rect 18500 290 18684 307
rect 18729 290 18913 307
rect 18958 290 19142 307
rect 19187 290 19371 307
rect 19416 290 19600 307
rect 19645 290 19829 307
rect 19874 290 20058 307
rect 20103 290 20287 307
rect 23118 1545 23302 1562
rect 23347 1545 23531 1562
rect 23576 1545 23760 1562
rect 23805 1545 23989 1562
rect 24034 1545 24218 1562
rect 24263 1545 24447 1562
rect 24492 1545 24676 1562
rect 24721 1545 24905 1562
rect 24950 1545 25134 1562
rect 25179 1545 25363 1562
rect 25408 1545 25592 1562
rect 23118 290 23302 307
rect 23347 290 23531 307
rect 23576 290 23760 307
rect 23805 290 23989 307
rect 24034 290 24218 307
rect 24263 290 24447 307
rect 24492 290 24676 307
rect 24721 290 24905 307
rect 24950 290 25134 307
rect 25179 290 25363 307
rect 25408 290 25592 307
rect 28382 1545 28566 1562
rect 28611 1545 28795 1562
rect 28840 1545 29024 1562
rect 29069 1545 29253 1562
rect 29298 1545 29482 1562
rect 29527 1545 29711 1562
rect 29756 1545 29940 1562
rect 29985 1545 30169 1562
rect 30214 1545 30398 1562
rect 30443 1545 30627 1562
rect 30672 1545 30856 1562
rect 28382 290 28566 307
rect 28611 290 28795 307
rect 28840 290 29024 307
rect 29069 290 29253 307
rect 29298 290 29482 307
rect 29527 290 29711 307
rect 29756 290 29940 307
rect 29985 290 30169 307
rect 30214 290 30398 307
rect 30443 290 30627 307
rect 30672 290 30856 307
<< locali >>
rect 9658 3852 10435 3854
rect 14962 3852 15739 3854
rect 20226 3852 21003 3854
rect 25531 3852 26308 3854
rect 30795 3852 31572 3854
rect 7691 3848 9870 3852
rect 7691 3844 8354 3848
rect 6337 3843 8354 3844
rect 6337 3842 8157 3843
rect 5331 3840 8157 3842
rect 5331 3839 7194 3840
rect 5331 3835 6958 3839
rect 5331 3834 6748 3835
rect 5331 3829 6037 3834
rect 5331 3823 5570 3829
rect 5331 3787 5399 3823
rect 5449 3787 5570 3823
rect 5331 3782 5570 3787
rect 5638 3827 6037 3829
rect 5638 3791 5817 3827
rect 5867 3791 6037 3827
rect 5638 3787 6037 3791
rect 6105 3833 6748 3834
rect 6105 3797 6272 3833
rect 6322 3797 6748 3833
rect 6105 3790 6748 3797
rect 6804 3794 6958 3835
rect 7014 3795 7194 3839
rect 7250 3835 8157 3840
rect 7250 3795 7417 3835
rect 7014 3794 7417 3795
rect 6804 3790 7417 3794
rect 7473 3834 8157 3835
rect 7473 3790 7639 3834
rect 6105 3789 7639 3790
rect 7695 3792 8157 3834
rect 8210 3797 8354 3843
rect 8407 3845 9414 3848
rect 8407 3838 8835 3845
rect 8407 3797 8584 3838
rect 8210 3792 8584 3797
rect 7695 3789 8584 3792
rect 6105 3788 8584 3789
rect 6105 3787 7706 3788
rect 8637 3794 8835 3838
rect 8888 3838 9414 3845
rect 8888 3794 9064 3838
rect 8637 3788 9064 3794
rect 9117 3790 9414 3838
rect 9462 3841 9870 3848
rect 9462 3795 9624 3841
rect 9669 3795 9870 3841
rect 9462 3794 9870 3795
rect 9918 3851 10435 3852
rect 9918 3842 10334 3851
rect 9918 3796 10097 3842
rect 10142 3796 10334 3842
rect 9918 3794 10334 3796
rect 9462 3793 10334 3794
rect 10382 3793 10435 3851
rect 12995 3848 15174 3852
rect 12995 3844 13658 3848
rect 11641 3843 13658 3844
rect 11641 3842 13461 3843
rect 9462 3791 10435 3793
rect 10635 3840 13461 3842
rect 10635 3839 12498 3840
rect 10635 3835 12262 3839
rect 10635 3834 12052 3835
rect 10635 3829 11341 3834
rect 10635 3823 10874 3829
rect 9462 3790 9726 3791
rect 9117 3788 9726 3790
rect 10635 3787 10703 3823
rect 10753 3787 10874 3823
rect 5638 3785 7706 3787
rect 5638 3782 6386 3785
rect 10635 3782 10874 3787
rect 10942 3827 11341 3829
rect 10942 3791 11121 3827
rect 11171 3791 11341 3827
rect 10942 3787 11341 3791
rect 11409 3833 12052 3834
rect 11409 3797 11576 3833
rect 11626 3797 12052 3833
rect 11409 3790 12052 3797
rect 12108 3794 12262 3835
rect 12318 3795 12498 3839
rect 12554 3835 13461 3840
rect 12554 3795 12721 3835
rect 12318 3794 12721 3795
rect 12108 3790 12721 3794
rect 12777 3834 13461 3835
rect 12777 3790 12943 3834
rect 11409 3789 12943 3790
rect 12999 3792 13461 3834
rect 13514 3797 13658 3843
rect 13711 3845 14718 3848
rect 13711 3838 14139 3845
rect 13711 3797 13888 3838
rect 13514 3792 13888 3797
rect 12999 3789 13888 3792
rect 11409 3788 13888 3789
rect 11409 3787 13010 3788
rect 13941 3794 14139 3838
rect 14192 3838 14718 3845
rect 14192 3794 14368 3838
rect 13941 3788 14368 3794
rect 14421 3790 14718 3838
rect 14766 3841 15174 3848
rect 14766 3795 14928 3841
rect 14973 3795 15174 3841
rect 14766 3794 15174 3795
rect 15222 3851 15739 3852
rect 15222 3842 15638 3851
rect 15222 3796 15401 3842
rect 15446 3796 15638 3842
rect 15222 3794 15638 3796
rect 14766 3793 15638 3794
rect 15686 3793 15739 3851
rect 18259 3848 20438 3852
rect 18259 3844 18922 3848
rect 16905 3843 18922 3844
rect 16905 3842 18725 3843
rect 14766 3791 15739 3793
rect 15899 3840 18725 3842
rect 15899 3839 17762 3840
rect 15899 3835 17526 3839
rect 15899 3834 17316 3835
rect 15899 3829 16605 3834
rect 15899 3823 16138 3829
rect 14766 3790 15030 3791
rect 14421 3788 15030 3790
rect 15899 3787 15967 3823
rect 16017 3787 16138 3823
rect 10942 3785 13010 3787
rect 10942 3782 11690 3785
rect 15899 3782 16138 3787
rect 16206 3827 16605 3829
rect 16206 3791 16385 3827
rect 16435 3791 16605 3827
rect 16206 3787 16605 3791
rect 16673 3833 17316 3834
rect 16673 3797 16840 3833
rect 16890 3797 17316 3833
rect 16673 3790 17316 3797
rect 17372 3794 17526 3835
rect 17582 3795 17762 3839
rect 17818 3835 18725 3840
rect 17818 3795 17985 3835
rect 17582 3794 17985 3795
rect 17372 3790 17985 3794
rect 18041 3834 18725 3835
rect 18041 3790 18207 3834
rect 16673 3789 18207 3790
rect 18263 3792 18725 3834
rect 18778 3797 18922 3843
rect 18975 3845 19982 3848
rect 18975 3838 19403 3845
rect 18975 3797 19152 3838
rect 18778 3792 19152 3797
rect 18263 3789 19152 3792
rect 16673 3788 19152 3789
rect 16673 3787 18274 3788
rect 19205 3794 19403 3838
rect 19456 3838 19982 3845
rect 19456 3794 19632 3838
rect 19205 3788 19632 3794
rect 19685 3790 19982 3838
rect 20030 3841 20438 3848
rect 20030 3795 20192 3841
rect 20237 3795 20438 3841
rect 20030 3794 20438 3795
rect 20486 3851 21003 3852
rect 20486 3842 20902 3851
rect 20486 3796 20665 3842
rect 20710 3796 20902 3842
rect 20486 3794 20902 3796
rect 20030 3793 20902 3794
rect 20950 3793 21003 3851
rect 23564 3848 25743 3852
rect 23564 3844 24227 3848
rect 22210 3843 24227 3844
rect 22210 3842 24030 3843
rect 20030 3791 21003 3793
rect 21204 3840 24030 3842
rect 21204 3839 23067 3840
rect 21204 3835 22831 3839
rect 21204 3834 22621 3835
rect 21204 3829 21910 3834
rect 21204 3823 21443 3829
rect 20030 3790 20294 3791
rect 19685 3788 20294 3790
rect 21204 3787 21272 3823
rect 21322 3787 21443 3823
rect 16206 3785 18274 3787
rect 16206 3782 16954 3785
rect 21204 3782 21443 3787
rect 21511 3827 21910 3829
rect 21511 3791 21690 3827
rect 21740 3791 21910 3827
rect 21511 3787 21910 3791
rect 21978 3833 22621 3834
rect 21978 3797 22145 3833
rect 22195 3797 22621 3833
rect 21978 3790 22621 3797
rect 22677 3794 22831 3835
rect 22887 3795 23067 3839
rect 23123 3835 24030 3840
rect 23123 3795 23290 3835
rect 22887 3794 23290 3795
rect 22677 3790 23290 3794
rect 23346 3834 24030 3835
rect 23346 3790 23512 3834
rect 21978 3789 23512 3790
rect 23568 3792 24030 3834
rect 24083 3797 24227 3843
rect 24280 3845 25287 3848
rect 24280 3838 24708 3845
rect 24280 3797 24457 3838
rect 24083 3792 24457 3797
rect 23568 3789 24457 3792
rect 21978 3788 24457 3789
rect 21978 3787 23579 3788
rect 24510 3794 24708 3838
rect 24761 3838 25287 3845
rect 24761 3794 24937 3838
rect 24510 3788 24937 3794
rect 24990 3790 25287 3838
rect 25335 3841 25743 3848
rect 25335 3795 25497 3841
rect 25542 3795 25743 3841
rect 25335 3794 25743 3795
rect 25791 3851 26308 3852
rect 25791 3842 26207 3851
rect 25791 3796 25970 3842
rect 26015 3796 26207 3842
rect 25791 3794 26207 3796
rect 25335 3793 26207 3794
rect 26255 3793 26308 3851
rect 28828 3848 31007 3852
rect 28828 3844 29491 3848
rect 27474 3843 29491 3844
rect 27474 3842 29294 3843
rect 25335 3791 26308 3793
rect 26468 3840 29294 3842
rect 26468 3839 28331 3840
rect 26468 3835 28095 3839
rect 26468 3834 27885 3835
rect 26468 3829 27174 3834
rect 26468 3823 26707 3829
rect 25335 3790 25599 3791
rect 24990 3788 25599 3790
rect 26468 3787 26536 3823
rect 26586 3787 26707 3823
rect 21511 3785 23579 3787
rect 21511 3782 22259 3785
rect 26468 3782 26707 3787
rect 26775 3827 27174 3829
rect 26775 3791 26954 3827
rect 27004 3791 27174 3827
rect 26775 3787 27174 3791
rect 27242 3833 27885 3834
rect 27242 3797 27409 3833
rect 27459 3797 27885 3833
rect 27242 3790 27885 3797
rect 27941 3794 28095 3835
rect 28151 3795 28331 3839
rect 28387 3835 29294 3840
rect 28387 3795 28554 3835
rect 28151 3794 28554 3795
rect 27941 3790 28554 3794
rect 28610 3834 29294 3835
rect 28610 3790 28776 3834
rect 27242 3789 28776 3790
rect 28832 3792 29294 3834
rect 29347 3797 29491 3843
rect 29544 3845 30551 3848
rect 29544 3838 29972 3845
rect 29544 3797 29721 3838
rect 29347 3792 29721 3797
rect 28832 3789 29721 3792
rect 27242 3788 29721 3789
rect 27242 3787 28843 3788
rect 29774 3794 29972 3838
rect 30025 3838 30551 3845
rect 30025 3794 30201 3838
rect 29774 3788 30201 3794
rect 30254 3790 30551 3838
rect 30599 3841 31007 3848
rect 30599 3795 30761 3841
rect 30806 3795 31007 3841
rect 30599 3794 31007 3795
rect 31055 3851 31572 3852
rect 31055 3842 31471 3851
rect 31055 3796 31234 3842
rect 31279 3796 31471 3842
rect 31055 3794 31471 3796
rect 30599 3793 31471 3794
rect 31519 3793 31572 3851
rect 30599 3791 31572 3793
rect 30599 3790 30863 3791
rect 30254 3788 30863 3790
rect 26775 3785 28843 3787
rect 26775 3782 27523 3785
rect 5323 3693 5371 3697
rect 5323 3680 5366 3693
rect 6322 3680 6370 3697
rect 5323 3649 5340 3680
rect 6353 3649 6370 3680
rect 5403 3629 5411 3646
rect 5595 3629 5603 3646
rect 5632 3629 5640 3646
rect 5824 3629 5832 3646
rect 5861 3629 5869 3646
rect 6053 3629 6061 3646
rect 6090 3629 6098 3646
rect 6282 3629 6290 3646
rect 5380 3599 5397 3607
rect 5609 3599 5626 3607
rect 5838 3599 5855 3607
rect 5380 2603 5397 2611
rect 5609 2603 5626 2611
rect 6067 3599 6084 3607
rect 6296 3599 6313 3607
rect 5838 2603 5855 2611
rect 6067 2603 6084 2611
rect 6296 2603 6313 2611
rect 5403 2580 5411 2582
rect 5403 2565 5407 2580
rect 5595 2565 5603 2582
rect 5632 2580 5640 2582
rect 5632 2565 5636 2580
rect 5824 2565 5832 2582
rect 5861 2580 5869 2582
rect 5861 2565 5865 2580
rect 6053 2565 6061 2582
rect 6090 2580 6098 2582
rect 6090 2565 6094 2580
rect 6282 2565 6290 2582
rect 5323 2531 5340 2562
rect 6353 2531 6370 2562
rect 5323 2514 5371 2531
rect 6322 2514 6370 2531
rect 6700 3677 6748 3694
rect 7699 3677 7747 3694
rect 10627 3693 10675 3697
rect 6700 3646 6717 3677
rect 7730 3646 7747 3677
rect 6780 3626 6788 3643
rect 6972 3626 6980 3643
rect 7009 3626 7017 3643
rect 7201 3626 7209 3643
rect 7238 3626 7246 3643
rect 7430 3626 7438 3643
rect 7467 3626 7475 3643
rect 7659 3626 7667 3643
rect 6757 3596 6774 3604
rect 6986 3596 7003 3604
rect 7215 3596 7232 3604
rect 6757 2600 6774 2608
rect 6986 2600 7003 2608
rect 7215 2600 7232 2608
rect 7444 3596 7461 3604
rect 7673 3596 7690 3604
rect 7444 2600 7461 2608
rect 7673 2600 7690 2608
rect 6780 2562 6788 2579
rect 6972 2562 6980 2579
rect 7009 2562 7017 2579
rect 7201 2562 7209 2579
rect 7238 2562 7246 2579
rect 7430 2562 7438 2579
rect 7467 2562 7475 2579
rect 7659 2562 7667 2579
rect 6700 2528 6717 2559
rect 7730 2528 7747 2559
rect 6700 2511 6748 2528
rect 7699 2511 7747 2528
rect 8108 3664 8156 3681
rect 9107 3664 9155 3681
rect 8108 3633 8125 3664
rect 9138 3633 9155 3664
rect 8188 3613 8196 3630
rect 8380 3613 8388 3630
rect 8417 3613 8425 3630
rect 8609 3613 8617 3630
rect 8646 3613 8654 3630
rect 8838 3613 8846 3630
rect 8875 3613 8883 3630
rect 9067 3613 9075 3630
rect 8165 3583 8182 3591
rect 8394 3583 8411 3591
rect 8165 2587 8182 2595
rect 8623 3583 8640 3591
rect 8852 3583 8869 3591
rect 8394 2587 8411 2595
rect 8623 2587 8640 2595
rect 9081 3583 9098 3591
rect 8852 2587 8869 2595
rect 9081 2587 9098 2595
rect 8188 2549 8196 2566
rect 8380 2549 8388 2566
rect 8417 2549 8425 2566
rect 8609 2549 8617 2566
rect 8646 2549 8654 2566
rect 8838 2549 8846 2566
rect 8875 2549 8883 2566
rect 9067 2549 9075 2566
rect 8108 2515 8125 2546
rect 9138 2515 9155 2546
rect 8108 2498 8156 2515
rect 9107 2498 9155 2515
rect 9370 3675 9418 3692
rect 10369 3675 10417 3692
rect 9370 3644 9387 3675
rect 10400 3644 10417 3675
rect 9450 3624 9458 3641
rect 9642 3624 9650 3641
rect 9679 3624 9687 3641
rect 9871 3624 9879 3641
rect 9908 3624 9916 3641
rect 10100 3624 10108 3641
rect 10137 3624 10145 3641
rect 10329 3624 10337 3641
rect 9427 3594 9444 3602
rect 9656 3594 9673 3602
rect 9885 3594 9902 3602
rect 10114 3594 10131 3602
rect 9427 2598 9444 2606
rect 9656 2598 9673 2606
rect 10343 3594 10360 3602
rect 9885 2598 9902 2606
rect 10114 2598 10131 2606
rect 10343 2598 10360 2606
rect 9450 2560 9458 2577
rect 9642 2560 9650 2577
rect 9679 2560 9687 2577
rect 9871 2560 9879 2577
rect 9908 2560 9916 2577
rect 10100 2560 10108 2577
rect 10137 2560 10145 2577
rect 10329 2560 10337 2577
rect 9370 2526 9387 2557
rect 10400 2526 10417 2557
rect 9370 2509 9418 2526
rect 10369 2509 10417 2526
rect 10627 3680 10670 3693
rect 11626 3680 11674 3697
rect 10627 3649 10644 3680
rect 11657 3649 11674 3680
rect 10707 3629 10715 3646
rect 10899 3629 10907 3646
rect 10936 3629 10944 3646
rect 11128 3629 11136 3646
rect 11165 3629 11173 3646
rect 11357 3629 11365 3646
rect 11394 3629 11402 3646
rect 11586 3629 11594 3646
rect 10684 3599 10701 3607
rect 10913 3599 10930 3607
rect 11142 3599 11159 3607
rect 10684 2603 10701 2611
rect 10913 2603 10930 2611
rect 11371 3599 11388 3607
rect 11600 3599 11617 3607
rect 11142 2603 11159 2611
rect 11371 2603 11388 2611
rect 11600 2603 11617 2611
rect 10707 2580 10715 2582
rect 10707 2565 10711 2580
rect 10899 2565 10907 2582
rect 10936 2580 10944 2582
rect 10936 2565 10940 2580
rect 11128 2565 11136 2582
rect 11165 2580 11173 2582
rect 11165 2565 11169 2580
rect 11357 2565 11365 2582
rect 11394 2580 11402 2582
rect 11394 2565 11398 2580
rect 11586 2565 11594 2582
rect 10627 2531 10644 2562
rect 11657 2531 11674 2562
rect 10627 2514 10675 2531
rect 11626 2514 11674 2531
rect 12004 3677 12052 3694
rect 13003 3677 13051 3694
rect 15891 3693 15939 3697
rect 12004 3646 12021 3677
rect 13034 3646 13051 3677
rect 12084 3626 12092 3643
rect 12276 3626 12284 3643
rect 12313 3626 12321 3643
rect 12505 3626 12513 3643
rect 12542 3626 12550 3643
rect 12734 3626 12742 3643
rect 12771 3626 12779 3643
rect 12963 3626 12971 3643
rect 12061 3596 12078 3604
rect 12290 3596 12307 3604
rect 12519 3596 12536 3604
rect 12061 2600 12078 2608
rect 12290 2600 12307 2608
rect 12519 2600 12536 2608
rect 12748 3596 12765 3604
rect 12977 3596 12994 3604
rect 12748 2600 12765 2608
rect 12977 2600 12994 2608
rect 12084 2562 12092 2579
rect 12276 2562 12284 2579
rect 12313 2562 12321 2579
rect 12505 2562 12513 2579
rect 12542 2562 12550 2579
rect 12734 2562 12742 2579
rect 12771 2562 12779 2579
rect 12963 2562 12971 2579
rect 12004 2528 12021 2559
rect 13034 2528 13051 2559
rect 12004 2511 12052 2528
rect 13003 2511 13051 2528
rect 13412 3664 13460 3681
rect 14411 3664 14459 3681
rect 13412 3633 13429 3664
rect 14442 3633 14459 3664
rect 13492 3613 13500 3630
rect 13684 3613 13692 3630
rect 13721 3613 13729 3630
rect 13913 3613 13921 3630
rect 13950 3613 13958 3630
rect 14142 3613 14150 3630
rect 14179 3613 14187 3630
rect 14371 3613 14379 3630
rect 13469 3583 13486 3591
rect 13698 3583 13715 3591
rect 13469 2587 13486 2595
rect 13927 3583 13944 3591
rect 14156 3583 14173 3591
rect 13698 2587 13715 2595
rect 13927 2587 13944 2595
rect 14385 3583 14402 3591
rect 14156 2587 14173 2595
rect 14385 2587 14402 2595
rect 13492 2549 13500 2566
rect 13684 2549 13692 2566
rect 13721 2549 13729 2566
rect 13913 2549 13921 2566
rect 13950 2549 13958 2566
rect 14142 2549 14150 2566
rect 14179 2549 14187 2566
rect 14371 2549 14379 2566
rect 13412 2515 13429 2546
rect 14442 2515 14459 2546
rect 13412 2498 13460 2515
rect 14411 2498 14459 2515
rect 14674 3675 14722 3692
rect 15673 3675 15721 3692
rect 14674 3644 14691 3675
rect 15704 3644 15721 3675
rect 14754 3624 14762 3641
rect 14946 3624 14954 3641
rect 14983 3624 14991 3641
rect 15175 3624 15183 3641
rect 15212 3624 15220 3641
rect 15404 3624 15412 3641
rect 15441 3624 15449 3641
rect 15633 3624 15641 3641
rect 14731 3594 14748 3602
rect 14960 3594 14977 3602
rect 15189 3594 15206 3602
rect 15418 3594 15435 3602
rect 14731 2598 14748 2606
rect 14960 2598 14977 2606
rect 15647 3594 15664 3602
rect 15189 2598 15206 2606
rect 15418 2598 15435 2606
rect 15647 2598 15664 2606
rect 14754 2560 14762 2577
rect 14946 2560 14954 2577
rect 14983 2560 14991 2577
rect 15175 2560 15183 2577
rect 15212 2560 15220 2577
rect 15404 2560 15412 2577
rect 15441 2560 15449 2577
rect 15633 2560 15641 2577
rect 14674 2526 14691 2557
rect 15704 2526 15721 2557
rect 14674 2509 14722 2526
rect 15673 2509 15721 2526
rect 15891 3680 15934 3693
rect 16890 3680 16938 3697
rect 15891 3649 15908 3680
rect 16921 3649 16938 3680
rect 15971 3629 15979 3646
rect 16163 3629 16171 3646
rect 16200 3629 16208 3646
rect 16392 3629 16400 3646
rect 16429 3629 16437 3646
rect 16621 3629 16629 3646
rect 16658 3629 16666 3646
rect 16850 3629 16858 3646
rect 15948 3599 15965 3607
rect 16177 3599 16194 3607
rect 16406 3599 16423 3607
rect 15948 2603 15965 2611
rect 16177 2603 16194 2611
rect 16635 3599 16652 3607
rect 16864 3599 16881 3607
rect 16406 2603 16423 2611
rect 16635 2603 16652 2611
rect 16864 2603 16881 2611
rect 15971 2580 15979 2582
rect 15971 2565 15975 2580
rect 16163 2565 16171 2582
rect 16200 2580 16208 2582
rect 16200 2565 16204 2580
rect 16392 2565 16400 2582
rect 16429 2580 16437 2582
rect 16429 2565 16433 2580
rect 16621 2565 16629 2582
rect 16658 2580 16666 2582
rect 16658 2565 16662 2580
rect 16850 2565 16858 2582
rect 15891 2531 15908 2562
rect 16921 2531 16938 2562
rect 15891 2514 15939 2531
rect 16890 2514 16938 2531
rect 17268 3677 17316 3694
rect 18267 3677 18315 3694
rect 21196 3693 21244 3697
rect 17268 3646 17285 3677
rect 18298 3646 18315 3677
rect 17348 3626 17356 3643
rect 17540 3626 17548 3643
rect 17577 3626 17585 3643
rect 17769 3626 17777 3643
rect 17806 3626 17814 3643
rect 17998 3626 18006 3643
rect 18035 3626 18043 3643
rect 18227 3626 18235 3643
rect 17325 3596 17342 3604
rect 17554 3596 17571 3604
rect 17783 3596 17800 3604
rect 17325 2600 17342 2608
rect 17554 2600 17571 2608
rect 17783 2600 17800 2608
rect 18012 3596 18029 3604
rect 18241 3596 18258 3604
rect 18012 2600 18029 2608
rect 18241 2600 18258 2608
rect 17348 2562 17356 2579
rect 17540 2562 17548 2579
rect 17577 2562 17585 2579
rect 17769 2562 17777 2579
rect 17806 2562 17814 2579
rect 17998 2562 18006 2579
rect 18035 2562 18043 2579
rect 18227 2562 18235 2579
rect 17268 2528 17285 2559
rect 18298 2528 18315 2559
rect 17268 2511 17316 2528
rect 18267 2511 18315 2528
rect 18676 3664 18724 3681
rect 19675 3664 19723 3681
rect 18676 3633 18693 3664
rect 19706 3633 19723 3664
rect 18756 3613 18764 3630
rect 18948 3613 18956 3630
rect 18985 3613 18993 3630
rect 19177 3613 19185 3630
rect 19214 3613 19222 3630
rect 19406 3613 19414 3630
rect 19443 3613 19451 3630
rect 19635 3613 19643 3630
rect 18733 3583 18750 3591
rect 18962 3583 18979 3591
rect 18733 2587 18750 2595
rect 19191 3583 19208 3591
rect 19420 3583 19437 3591
rect 18962 2587 18979 2595
rect 19191 2587 19208 2595
rect 19649 3583 19666 3591
rect 19420 2587 19437 2595
rect 19649 2587 19666 2595
rect 18756 2549 18764 2566
rect 18948 2549 18956 2566
rect 18985 2549 18993 2566
rect 19177 2549 19185 2566
rect 19214 2549 19222 2566
rect 19406 2549 19414 2566
rect 19443 2549 19451 2566
rect 19635 2549 19643 2566
rect 18676 2515 18693 2546
rect 19706 2515 19723 2546
rect 18676 2498 18724 2515
rect 19675 2498 19723 2515
rect 19938 3675 19986 3692
rect 20937 3675 20985 3692
rect 19938 3644 19955 3675
rect 20968 3644 20985 3675
rect 20018 3624 20026 3641
rect 20210 3624 20218 3641
rect 20247 3624 20255 3641
rect 20439 3624 20447 3641
rect 20476 3624 20484 3641
rect 20668 3624 20676 3641
rect 20705 3624 20713 3641
rect 20897 3624 20905 3641
rect 19995 3594 20012 3602
rect 20224 3594 20241 3602
rect 20453 3594 20470 3602
rect 20682 3594 20699 3602
rect 19995 2598 20012 2606
rect 20224 2598 20241 2606
rect 20911 3594 20928 3602
rect 20453 2598 20470 2606
rect 20682 2598 20699 2606
rect 20911 2598 20928 2606
rect 20018 2560 20026 2577
rect 20210 2560 20218 2577
rect 20247 2560 20255 2577
rect 20439 2560 20447 2577
rect 20476 2560 20484 2577
rect 20668 2560 20676 2577
rect 20705 2560 20713 2577
rect 20897 2560 20905 2577
rect 19938 2526 19955 2557
rect 20968 2526 20985 2557
rect 19938 2509 19986 2526
rect 20937 2509 20985 2526
rect 21196 3680 21239 3693
rect 22195 3680 22243 3697
rect 21196 3649 21213 3680
rect 22226 3649 22243 3680
rect 21276 3629 21284 3646
rect 21468 3629 21476 3646
rect 21505 3629 21513 3646
rect 21697 3629 21705 3646
rect 21734 3629 21742 3646
rect 21926 3629 21934 3646
rect 21963 3629 21971 3646
rect 22155 3629 22163 3646
rect 21253 3599 21270 3607
rect 21482 3599 21499 3607
rect 21711 3599 21728 3607
rect 21253 2603 21270 2611
rect 21482 2603 21499 2611
rect 21940 3599 21957 3607
rect 22169 3599 22186 3607
rect 21711 2603 21728 2611
rect 21940 2603 21957 2611
rect 22169 2603 22186 2611
rect 21276 2580 21284 2582
rect 21276 2565 21280 2580
rect 21468 2565 21476 2582
rect 21505 2580 21513 2582
rect 21505 2565 21509 2580
rect 21697 2565 21705 2582
rect 21734 2580 21742 2582
rect 21734 2565 21738 2580
rect 21926 2565 21934 2582
rect 21963 2580 21971 2582
rect 21963 2565 21967 2580
rect 22155 2565 22163 2582
rect 21196 2531 21213 2562
rect 22226 2531 22243 2562
rect 21196 2514 21244 2531
rect 22195 2514 22243 2531
rect 22573 3677 22621 3694
rect 23572 3677 23620 3694
rect 26460 3693 26508 3697
rect 22573 3646 22590 3677
rect 23603 3646 23620 3677
rect 22653 3626 22661 3643
rect 22845 3626 22853 3643
rect 22882 3626 22890 3643
rect 23074 3626 23082 3643
rect 23111 3626 23119 3643
rect 23303 3626 23311 3643
rect 23340 3626 23348 3643
rect 23532 3626 23540 3643
rect 22630 3596 22647 3604
rect 22859 3596 22876 3604
rect 23088 3596 23105 3604
rect 22630 2600 22647 2608
rect 22859 2600 22876 2608
rect 23088 2600 23105 2608
rect 23317 3596 23334 3604
rect 23546 3596 23563 3604
rect 23317 2600 23334 2608
rect 23546 2600 23563 2608
rect 22653 2562 22661 2579
rect 22845 2562 22853 2579
rect 22882 2562 22890 2579
rect 23074 2562 23082 2579
rect 23111 2562 23119 2579
rect 23303 2562 23311 2579
rect 23340 2562 23348 2579
rect 23532 2562 23540 2579
rect 22573 2528 22590 2559
rect 23603 2528 23620 2559
rect 22573 2511 22621 2528
rect 23572 2511 23620 2528
rect 23981 3664 24029 3681
rect 24980 3664 25028 3681
rect 23981 3633 23998 3664
rect 25011 3633 25028 3664
rect 24061 3613 24069 3630
rect 24253 3613 24261 3630
rect 24290 3613 24298 3630
rect 24482 3613 24490 3630
rect 24519 3613 24527 3630
rect 24711 3613 24719 3630
rect 24748 3613 24756 3630
rect 24940 3613 24948 3630
rect 24038 3583 24055 3591
rect 24267 3583 24284 3591
rect 24038 2587 24055 2595
rect 24496 3583 24513 3591
rect 24725 3583 24742 3591
rect 24267 2587 24284 2595
rect 24496 2587 24513 2595
rect 24954 3583 24971 3591
rect 24725 2587 24742 2595
rect 24954 2587 24971 2595
rect 24061 2549 24069 2566
rect 24253 2549 24261 2566
rect 24290 2549 24298 2566
rect 24482 2549 24490 2566
rect 24519 2549 24527 2566
rect 24711 2549 24719 2566
rect 24748 2549 24756 2566
rect 24940 2549 24948 2566
rect 23981 2515 23998 2546
rect 25011 2515 25028 2546
rect 23981 2498 24029 2515
rect 24980 2498 25028 2515
rect 25243 3675 25291 3692
rect 26242 3675 26290 3692
rect 25243 3644 25260 3675
rect 26273 3644 26290 3675
rect 25323 3624 25331 3641
rect 25515 3624 25523 3641
rect 25552 3624 25560 3641
rect 25744 3624 25752 3641
rect 25781 3624 25789 3641
rect 25973 3624 25981 3641
rect 26010 3624 26018 3641
rect 26202 3624 26210 3641
rect 25300 3594 25317 3602
rect 25529 3594 25546 3602
rect 25758 3594 25775 3602
rect 25987 3594 26004 3602
rect 25300 2598 25317 2606
rect 25529 2598 25546 2606
rect 26216 3594 26233 3602
rect 25758 2598 25775 2606
rect 25987 2598 26004 2606
rect 26216 2598 26233 2606
rect 25323 2560 25331 2577
rect 25515 2560 25523 2577
rect 25552 2560 25560 2577
rect 25744 2560 25752 2577
rect 25781 2560 25789 2577
rect 25973 2560 25981 2577
rect 26010 2560 26018 2577
rect 26202 2560 26210 2577
rect 25243 2526 25260 2557
rect 26273 2526 26290 2557
rect 25243 2509 25291 2526
rect 26242 2509 26290 2526
rect 26460 3680 26503 3693
rect 27459 3680 27507 3697
rect 26460 3649 26477 3680
rect 27490 3649 27507 3680
rect 26540 3629 26548 3646
rect 26732 3629 26740 3646
rect 26769 3629 26777 3646
rect 26961 3629 26969 3646
rect 26998 3629 27006 3646
rect 27190 3629 27198 3646
rect 27227 3629 27235 3646
rect 27419 3629 27427 3646
rect 26517 3599 26534 3607
rect 26746 3599 26763 3607
rect 26975 3599 26992 3607
rect 26517 2603 26534 2611
rect 26746 2603 26763 2611
rect 27204 3599 27221 3607
rect 27433 3599 27450 3607
rect 26975 2603 26992 2611
rect 27204 2603 27221 2611
rect 27433 2603 27450 2611
rect 26540 2580 26548 2582
rect 26540 2565 26544 2580
rect 26732 2565 26740 2582
rect 26769 2580 26777 2582
rect 26769 2565 26773 2580
rect 26961 2565 26969 2582
rect 26998 2580 27006 2582
rect 26998 2565 27002 2580
rect 27190 2565 27198 2582
rect 27227 2580 27235 2582
rect 27227 2565 27231 2580
rect 27419 2565 27427 2582
rect 26460 2531 26477 2562
rect 27490 2531 27507 2562
rect 26460 2514 26508 2531
rect 27459 2514 27507 2531
rect 27837 3677 27885 3694
rect 28836 3677 28884 3694
rect 27837 3646 27854 3677
rect 28867 3646 28884 3677
rect 27917 3626 27925 3643
rect 28109 3626 28117 3643
rect 28146 3626 28154 3643
rect 28338 3626 28346 3643
rect 28375 3626 28383 3643
rect 28567 3626 28575 3643
rect 28604 3626 28612 3643
rect 28796 3626 28804 3643
rect 27894 3596 27911 3604
rect 28123 3596 28140 3604
rect 28352 3596 28369 3604
rect 27894 2600 27911 2608
rect 28123 2600 28140 2608
rect 28352 2600 28369 2608
rect 28581 3596 28598 3604
rect 28810 3596 28827 3604
rect 28581 2600 28598 2608
rect 28810 2600 28827 2608
rect 27917 2562 27925 2579
rect 28109 2562 28117 2579
rect 28146 2562 28154 2579
rect 28338 2562 28346 2579
rect 28375 2562 28383 2579
rect 28567 2562 28575 2579
rect 28604 2562 28612 2579
rect 28796 2562 28804 2579
rect 27837 2528 27854 2559
rect 28867 2528 28884 2559
rect 27837 2511 27885 2528
rect 28836 2511 28884 2528
rect 29245 3664 29293 3681
rect 30244 3664 30292 3681
rect 29245 3633 29262 3664
rect 30275 3633 30292 3664
rect 29325 3613 29333 3630
rect 29517 3613 29525 3630
rect 29554 3613 29562 3630
rect 29746 3613 29754 3630
rect 29783 3613 29791 3630
rect 29975 3613 29983 3630
rect 30012 3613 30020 3630
rect 30204 3613 30212 3630
rect 29302 3583 29319 3591
rect 29531 3583 29548 3591
rect 29302 2587 29319 2595
rect 29760 3583 29777 3591
rect 29989 3583 30006 3591
rect 29531 2587 29548 2595
rect 29760 2587 29777 2595
rect 30218 3583 30235 3591
rect 29989 2587 30006 2595
rect 30218 2587 30235 2595
rect 29325 2549 29333 2566
rect 29517 2549 29525 2566
rect 29554 2549 29562 2566
rect 29746 2549 29754 2566
rect 29783 2549 29791 2566
rect 29975 2549 29983 2566
rect 30012 2549 30020 2566
rect 30204 2549 30212 2566
rect 29245 2515 29262 2546
rect 30275 2515 30292 2546
rect 29245 2498 29293 2515
rect 30244 2498 30292 2515
rect 30507 3675 30555 3692
rect 31506 3675 31554 3692
rect 30507 3644 30524 3675
rect 31537 3644 31554 3675
rect 30587 3624 30595 3641
rect 30779 3624 30787 3641
rect 30816 3624 30824 3641
rect 31008 3624 31016 3641
rect 31045 3624 31053 3641
rect 31237 3624 31245 3641
rect 31274 3624 31282 3641
rect 31466 3624 31474 3641
rect 30564 3594 30581 3602
rect 30793 3594 30810 3602
rect 31022 3594 31039 3602
rect 31251 3594 31268 3602
rect 30564 2598 30581 2606
rect 30793 2598 30810 2606
rect 31480 3594 31497 3602
rect 31022 2598 31039 2606
rect 31251 2598 31268 2606
rect 31480 2598 31497 2606
rect 30587 2560 30595 2577
rect 30779 2560 30787 2577
rect 30816 2560 30824 2577
rect 31008 2560 31016 2577
rect 31045 2560 31053 2577
rect 31237 2560 31245 2577
rect 31274 2560 31282 2577
rect 31466 2560 31474 2577
rect 30507 2526 30524 2557
rect 31537 2526 31554 2557
rect 30507 2509 30555 2526
rect 31506 2509 31554 2526
rect 5953 2101 6001 2118
rect 7079 2101 7127 2118
rect 5953 2070 5970 2101
rect 7110 2070 7127 2101
rect 6004 2039 6021 2047
rect 6038 2044 6046 2061
rect 7034 2044 7042 2061
rect 6004 2014 6021 2022
rect 7059 2039 7076 2047
rect 6038 2000 6046 2017
rect 7034 2000 7042 2017
rect 7059 2014 7076 2022
rect 5953 1960 5970 1991
rect 7110 1960 7127 1991
rect 5953 1943 6001 1960
rect 7079 1943 7127 1960
rect 8678 2106 8726 2123
rect 9804 2106 9852 2123
rect 8678 2075 8695 2106
rect 9835 2075 9852 2106
rect 8729 2044 8746 2052
rect 8763 2049 8771 2066
rect 9759 2049 9767 2066
rect 8729 2019 8746 2027
rect 9784 2044 9801 2052
rect 8763 2005 8771 2022
rect 9759 2005 9767 2022
rect 9784 2019 9801 2027
rect 8678 1965 8695 1996
rect 9835 1965 9852 1996
rect 8678 1948 8726 1965
rect 9804 1948 9852 1965
rect 11257 2101 11305 2118
rect 12383 2101 12431 2118
rect 11257 2070 11274 2101
rect 12414 2070 12431 2101
rect 11308 2039 11325 2047
rect 11342 2044 11350 2061
rect 12338 2044 12346 2061
rect 11308 2014 11325 2022
rect 12363 2039 12380 2047
rect 11342 2000 11350 2017
rect 12338 2000 12346 2017
rect 12363 2014 12380 2022
rect 11257 1960 11274 1991
rect 12414 1960 12431 1991
rect 11257 1943 11305 1960
rect 12383 1943 12431 1960
rect 13982 2106 14030 2123
rect 15108 2106 15156 2123
rect 13982 2075 13999 2106
rect 15139 2075 15156 2106
rect 14033 2044 14050 2052
rect 14067 2049 14075 2066
rect 15063 2049 15071 2066
rect 14033 2019 14050 2027
rect 15088 2044 15105 2052
rect 14067 2005 14075 2022
rect 15063 2005 15071 2022
rect 15088 2019 15105 2027
rect 13982 1965 13999 1996
rect 15139 1965 15156 1996
rect 13982 1948 14030 1965
rect 15108 1948 15156 1965
rect 16521 2101 16569 2118
rect 17647 2101 17695 2118
rect 16521 2070 16538 2101
rect 17678 2070 17695 2101
rect 16572 2039 16589 2047
rect 16606 2044 16614 2061
rect 17602 2044 17610 2061
rect 16572 2014 16589 2022
rect 17627 2039 17644 2047
rect 16606 2000 16614 2017
rect 17602 2000 17610 2017
rect 17627 2014 17644 2022
rect 16521 1960 16538 1991
rect 17678 1960 17695 1991
rect 16521 1943 16569 1960
rect 17647 1943 17695 1960
rect 19246 2106 19294 2123
rect 20372 2106 20420 2123
rect 19246 2075 19263 2106
rect 20403 2075 20420 2106
rect 19297 2044 19314 2052
rect 19331 2049 19339 2066
rect 20327 2049 20335 2066
rect 19297 2019 19314 2027
rect 20352 2044 20369 2052
rect 19331 2005 19339 2022
rect 20327 2005 20335 2022
rect 20352 2019 20369 2027
rect 19246 1965 19263 1996
rect 20403 1965 20420 1996
rect 19246 1948 19294 1965
rect 20372 1948 20420 1965
rect 21826 2101 21874 2118
rect 22952 2101 23000 2118
rect 21826 2070 21843 2101
rect 22983 2070 23000 2101
rect 21877 2039 21894 2047
rect 21911 2044 21919 2061
rect 22907 2044 22915 2061
rect 21877 2014 21894 2022
rect 22932 2039 22949 2047
rect 21911 2000 21919 2017
rect 22907 2000 22915 2017
rect 22932 2014 22949 2022
rect 21826 1960 21843 1991
rect 22983 1960 23000 1991
rect 21826 1943 21874 1960
rect 22952 1943 23000 1960
rect 24551 2106 24599 2123
rect 25677 2106 25725 2123
rect 24551 2075 24568 2106
rect 25708 2075 25725 2106
rect 24602 2044 24619 2052
rect 24636 2049 24644 2066
rect 25632 2049 25640 2066
rect 24602 2019 24619 2027
rect 25657 2044 25674 2052
rect 24636 2005 24644 2022
rect 25632 2005 25640 2022
rect 25657 2019 25674 2027
rect 24551 1965 24568 1996
rect 25708 1965 25725 1996
rect 24551 1948 24599 1965
rect 25677 1948 25725 1965
rect 27090 2101 27138 2118
rect 28216 2101 28264 2118
rect 27090 2070 27107 2101
rect 28247 2070 28264 2101
rect 27141 2039 27158 2047
rect 27175 2044 27183 2061
rect 28171 2044 28179 2061
rect 27141 2014 27158 2022
rect 28196 2039 28213 2047
rect 27175 2000 27183 2017
rect 28171 2000 28179 2017
rect 28196 2014 28213 2022
rect 27090 1960 27107 1991
rect 28247 1960 28264 1991
rect 27090 1943 27138 1960
rect 28216 1943 28264 1960
rect 29815 2106 29863 2123
rect 30941 2106 30989 2123
rect 29815 2075 29832 2106
rect 30972 2075 30989 2106
rect 29866 2044 29883 2052
rect 29900 2049 29908 2066
rect 30896 2049 30904 2066
rect 29866 2019 29883 2027
rect 30921 2044 30938 2052
rect 29900 2005 29908 2022
rect 30896 2005 30904 2022
rect 30921 2019 30938 2027
rect 29815 1965 29832 1996
rect 30972 1965 30989 1996
rect 29815 1948 29863 1965
rect 30941 1948 30989 1965
rect 7157 1596 7205 1613
rect 9759 1596 9807 1613
rect 7157 1565 7174 1596
rect 9790 1565 9807 1596
rect 7237 1545 7245 1562
rect 7429 1545 7437 1562
rect 7466 1545 7474 1562
rect 7658 1545 7666 1562
rect 7695 1545 7703 1562
rect 7887 1545 7895 1562
rect 7924 1545 7932 1562
rect 8116 1545 8124 1562
rect 8153 1545 8161 1562
rect 8345 1545 8353 1562
rect 8382 1545 8390 1562
rect 8574 1545 8582 1562
rect 8611 1545 8619 1562
rect 8803 1545 8811 1562
rect 8840 1545 8848 1562
rect 9032 1545 9040 1562
rect 9069 1545 9077 1562
rect 9261 1545 9269 1562
rect 9298 1545 9306 1562
rect 9490 1545 9498 1562
rect 9527 1545 9535 1562
rect 9719 1545 9727 1562
rect 7214 1520 7231 1528
rect 7443 1520 7460 1528
rect 7672 1520 7689 1528
rect 7901 1520 7918 1528
rect 7214 324 7231 332
rect 7443 324 7460 332
rect 8130 1520 8147 1528
rect 8359 1520 8376 1528
rect 7672 324 7689 332
rect 7901 324 7918 332
rect 8588 1520 8605 1528
rect 8817 1520 8834 1528
rect 8130 324 8147 332
rect 8359 324 8376 332
rect 9046 1520 9063 1528
rect 8588 324 8605 332
rect 8817 324 8834 332
rect 9275 1520 9292 1528
rect 9504 1520 9521 1528
rect 9733 1520 9750 1528
rect 9046 324 9063 332
rect 9275 324 9292 332
rect 9504 324 9521 332
rect 9733 324 9750 332
rect 7237 290 7245 307
rect 7429 290 7437 307
rect 7466 290 7474 307
rect 7658 290 7666 307
rect 7695 290 7703 307
rect 7887 290 7895 307
rect 7924 290 7932 307
rect 8116 290 8124 307
rect 8153 290 8161 307
rect 8345 290 8353 307
rect 8382 290 8390 307
rect 8574 290 8582 307
rect 8611 290 8619 307
rect 8803 290 8811 307
rect 8840 290 8848 307
rect 9032 290 9040 307
rect 9069 290 9077 307
rect 9261 290 9269 307
rect 9298 290 9306 307
rect 9490 290 9498 307
rect 9527 290 9535 307
rect 9719 290 9727 307
rect 7157 256 7174 287
rect 9790 256 9807 287
rect 7157 239 7205 256
rect 9759 239 9807 256
rect 12461 1596 12509 1613
rect 15063 1596 15111 1613
rect 12461 1565 12478 1596
rect 15094 1565 15111 1596
rect 12541 1545 12549 1562
rect 12733 1545 12741 1562
rect 12770 1545 12778 1562
rect 12962 1545 12970 1562
rect 12999 1545 13007 1562
rect 13191 1545 13199 1562
rect 13228 1545 13236 1562
rect 13420 1545 13428 1562
rect 13457 1545 13465 1562
rect 13649 1545 13657 1562
rect 13686 1545 13694 1562
rect 13878 1545 13886 1562
rect 13915 1545 13923 1562
rect 14107 1545 14115 1562
rect 14144 1545 14152 1562
rect 14336 1545 14344 1562
rect 14373 1545 14381 1562
rect 14565 1545 14573 1562
rect 14602 1545 14610 1562
rect 14794 1545 14802 1562
rect 14831 1545 14839 1562
rect 15023 1545 15031 1562
rect 12518 1520 12535 1528
rect 12747 1520 12764 1528
rect 12976 1520 12993 1528
rect 13205 1520 13222 1528
rect 12518 324 12535 332
rect 12747 324 12764 332
rect 13434 1520 13451 1528
rect 13663 1520 13680 1528
rect 12976 324 12993 332
rect 13205 324 13222 332
rect 13892 1520 13909 1528
rect 14121 1520 14138 1528
rect 13434 324 13451 332
rect 13663 324 13680 332
rect 14350 1520 14367 1528
rect 13892 324 13909 332
rect 14121 324 14138 332
rect 14579 1520 14596 1528
rect 14808 1520 14825 1528
rect 15037 1520 15054 1528
rect 14350 324 14367 332
rect 14579 324 14596 332
rect 14808 324 14825 332
rect 15037 324 15054 332
rect 12541 290 12549 307
rect 12733 290 12741 307
rect 12770 290 12778 307
rect 12962 290 12970 307
rect 12999 290 13007 307
rect 13191 290 13199 307
rect 13228 290 13236 307
rect 13420 290 13428 307
rect 13457 290 13465 307
rect 13649 290 13657 307
rect 13686 290 13694 307
rect 13878 290 13886 307
rect 13915 290 13923 307
rect 14107 290 14115 307
rect 14144 290 14152 307
rect 14336 290 14344 307
rect 14373 290 14381 307
rect 14565 290 14573 307
rect 14602 290 14610 307
rect 14794 290 14802 307
rect 14831 290 14839 307
rect 15023 290 15031 307
rect 12461 256 12478 287
rect 15094 256 15111 287
rect 12461 239 12509 256
rect 15063 239 15111 256
rect 17725 1596 17773 1613
rect 20327 1596 20375 1613
rect 17725 1565 17742 1596
rect 20358 1565 20375 1596
rect 17805 1545 17813 1562
rect 17997 1545 18005 1562
rect 18034 1545 18042 1562
rect 18226 1545 18234 1562
rect 18263 1545 18271 1562
rect 18455 1545 18463 1562
rect 18492 1545 18500 1562
rect 18684 1545 18692 1562
rect 18721 1545 18729 1562
rect 18913 1545 18921 1562
rect 18950 1545 18958 1562
rect 19142 1545 19150 1562
rect 19179 1545 19187 1562
rect 19371 1545 19379 1562
rect 19408 1545 19416 1562
rect 19600 1545 19608 1562
rect 19637 1545 19645 1562
rect 19829 1545 19837 1562
rect 19866 1545 19874 1562
rect 20058 1545 20066 1562
rect 20095 1545 20103 1562
rect 20287 1545 20295 1562
rect 17782 1520 17799 1528
rect 18011 1520 18028 1528
rect 18240 1520 18257 1528
rect 18469 1520 18486 1528
rect 17782 324 17799 332
rect 18011 324 18028 332
rect 18698 1520 18715 1528
rect 18927 1520 18944 1528
rect 18240 324 18257 332
rect 18469 324 18486 332
rect 19156 1520 19173 1528
rect 19385 1520 19402 1528
rect 18698 324 18715 332
rect 18927 324 18944 332
rect 19614 1520 19631 1528
rect 19156 324 19173 332
rect 19385 324 19402 332
rect 19843 1520 19860 1528
rect 20072 1520 20089 1528
rect 20301 1520 20318 1528
rect 19614 324 19631 332
rect 19843 324 19860 332
rect 20072 324 20089 332
rect 20301 324 20318 332
rect 17805 290 17813 307
rect 17997 290 18005 307
rect 18034 290 18042 307
rect 18226 290 18234 307
rect 18263 290 18271 307
rect 18455 290 18463 307
rect 18492 290 18500 307
rect 18684 290 18692 307
rect 18721 290 18729 307
rect 18913 290 18921 307
rect 18950 290 18958 307
rect 19142 290 19150 307
rect 19179 290 19187 307
rect 19371 290 19379 307
rect 19408 290 19416 307
rect 19600 290 19608 307
rect 19637 290 19645 307
rect 19829 290 19837 307
rect 19866 290 19874 307
rect 20058 290 20066 307
rect 20095 290 20103 307
rect 20287 290 20295 307
rect 17725 256 17742 287
rect 20358 256 20375 287
rect 17725 239 17773 256
rect 20327 239 20375 256
rect 23030 1596 23078 1613
rect 25632 1596 25680 1613
rect 23030 1565 23047 1596
rect 25663 1565 25680 1596
rect 23110 1545 23118 1562
rect 23302 1545 23310 1562
rect 23339 1545 23347 1562
rect 23531 1545 23539 1562
rect 23568 1545 23576 1562
rect 23760 1545 23768 1562
rect 23797 1545 23805 1562
rect 23989 1545 23997 1562
rect 24026 1545 24034 1562
rect 24218 1545 24226 1562
rect 24255 1545 24263 1562
rect 24447 1545 24455 1562
rect 24484 1545 24492 1562
rect 24676 1545 24684 1562
rect 24713 1545 24721 1562
rect 24905 1545 24913 1562
rect 24942 1545 24950 1562
rect 25134 1545 25142 1562
rect 25171 1545 25179 1562
rect 25363 1545 25371 1562
rect 25400 1545 25408 1562
rect 25592 1545 25600 1562
rect 23087 1520 23104 1528
rect 23316 1520 23333 1528
rect 23545 1520 23562 1528
rect 23774 1520 23791 1528
rect 23087 324 23104 332
rect 23316 324 23333 332
rect 24003 1520 24020 1528
rect 24232 1520 24249 1528
rect 23545 324 23562 332
rect 23774 324 23791 332
rect 24461 1520 24478 1528
rect 24690 1520 24707 1528
rect 24003 324 24020 332
rect 24232 324 24249 332
rect 24919 1520 24936 1528
rect 24461 324 24478 332
rect 24690 324 24707 332
rect 25148 1520 25165 1528
rect 25377 1520 25394 1528
rect 25606 1520 25623 1528
rect 24919 324 24936 332
rect 25148 324 25165 332
rect 25377 324 25394 332
rect 25606 324 25623 332
rect 23110 290 23118 307
rect 23302 290 23310 307
rect 23339 290 23347 307
rect 23531 290 23539 307
rect 23568 290 23576 307
rect 23760 290 23768 307
rect 23797 290 23805 307
rect 23989 290 23997 307
rect 24026 290 24034 307
rect 24218 290 24226 307
rect 24255 290 24263 307
rect 24447 290 24455 307
rect 24484 290 24492 307
rect 24676 290 24684 307
rect 24713 290 24721 307
rect 24905 290 24913 307
rect 24942 290 24950 307
rect 25134 290 25142 307
rect 25171 290 25179 307
rect 25363 290 25371 307
rect 25400 290 25408 307
rect 25592 290 25600 307
rect 23030 256 23047 287
rect 25663 256 25680 287
rect 23030 239 23078 256
rect 25632 239 25680 256
rect 28294 1596 28342 1613
rect 30896 1596 30944 1613
rect 28294 1565 28311 1596
rect 30927 1565 30944 1596
rect 28374 1545 28382 1562
rect 28566 1545 28574 1562
rect 28603 1545 28611 1562
rect 28795 1545 28803 1562
rect 28832 1545 28840 1562
rect 29024 1545 29032 1562
rect 29061 1545 29069 1562
rect 29253 1545 29261 1562
rect 29290 1545 29298 1562
rect 29482 1545 29490 1562
rect 29519 1545 29527 1562
rect 29711 1545 29719 1562
rect 29748 1545 29756 1562
rect 29940 1545 29948 1562
rect 29977 1545 29985 1562
rect 30169 1545 30177 1562
rect 30206 1545 30214 1562
rect 30398 1545 30406 1562
rect 30435 1545 30443 1562
rect 30627 1545 30635 1562
rect 30664 1545 30672 1562
rect 30856 1545 30864 1562
rect 28351 1520 28368 1528
rect 28580 1520 28597 1528
rect 28809 1520 28826 1528
rect 29038 1520 29055 1528
rect 28351 324 28368 332
rect 28580 324 28597 332
rect 29267 1520 29284 1528
rect 29496 1520 29513 1528
rect 28809 324 28826 332
rect 29038 324 29055 332
rect 29725 1520 29742 1528
rect 29954 1520 29971 1528
rect 29267 324 29284 332
rect 29496 324 29513 332
rect 30183 1520 30200 1528
rect 29725 324 29742 332
rect 29954 324 29971 332
rect 30412 1520 30429 1528
rect 30641 1520 30658 1528
rect 30870 1520 30887 1528
rect 30183 324 30200 332
rect 30412 324 30429 332
rect 30641 324 30658 332
rect 30870 324 30887 332
rect 28374 290 28382 307
rect 28566 290 28574 307
rect 28603 290 28611 307
rect 28795 290 28803 307
rect 28832 290 28840 307
rect 29024 290 29032 307
rect 29061 290 29069 307
rect 29253 290 29261 307
rect 29290 290 29298 307
rect 29482 290 29490 307
rect 29519 290 29527 307
rect 29711 290 29719 307
rect 29748 290 29756 307
rect 29940 290 29948 307
rect 29977 290 29985 307
rect 30169 290 30177 307
rect 30206 290 30214 307
rect 30398 290 30406 307
rect 30435 290 30443 307
rect 30627 290 30635 307
rect 30664 290 30672 307
rect 30856 290 30864 307
rect 28294 256 28311 287
rect 30927 256 30944 287
rect 28294 239 28342 256
rect 30896 239 30944 256
rect 7135 139 9874 140
rect 7135 136 8574 139
rect 7135 82 7186 136
rect 7243 132 8104 136
rect 7243 129 7861 132
rect 7243 82 7414 129
rect 7135 71 7414 82
rect 7493 128 7861 129
rect 7493 74 7659 128
rect 7716 74 7861 128
rect 7940 82 8104 132
rect 8161 85 8574 136
rect 8631 136 9485 139
rect 8631 132 9038 136
rect 8631 85 8746 132
rect 8161 82 8746 85
rect 7940 74 8746 82
rect 8825 82 9038 132
rect 9095 134 9485 136
rect 9095 82 9295 134
rect 8825 76 9295 82
rect 9374 85 9485 134
rect 9542 85 9874 139
rect 9374 76 9874 85
rect 8825 74 9874 76
rect 7493 71 9874 74
rect 7135 65 9874 71
rect 12439 139 15178 140
rect 12439 136 13878 139
rect 12439 82 12490 136
rect 12547 132 13408 136
rect 12547 129 13165 132
rect 12547 82 12718 129
rect 12439 71 12718 82
rect 12797 128 13165 129
rect 12797 74 12963 128
rect 13020 74 13165 128
rect 13244 82 13408 132
rect 13465 85 13878 136
rect 13935 136 14789 139
rect 13935 132 14342 136
rect 13935 85 14050 132
rect 13465 82 14050 85
rect 13244 74 14050 82
rect 14129 82 14342 132
rect 14399 134 14789 136
rect 14399 82 14599 134
rect 14129 76 14599 82
rect 14678 85 14789 134
rect 14846 85 15178 139
rect 14678 76 15178 85
rect 14129 74 15178 76
rect 12797 71 15178 74
rect 12439 65 15178 71
rect 17703 139 20442 140
rect 17703 136 19142 139
rect 17703 82 17754 136
rect 17811 132 18672 136
rect 17811 129 18429 132
rect 17811 82 17982 129
rect 17703 71 17982 82
rect 18061 128 18429 129
rect 18061 74 18227 128
rect 18284 74 18429 128
rect 18508 82 18672 132
rect 18729 85 19142 136
rect 19199 136 20053 139
rect 19199 132 19606 136
rect 19199 85 19314 132
rect 18729 82 19314 85
rect 18508 74 19314 82
rect 19393 82 19606 132
rect 19663 134 20053 136
rect 19663 82 19863 134
rect 19393 76 19863 82
rect 19942 85 20053 134
rect 20110 85 20442 139
rect 19942 76 20442 85
rect 19393 74 20442 76
rect 18061 71 20442 74
rect 17703 65 20442 71
rect 23008 139 25747 140
rect 23008 136 24447 139
rect 23008 82 23059 136
rect 23116 132 23977 136
rect 23116 129 23734 132
rect 23116 82 23287 129
rect 23008 71 23287 82
rect 23366 128 23734 129
rect 23366 74 23532 128
rect 23589 74 23734 128
rect 23813 82 23977 132
rect 24034 85 24447 136
rect 24504 136 25358 139
rect 24504 132 24911 136
rect 24504 85 24619 132
rect 24034 82 24619 85
rect 23813 74 24619 82
rect 24698 82 24911 132
rect 24968 134 25358 136
rect 24968 82 25168 134
rect 24698 76 25168 82
rect 25247 85 25358 134
rect 25415 85 25747 139
rect 25247 76 25747 85
rect 24698 74 25747 76
rect 23366 71 25747 74
rect 23008 65 25747 71
rect 28272 139 31011 140
rect 28272 136 29711 139
rect 28272 82 28323 136
rect 28380 132 29241 136
rect 28380 129 28998 132
rect 28380 82 28551 129
rect 28272 71 28551 82
rect 28630 128 28998 129
rect 28630 74 28796 128
rect 28853 74 28998 128
rect 29077 82 29241 132
rect 29298 85 29711 136
rect 29768 136 30622 139
rect 29768 132 30175 136
rect 29768 85 29883 132
rect 29298 82 29883 85
rect 29077 74 29883 82
rect 29962 82 30175 132
rect 30232 134 30622 136
rect 30232 82 30432 134
rect 29962 76 30432 82
rect 30511 85 30622 134
rect 30679 85 31011 139
rect 30511 76 31011 85
rect 29962 74 31011 76
rect 28630 71 31011 74
rect 28272 65 31011 71
<< viali >>
rect 5399 3787 5449 3823
rect 5817 3791 5867 3827
rect 6272 3797 6322 3833
rect 6748 3790 6804 3835
rect 7194 3795 7250 3840
rect 7639 3789 7695 3834
rect 8157 3792 8210 3843
rect 8584 3787 8637 3838
rect 9064 3787 9117 3838
rect 9414 3790 9462 3848
rect 9870 3794 9918 3852
rect 10334 3793 10382 3851
rect 10703 3787 10753 3823
rect 11121 3791 11171 3827
rect 11576 3797 11626 3833
rect 12052 3790 12108 3835
rect 12498 3795 12554 3840
rect 12943 3789 12999 3834
rect 13461 3792 13514 3843
rect 13888 3787 13941 3838
rect 14368 3787 14421 3838
rect 14718 3790 14766 3848
rect 15174 3794 15222 3852
rect 15638 3793 15686 3851
rect 15967 3787 16017 3823
rect 16385 3791 16435 3827
rect 16840 3797 16890 3833
rect 17316 3790 17372 3835
rect 17762 3795 17818 3840
rect 18207 3789 18263 3834
rect 18725 3792 18778 3843
rect 19152 3787 19205 3838
rect 19632 3787 19685 3838
rect 19982 3790 20030 3848
rect 20438 3794 20486 3852
rect 20902 3793 20950 3851
rect 21272 3787 21322 3823
rect 21690 3791 21740 3827
rect 22145 3797 22195 3833
rect 22621 3790 22677 3835
rect 23067 3795 23123 3840
rect 23512 3789 23568 3834
rect 24030 3792 24083 3843
rect 24457 3787 24510 3838
rect 24937 3787 24990 3838
rect 25287 3790 25335 3848
rect 25743 3794 25791 3852
rect 26207 3793 26255 3851
rect 26536 3787 26586 3823
rect 26954 3791 27004 3827
rect 27409 3797 27459 3833
rect 27885 3790 27941 3835
rect 28331 3795 28387 3840
rect 28776 3789 28832 3834
rect 29294 3792 29347 3843
rect 29721 3787 29774 3838
rect 30201 3787 30254 3838
rect 30551 3790 30599 3848
rect 31007 3794 31055 3852
rect 31471 3793 31519 3851
rect 5366 3680 5371 3693
rect 5371 3680 5402 3693
rect 7126 3694 7164 3704
rect 5366 3675 5402 3680
rect 5376 3510 5380 3546
rect 5380 3510 5393 3546
rect 5837 3508 5838 3544
rect 5838 3508 5854 3544
rect 5608 3353 5609 3389
rect 5609 3353 5625 3389
rect 6294 3508 6296 3544
rect 6296 3508 6311 3544
rect 6063 3353 6067 3392
rect 6067 3353 6081 3392
rect 5407 2565 5411 2580
rect 5411 2565 5591 2580
rect 5636 2565 5640 2580
rect 5640 2565 5820 2580
rect 5865 2565 5869 2580
rect 5869 2565 6049 2580
rect 6094 2565 6098 2580
rect 6098 2565 6278 2580
rect 5407 2563 5591 2565
rect 5636 2563 5820 2565
rect 5865 2563 6049 2565
rect 6094 2563 6278 2565
rect 7126 3682 7164 3694
rect 9728 3692 9761 3697
rect 8378 3681 8413 3686
rect 6788 3626 6972 3643
rect 7017 3626 7201 3643
rect 7246 3626 7430 3643
rect 7475 3626 7659 3643
rect 6754 3511 6757 3552
rect 6757 3511 6772 3552
rect 7213 3508 7215 3549
rect 7215 3508 7231 3549
rect 6983 3402 6986 3443
rect 6986 3402 7001 3443
rect 7670 3508 7673 3549
rect 7673 3508 7688 3549
rect 7447 3399 7461 3440
rect 7461 3399 7465 3440
rect 8378 3664 8413 3681
rect 8378 3663 8413 3664
rect 8196 3613 8380 3630
rect 8425 3613 8609 3630
rect 8654 3613 8838 3630
rect 8883 3613 9067 3630
rect 8164 3503 8165 3549
rect 8165 3503 8182 3549
rect 8182 3503 8189 3549
rect 8624 3504 8640 3547
rect 8640 3504 8644 3547
rect 8395 3360 8411 3403
rect 8411 3360 8415 3403
rect 9080 3508 9081 3551
rect 9081 3508 9098 3551
rect 9098 3508 9100 3551
rect 8853 3360 8869 3403
rect 8869 3360 8873 3403
rect 9728 3675 9761 3692
rect 9429 3505 9444 3536
rect 9444 3505 9447 3536
rect 9890 3504 9902 3550
rect 9902 3504 9909 3550
rect 9646 3307 9656 3360
rect 9656 3307 9673 3360
rect 9673 3307 9680 3360
rect 10344 3509 10360 3555
rect 10360 3509 10363 3555
rect 10107 3311 10114 3364
rect 10114 3311 10131 3364
rect 10131 3311 10141 3364
rect 9458 2560 9642 2577
rect 9687 2560 9871 2577
rect 9916 2560 10100 2577
rect 10145 2560 10329 2577
rect 10670 3680 10675 3693
rect 10675 3680 10706 3693
rect 12430 3694 12468 3704
rect 10670 3675 10706 3680
rect 10680 3510 10684 3546
rect 10684 3510 10697 3546
rect 11141 3508 11142 3544
rect 11142 3508 11158 3544
rect 10912 3353 10913 3389
rect 10913 3353 10929 3389
rect 11598 3508 11600 3544
rect 11600 3508 11615 3544
rect 11367 3353 11371 3392
rect 11371 3353 11385 3392
rect 10711 2565 10715 2580
rect 10715 2565 10895 2580
rect 10940 2565 10944 2580
rect 10944 2565 11124 2580
rect 11169 2565 11173 2580
rect 11173 2565 11353 2580
rect 11398 2565 11402 2580
rect 11402 2565 11582 2580
rect 10711 2563 10895 2565
rect 10940 2563 11124 2565
rect 11169 2563 11353 2565
rect 11398 2563 11582 2565
rect 12430 3682 12468 3694
rect 15032 3692 15065 3697
rect 13682 3681 13717 3686
rect 12092 3626 12276 3643
rect 12321 3626 12505 3643
rect 12550 3626 12734 3643
rect 12779 3626 12963 3643
rect 12058 3511 12061 3552
rect 12061 3511 12076 3552
rect 12517 3508 12519 3549
rect 12519 3508 12535 3549
rect 12287 3402 12290 3443
rect 12290 3402 12305 3443
rect 12974 3508 12977 3549
rect 12977 3508 12992 3549
rect 12751 3399 12765 3440
rect 12765 3399 12769 3440
rect 13682 3664 13717 3681
rect 13682 3663 13717 3664
rect 13500 3613 13684 3630
rect 13729 3613 13913 3630
rect 13958 3613 14142 3630
rect 14187 3613 14371 3630
rect 13468 3503 13469 3549
rect 13469 3503 13486 3549
rect 13486 3503 13493 3549
rect 13928 3504 13944 3547
rect 13944 3504 13948 3547
rect 13699 3360 13715 3403
rect 13715 3360 13719 3403
rect 14384 3508 14385 3551
rect 14385 3508 14402 3551
rect 14402 3508 14404 3551
rect 14157 3360 14173 3403
rect 14173 3360 14177 3403
rect 15032 3675 15065 3692
rect 14733 3505 14748 3536
rect 14748 3505 14751 3536
rect 15194 3504 15206 3550
rect 15206 3504 15213 3550
rect 14950 3307 14960 3360
rect 14960 3307 14977 3360
rect 14977 3307 14984 3360
rect 15648 3509 15664 3555
rect 15664 3509 15667 3555
rect 15411 3311 15418 3364
rect 15418 3311 15435 3364
rect 15435 3311 15445 3364
rect 14762 2560 14946 2577
rect 14991 2560 15175 2577
rect 15220 2560 15404 2577
rect 15449 2560 15633 2577
rect 15934 3680 15939 3693
rect 15939 3680 15970 3693
rect 17694 3694 17732 3704
rect 15934 3675 15970 3680
rect 15944 3510 15948 3546
rect 15948 3510 15961 3546
rect 16405 3508 16406 3544
rect 16406 3508 16422 3544
rect 16176 3353 16177 3389
rect 16177 3353 16193 3389
rect 16862 3508 16864 3544
rect 16864 3508 16879 3544
rect 16631 3353 16635 3392
rect 16635 3353 16649 3392
rect 15975 2565 15979 2580
rect 15979 2565 16159 2580
rect 16204 2565 16208 2580
rect 16208 2565 16388 2580
rect 16433 2565 16437 2580
rect 16437 2565 16617 2580
rect 16662 2565 16666 2580
rect 16666 2565 16846 2580
rect 15975 2563 16159 2565
rect 16204 2563 16388 2565
rect 16433 2563 16617 2565
rect 16662 2563 16846 2565
rect 17694 3682 17732 3694
rect 20296 3692 20329 3697
rect 18946 3681 18981 3686
rect 17356 3626 17540 3643
rect 17585 3626 17769 3643
rect 17814 3626 17998 3643
rect 18043 3626 18227 3643
rect 17322 3511 17325 3552
rect 17325 3511 17340 3552
rect 17781 3508 17783 3549
rect 17783 3508 17799 3549
rect 17551 3402 17554 3443
rect 17554 3402 17569 3443
rect 18238 3508 18241 3549
rect 18241 3508 18256 3549
rect 18015 3399 18029 3440
rect 18029 3399 18033 3440
rect 18946 3664 18981 3681
rect 18946 3663 18981 3664
rect 18764 3613 18948 3630
rect 18993 3613 19177 3630
rect 19222 3613 19406 3630
rect 19451 3613 19635 3630
rect 18732 3503 18733 3549
rect 18733 3503 18750 3549
rect 18750 3503 18757 3549
rect 19192 3504 19208 3547
rect 19208 3504 19212 3547
rect 18963 3360 18979 3403
rect 18979 3360 18983 3403
rect 19648 3508 19649 3551
rect 19649 3508 19666 3551
rect 19666 3508 19668 3551
rect 19421 3360 19437 3403
rect 19437 3360 19441 3403
rect 20296 3675 20329 3692
rect 19997 3505 20012 3536
rect 20012 3505 20015 3536
rect 20458 3504 20470 3550
rect 20470 3504 20477 3550
rect 20214 3307 20224 3360
rect 20224 3307 20241 3360
rect 20241 3307 20248 3360
rect 20912 3509 20928 3555
rect 20928 3509 20931 3555
rect 20675 3311 20682 3364
rect 20682 3311 20699 3364
rect 20699 3311 20709 3364
rect 20026 2560 20210 2577
rect 20255 2560 20439 2577
rect 20484 2560 20668 2577
rect 20713 2560 20897 2577
rect 21239 3680 21244 3693
rect 21244 3680 21275 3693
rect 22999 3694 23037 3704
rect 21239 3675 21275 3680
rect 21249 3510 21253 3546
rect 21253 3510 21266 3546
rect 21710 3508 21711 3544
rect 21711 3508 21727 3544
rect 21481 3353 21482 3389
rect 21482 3353 21498 3389
rect 22167 3508 22169 3544
rect 22169 3508 22184 3544
rect 21936 3353 21940 3392
rect 21940 3353 21954 3392
rect 21280 2565 21284 2580
rect 21284 2565 21464 2580
rect 21509 2565 21513 2580
rect 21513 2565 21693 2580
rect 21738 2565 21742 2580
rect 21742 2565 21922 2580
rect 21967 2565 21971 2580
rect 21971 2565 22151 2580
rect 21280 2563 21464 2565
rect 21509 2563 21693 2565
rect 21738 2563 21922 2565
rect 21967 2563 22151 2565
rect 22999 3682 23037 3694
rect 25601 3692 25634 3697
rect 24251 3681 24286 3686
rect 22661 3626 22845 3643
rect 22890 3626 23074 3643
rect 23119 3626 23303 3643
rect 23348 3626 23532 3643
rect 22627 3511 22630 3552
rect 22630 3511 22645 3552
rect 23086 3508 23088 3549
rect 23088 3508 23104 3549
rect 22856 3402 22859 3443
rect 22859 3402 22874 3443
rect 23543 3508 23546 3549
rect 23546 3508 23561 3549
rect 23320 3399 23334 3440
rect 23334 3399 23338 3440
rect 24251 3664 24286 3681
rect 24251 3663 24286 3664
rect 24069 3613 24253 3630
rect 24298 3613 24482 3630
rect 24527 3613 24711 3630
rect 24756 3613 24940 3630
rect 24037 3503 24038 3549
rect 24038 3503 24055 3549
rect 24055 3503 24062 3549
rect 24497 3504 24513 3547
rect 24513 3504 24517 3547
rect 24268 3360 24284 3403
rect 24284 3360 24288 3403
rect 24953 3508 24954 3551
rect 24954 3508 24971 3551
rect 24971 3508 24973 3551
rect 24726 3360 24742 3403
rect 24742 3360 24746 3403
rect 25601 3675 25634 3692
rect 25302 3505 25317 3536
rect 25317 3505 25320 3536
rect 25763 3504 25775 3550
rect 25775 3504 25782 3550
rect 25519 3307 25529 3360
rect 25529 3307 25546 3360
rect 25546 3307 25553 3360
rect 26217 3509 26233 3555
rect 26233 3509 26236 3555
rect 25980 3311 25987 3364
rect 25987 3311 26004 3364
rect 26004 3311 26014 3364
rect 25331 2560 25515 2577
rect 25560 2560 25744 2577
rect 25789 2560 25973 2577
rect 26018 2560 26202 2577
rect 26503 3680 26508 3693
rect 26508 3680 26539 3693
rect 28263 3694 28301 3704
rect 26503 3675 26539 3680
rect 26513 3510 26517 3546
rect 26517 3510 26530 3546
rect 26974 3508 26975 3544
rect 26975 3508 26991 3544
rect 26745 3353 26746 3389
rect 26746 3353 26762 3389
rect 27431 3508 27433 3544
rect 27433 3508 27448 3544
rect 27200 3353 27204 3392
rect 27204 3353 27218 3392
rect 26544 2565 26548 2580
rect 26548 2565 26728 2580
rect 26773 2565 26777 2580
rect 26777 2565 26957 2580
rect 27002 2565 27006 2580
rect 27006 2565 27186 2580
rect 27231 2565 27235 2580
rect 27235 2565 27415 2580
rect 26544 2563 26728 2565
rect 26773 2563 26957 2565
rect 27002 2563 27186 2565
rect 27231 2563 27415 2565
rect 28263 3682 28301 3694
rect 30865 3692 30898 3697
rect 29515 3681 29550 3686
rect 27925 3626 28109 3643
rect 28154 3626 28338 3643
rect 28383 3626 28567 3643
rect 28612 3626 28796 3643
rect 27891 3511 27894 3552
rect 27894 3511 27909 3552
rect 28350 3508 28352 3549
rect 28352 3508 28368 3549
rect 28120 3402 28123 3443
rect 28123 3402 28138 3443
rect 28807 3508 28810 3549
rect 28810 3508 28825 3549
rect 28584 3399 28598 3440
rect 28598 3399 28602 3440
rect 29515 3664 29550 3681
rect 29515 3663 29550 3664
rect 29333 3613 29517 3630
rect 29562 3613 29746 3630
rect 29791 3613 29975 3630
rect 30020 3613 30204 3630
rect 29301 3503 29302 3549
rect 29302 3503 29319 3549
rect 29319 3503 29326 3549
rect 29761 3504 29777 3547
rect 29777 3504 29781 3547
rect 29532 3360 29548 3403
rect 29548 3360 29552 3403
rect 30217 3508 30218 3551
rect 30218 3508 30235 3551
rect 30235 3508 30237 3551
rect 29990 3360 30006 3403
rect 30006 3360 30010 3403
rect 30865 3675 30898 3692
rect 30566 3505 30581 3536
rect 30581 3505 30584 3536
rect 31027 3504 31039 3550
rect 31039 3504 31046 3550
rect 30783 3307 30793 3360
rect 30793 3307 30810 3360
rect 30810 3307 30817 3360
rect 31481 3509 31497 3555
rect 31497 3509 31500 3555
rect 31244 3311 31251 3364
rect 31251 3311 31268 3364
rect 31268 3311 31278 3364
rect 30595 2560 30779 2577
rect 30824 2560 31008 2577
rect 31053 2560 31237 2577
rect 31282 2560 31466 2577
rect 6492 2061 6562 2065
rect 6492 2047 6562 2061
rect 6004 2022 6021 2039
rect 6509 2000 6562 2017
rect 6509 1994 6562 2000
rect 6505 1960 6558 1963
rect 6505 1943 6558 1960
rect 9236 2066 9278 2071
rect 9236 2051 9278 2066
rect 9784 2027 9801 2044
rect 9236 2022 9276 2023
rect 9236 2005 9276 2022
rect 9236 2003 9276 2005
rect 9237 1965 9277 1970
rect 9237 1950 9277 1965
rect 11796 2061 11866 2065
rect 11796 2047 11866 2061
rect 11308 2022 11325 2039
rect 11813 2000 11866 2017
rect 11813 1994 11866 2000
rect 11809 1960 11862 1963
rect 11809 1943 11862 1960
rect 14540 2066 14582 2071
rect 14540 2051 14582 2066
rect 15088 2027 15105 2044
rect 14540 2022 14580 2023
rect 14540 2005 14580 2022
rect 14540 2003 14580 2005
rect 14541 1965 14581 1970
rect 14541 1950 14581 1965
rect 17060 2061 17130 2065
rect 17060 2047 17130 2061
rect 16572 2022 16589 2039
rect 17077 2000 17130 2017
rect 17077 1994 17130 2000
rect 17073 1960 17126 1963
rect 17073 1943 17126 1960
rect 19804 2066 19846 2071
rect 19804 2051 19846 2066
rect 20352 2027 20369 2044
rect 19804 2022 19844 2023
rect 19804 2005 19844 2022
rect 19804 2003 19844 2005
rect 19805 1965 19845 1970
rect 19805 1950 19845 1965
rect 22365 2061 22435 2065
rect 22365 2047 22435 2061
rect 21877 2022 21894 2039
rect 22382 2000 22435 2017
rect 22382 1994 22435 2000
rect 22378 1960 22431 1963
rect 22378 1943 22431 1960
rect 25109 2066 25151 2071
rect 25109 2051 25151 2066
rect 25657 2027 25674 2044
rect 25109 2022 25149 2023
rect 25109 2005 25149 2022
rect 25109 2003 25149 2005
rect 25110 1965 25150 1970
rect 25110 1950 25150 1965
rect 27629 2061 27699 2065
rect 27629 2047 27699 2061
rect 27141 2022 27158 2039
rect 27646 2000 27699 2017
rect 27646 1994 27699 2000
rect 27642 1960 27695 1963
rect 27642 1943 27695 1960
rect 30373 2066 30415 2071
rect 30373 2051 30415 2066
rect 30921 2027 30938 2044
rect 30373 2022 30413 2023
rect 30373 2005 30413 2022
rect 30373 2003 30413 2005
rect 30374 1965 30414 1970
rect 30374 1950 30414 1965
rect 6505 1940 6558 1943
rect 11809 1940 11862 1943
rect 17073 1940 17126 1943
rect 22378 1940 22431 1943
rect 27642 1940 27695 1943
rect 7211 1431 7214 1479
rect 7214 1431 7231 1479
rect 7231 1431 7235 1479
rect 7669 1427 7672 1475
rect 7672 1427 7689 1475
rect 7689 1427 7693 1475
rect 7427 1323 7443 1378
rect 7443 1323 7460 1378
rect 7460 1323 7462 1378
rect 8128 1433 8130 1481
rect 8130 1433 8147 1481
rect 8147 1433 8152 1481
rect 7889 1329 7901 1384
rect 7901 1329 7918 1384
rect 7918 1329 7924 1384
rect 8582 1437 8588 1485
rect 8588 1437 8605 1485
rect 8605 1437 8606 1485
rect 8348 1335 8359 1390
rect 8359 1335 8376 1390
rect 8376 1335 8383 1390
rect 9035 1434 9046 1482
rect 9046 1434 9059 1482
rect 8810 1335 8817 1390
rect 8817 1335 8834 1390
rect 8834 1335 8845 1390
rect 9501 1434 9504 1482
rect 9504 1434 9521 1482
rect 9521 1434 9525 1482
rect 9272 1329 9275 1384
rect 9275 1329 9292 1384
rect 9292 1329 9307 1384
rect 9720 1338 9733 1393
rect 9733 1338 9750 1393
rect 9750 1338 9755 1393
rect 7245 290 7429 307
rect 7474 290 7658 307
rect 7703 290 7887 307
rect 7932 290 8116 307
rect 8161 290 8345 307
rect 8390 290 8574 307
rect 8619 290 8803 307
rect 8848 290 9032 307
rect 9077 290 9261 307
rect 9306 290 9490 307
rect 9535 290 9719 307
rect 9172 239 9223 252
rect 12515 1431 12518 1479
rect 12518 1431 12535 1479
rect 12535 1431 12539 1479
rect 12973 1427 12976 1475
rect 12976 1427 12993 1475
rect 12993 1427 12997 1475
rect 12731 1323 12747 1378
rect 12747 1323 12764 1378
rect 12764 1323 12766 1378
rect 13432 1433 13434 1481
rect 13434 1433 13451 1481
rect 13451 1433 13456 1481
rect 13193 1329 13205 1384
rect 13205 1329 13222 1384
rect 13222 1329 13228 1384
rect 13886 1437 13892 1485
rect 13892 1437 13909 1485
rect 13909 1437 13910 1485
rect 13652 1335 13663 1390
rect 13663 1335 13680 1390
rect 13680 1335 13687 1390
rect 14339 1434 14350 1482
rect 14350 1434 14363 1482
rect 14114 1335 14121 1390
rect 14121 1335 14138 1390
rect 14138 1335 14149 1390
rect 14805 1434 14808 1482
rect 14808 1434 14825 1482
rect 14825 1434 14829 1482
rect 14576 1329 14579 1384
rect 14579 1329 14596 1384
rect 14596 1329 14611 1384
rect 15024 1338 15037 1393
rect 15037 1338 15054 1393
rect 15054 1338 15059 1393
rect 12549 290 12733 307
rect 12778 290 12962 307
rect 13007 290 13191 307
rect 13236 290 13420 307
rect 13465 290 13649 307
rect 13694 290 13878 307
rect 13923 290 14107 307
rect 14152 290 14336 307
rect 14381 290 14565 307
rect 14610 290 14794 307
rect 14839 290 15023 307
rect 14476 239 14527 252
rect 17779 1431 17782 1479
rect 17782 1431 17799 1479
rect 17799 1431 17803 1479
rect 18237 1427 18240 1475
rect 18240 1427 18257 1475
rect 18257 1427 18261 1475
rect 17995 1323 18011 1378
rect 18011 1323 18028 1378
rect 18028 1323 18030 1378
rect 18696 1433 18698 1481
rect 18698 1433 18715 1481
rect 18715 1433 18720 1481
rect 18457 1329 18469 1384
rect 18469 1329 18486 1384
rect 18486 1329 18492 1384
rect 19150 1437 19156 1485
rect 19156 1437 19173 1485
rect 19173 1437 19174 1485
rect 18916 1335 18927 1390
rect 18927 1335 18944 1390
rect 18944 1335 18951 1390
rect 19603 1434 19614 1482
rect 19614 1434 19627 1482
rect 19378 1335 19385 1390
rect 19385 1335 19402 1390
rect 19402 1335 19413 1390
rect 20069 1434 20072 1482
rect 20072 1434 20089 1482
rect 20089 1434 20093 1482
rect 19840 1329 19843 1384
rect 19843 1329 19860 1384
rect 19860 1329 19875 1384
rect 20288 1338 20301 1393
rect 20301 1338 20318 1393
rect 20318 1338 20323 1393
rect 17813 290 17997 307
rect 18042 290 18226 307
rect 18271 290 18455 307
rect 18500 290 18684 307
rect 18729 290 18913 307
rect 18958 290 19142 307
rect 19187 290 19371 307
rect 19416 290 19600 307
rect 19645 290 19829 307
rect 19874 290 20058 307
rect 20103 290 20287 307
rect 19740 239 19791 252
rect 23084 1431 23087 1479
rect 23087 1431 23104 1479
rect 23104 1431 23108 1479
rect 23542 1427 23545 1475
rect 23545 1427 23562 1475
rect 23562 1427 23566 1475
rect 23300 1323 23316 1378
rect 23316 1323 23333 1378
rect 23333 1323 23335 1378
rect 24001 1433 24003 1481
rect 24003 1433 24020 1481
rect 24020 1433 24025 1481
rect 23762 1329 23774 1384
rect 23774 1329 23791 1384
rect 23791 1329 23797 1384
rect 24455 1437 24461 1485
rect 24461 1437 24478 1485
rect 24478 1437 24479 1485
rect 24221 1335 24232 1390
rect 24232 1335 24249 1390
rect 24249 1335 24256 1390
rect 24908 1434 24919 1482
rect 24919 1434 24932 1482
rect 24683 1335 24690 1390
rect 24690 1335 24707 1390
rect 24707 1335 24718 1390
rect 25374 1434 25377 1482
rect 25377 1434 25394 1482
rect 25394 1434 25398 1482
rect 25145 1329 25148 1384
rect 25148 1329 25165 1384
rect 25165 1329 25180 1384
rect 25593 1338 25606 1393
rect 25606 1338 25623 1393
rect 25623 1338 25628 1393
rect 23118 290 23302 307
rect 23347 290 23531 307
rect 23576 290 23760 307
rect 23805 290 23989 307
rect 24034 290 24218 307
rect 24263 290 24447 307
rect 24492 290 24676 307
rect 24721 290 24905 307
rect 24950 290 25134 307
rect 25179 290 25363 307
rect 25408 290 25592 307
rect 25045 239 25096 252
rect 28348 1431 28351 1479
rect 28351 1431 28368 1479
rect 28368 1431 28372 1479
rect 28806 1427 28809 1475
rect 28809 1427 28826 1475
rect 28826 1427 28830 1475
rect 28564 1323 28580 1378
rect 28580 1323 28597 1378
rect 28597 1323 28599 1378
rect 29265 1433 29267 1481
rect 29267 1433 29284 1481
rect 29284 1433 29289 1481
rect 29026 1329 29038 1384
rect 29038 1329 29055 1384
rect 29055 1329 29061 1384
rect 29719 1437 29725 1485
rect 29725 1437 29742 1485
rect 29742 1437 29743 1485
rect 29485 1335 29496 1390
rect 29496 1335 29513 1390
rect 29513 1335 29520 1390
rect 30172 1434 30183 1482
rect 30183 1434 30196 1482
rect 29947 1335 29954 1390
rect 29954 1335 29971 1390
rect 29971 1335 29982 1390
rect 30638 1434 30641 1482
rect 30641 1434 30658 1482
rect 30658 1434 30662 1482
rect 30409 1329 30412 1384
rect 30412 1329 30429 1384
rect 30429 1329 30444 1384
rect 30857 1338 30870 1393
rect 30870 1338 30887 1393
rect 30887 1338 30892 1393
rect 28382 290 28566 307
rect 28611 290 28795 307
rect 28840 290 29024 307
rect 29069 290 29253 307
rect 29298 290 29482 307
rect 29527 290 29711 307
rect 29756 290 29940 307
rect 29985 290 30169 307
rect 30214 290 30398 307
rect 30443 290 30627 307
rect 30672 290 30856 307
rect 30309 239 30360 252
rect 9172 235 9223 239
rect 14476 235 14527 239
rect 19740 235 19791 239
rect 25045 235 25096 239
rect 30309 235 30360 239
rect 7186 82 7243 136
rect 7659 74 7716 128
rect 8104 82 8161 136
rect 8574 85 8631 139
rect 9038 82 9095 136
rect 9485 85 9542 139
rect 12490 82 12547 136
rect 12963 74 13020 128
rect 13408 82 13465 136
rect 13878 85 13935 139
rect 14342 82 14399 136
rect 14789 85 14846 139
rect 17754 82 17811 136
rect 18227 74 18284 128
rect 18672 82 18729 136
rect 19142 85 19199 139
rect 19606 82 19663 136
rect 20053 85 20110 139
rect 23059 82 23116 136
rect 23532 74 23589 128
rect 23977 82 24034 136
rect 24447 85 24504 139
rect 24911 82 24968 136
rect 25358 85 25415 139
rect 28323 82 28380 136
rect 28796 74 28853 128
rect 29241 82 29298 136
rect 29711 85 29768 139
rect 30175 82 30232 136
rect 30622 85 30679 139
<< metal1 >>
rect 1528 4000 5744 4235
rect 1528 3852 31632 4000
rect 1528 3848 9870 3852
rect 1528 3843 8160 3848
rect 8187 3843 9414 3848
rect 1528 3840 8157 3843
rect 1528 3835 7194 3840
rect 1528 3833 6748 3835
rect 1528 3827 6272 3833
rect 1528 3823 5817 3827
rect 1528 3787 5399 3823
rect 5449 3791 5817 3823
rect 5867 3797 6272 3827
rect 6322 3797 6748 3833
rect 5867 3791 6748 3797
rect 5449 3790 6748 3791
rect 6804 3795 7194 3835
rect 7250 3834 8157 3840
rect 7250 3795 7639 3834
rect 6804 3790 7639 3795
rect 5449 3789 7639 3790
rect 7695 3792 8157 3834
rect 8210 3838 9414 3843
rect 8210 3792 8584 3838
rect 7695 3789 8584 3792
rect 5449 3787 8584 3789
rect 8637 3787 9064 3838
rect 9117 3790 9414 3838
rect 9462 3794 9870 3848
rect 9918 3851 15174 3852
rect 9918 3794 10334 3851
rect 9462 3793 10334 3794
rect 10382 3848 15174 3851
rect 10382 3843 13464 3848
rect 13491 3843 14718 3848
rect 10382 3840 13461 3843
rect 10382 3835 12498 3840
rect 10382 3833 12052 3835
rect 10382 3827 11576 3833
rect 10382 3823 11121 3827
rect 10382 3793 10703 3823
rect 9462 3790 10703 3793
rect 9117 3787 10703 3790
rect 10753 3791 11121 3823
rect 11171 3797 11576 3827
rect 11626 3797 12052 3833
rect 11171 3791 12052 3797
rect 10753 3790 12052 3791
rect 12108 3795 12498 3835
rect 12554 3834 13461 3840
rect 12554 3795 12943 3834
rect 12108 3790 12943 3795
rect 10753 3789 12943 3790
rect 12999 3792 13461 3834
rect 13514 3838 14718 3843
rect 13514 3792 13888 3838
rect 12999 3789 13888 3792
rect 10753 3787 13888 3789
rect 13941 3787 14368 3838
rect 14421 3790 14718 3838
rect 14766 3794 15174 3848
rect 15222 3851 20438 3852
rect 15222 3794 15638 3851
rect 14766 3793 15638 3794
rect 15686 3848 20438 3851
rect 15686 3843 18728 3848
rect 18755 3843 19982 3848
rect 15686 3840 18725 3843
rect 15686 3835 17762 3840
rect 15686 3833 17316 3835
rect 15686 3827 16840 3833
rect 15686 3823 16385 3827
rect 15686 3793 15967 3823
rect 14766 3790 15967 3793
rect 14421 3787 15967 3790
rect 16017 3791 16385 3823
rect 16435 3797 16840 3827
rect 16890 3797 17316 3833
rect 16435 3791 17316 3797
rect 16017 3790 17316 3791
rect 17372 3795 17762 3835
rect 17818 3834 18725 3840
rect 17818 3795 18207 3834
rect 17372 3790 18207 3795
rect 16017 3789 18207 3790
rect 18263 3792 18725 3834
rect 18778 3838 19982 3843
rect 18778 3792 19152 3838
rect 18263 3789 19152 3792
rect 16017 3787 19152 3789
rect 19205 3787 19632 3838
rect 19685 3790 19982 3838
rect 20030 3794 20438 3848
rect 20486 3851 25743 3852
rect 20486 3794 20902 3851
rect 20030 3793 20902 3794
rect 20950 3848 25743 3851
rect 20950 3843 24033 3848
rect 24060 3843 25287 3848
rect 20950 3840 24030 3843
rect 20950 3835 23067 3840
rect 20950 3833 22621 3835
rect 20950 3827 22145 3833
rect 20950 3823 21690 3827
rect 20950 3793 21272 3823
rect 20030 3790 21272 3793
rect 19685 3787 21272 3790
rect 21322 3791 21690 3823
rect 21740 3797 22145 3827
rect 22195 3797 22621 3833
rect 21740 3791 22621 3797
rect 21322 3790 22621 3791
rect 22677 3795 23067 3835
rect 23123 3834 24030 3840
rect 23123 3795 23512 3834
rect 22677 3790 23512 3795
rect 21322 3789 23512 3790
rect 23568 3792 24030 3834
rect 24083 3838 25287 3843
rect 24083 3792 24457 3838
rect 23568 3789 24457 3792
rect 21322 3787 24457 3789
rect 24510 3787 24937 3838
rect 24990 3790 25287 3838
rect 25335 3794 25743 3848
rect 25791 3851 31007 3852
rect 25791 3794 26207 3851
rect 25335 3793 26207 3794
rect 26255 3848 31007 3851
rect 26255 3843 29297 3848
rect 29324 3843 30551 3848
rect 26255 3840 29294 3843
rect 26255 3835 28331 3840
rect 26255 3833 27885 3835
rect 26255 3827 27409 3833
rect 26255 3823 26954 3827
rect 26255 3793 26536 3823
rect 25335 3790 26536 3793
rect 24990 3787 26536 3790
rect 26586 3791 26954 3823
rect 27004 3797 27409 3827
rect 27459 3797 27885 3833
rect 27004 3791 27885 3797
rect 26586 3790 27885 3791
rect 27941 3795 28331 3835
rect 28387 3834 29294 3840
rect 28387 3795 28776 3834
rect 27941 3790 28776 3795
rect 26586 3789 28776 3790
rect 28832 3792 29294 3834
rect 29347 3838 30551 3843
rect 29347 3792 29721 3838
rect 28832 3789 29721 3792
rect 26586 3787 29721 3789
rect 29774 3787 30201 3838
rect 30254 3790 30551 3838
rect 30599 3794 31007 3848
rect 31055 3851 31632 3852
rect 31055 3794 31471 3851
rect 30599 3793 31471 3794
rect 31519 3793 31632 3851
rect 30599 3790 31632 3793
rect 30254 3787 31632 3790
rect 1528 3761 31632 3787
rect 5274 3755 31632 3761
rect 5352 3693 5411 3755
rect 5352 3675 5366 3693
rect 5402 3675 5411 3693
rect 5352 3551 5411 3675
rect 7119 3704 7172 3755
rect 7119 3682 7126 3704
rect 7164 3682 7172 3704
rect 7119 3673 7172 3682
rect 8368 3686 8431 3755
rect 7861 3657 8005 3675
rect 8368 3663 8378 3686
rect 8413 3663 8431 3686
rect 8368 3659 8431 3663
rect 6768 3652 8172 3657
rect 6768 3643 7882 3652
rect 6768 3626 6788 3643
rect 6972 3626 7017 3643
rect 7201 3626 7246 3643
rect 7430 3626 7475 3643
rect 7659 3626 7882 3643
rect 6768 3610 7882 3626
rect 7757 3597 7882 3610
rect 7861 3592 7882 3597
rect 7986 3639 8172 3652
rect 7986 3630 9098 3639
rect 7986 3613 8196 3630
rect 8380 3613 8425 3630
rect 8609 3613 8654 3630
rect 8838 3613 8883 3630
rect 9067 3613 9098 3630
rect 7986 3597 9098 3613
rect 7986 3592 8005 3597
rect 7861 3571 8005 3592
rect 9418 3561 9459 3755
rect 9721 3750 10495 3755
rect 9721 3697 9770 3750
rect 9721 3675 9728 3697
rect 9761 3675 9770 3697
rect 9721 3668 9770 3675
rect 10656 3693 10715 3755
rect 10656 3675 10670 3693
rect 10706 3675 10715 3693
rect 6735 3552 7711 3559
rect 6047 3551 6192 3552
rect 5352 3546 6329 3551
rect 5352 3510 5376 3546
rect 5393 3544 6329 3546
rect 5393 3510 5837 3544
rect 5352 3508 5837 3510
rect 5854 3508 6294 3544
rect 6311 3508 6329 3544
rect 5352 3507 6329 3508
rect 5352 3503 6098 3507
rect 6140 3503 6329 3507
rect 6735 3547 6754 3552
rect 6772 3549 7711 3552
rect 6772 3547 7213 3549
rect 6735 3501 6750 3547
rect 6803 3508 7213 3547
rect 7231 3508 7670 3549
rect 7688 3508 7711 3549
rect 6803 3501 7711 3508
rect 6735 3494 7711 3501
rect 8145 3551 9126 3559
rect 8145 3549 9080 3551
rect 8145 3544 8164 3549
rect 8189 3547 9080 3549
rect 8145 3499 8159 3544
rect 8189 3504 8624 3547
rect 8644 3508 9080 3547
rect 9100 3508 9126 3551
rect 8644 3504 9126 3508
rect 8189 3503 9126 3504
rect 8186 3499 9126 3503
rect 8145 3493 9126 3499
rect 9416 3555 10372 3561
rect 9416 3550 10344 3555
rect 9416 3536 9890 3550
rect 9416 3505 9429 3536
rect 9447 3505 9890 3536
rect 9416 3504 9890 3505
rect 9909 3509 10344 3550
rect 10363 3509 10372 3555
rect 9909 3504 10372 3509
rect 9416 3485 10372 3504
rect 10656 3551 10715 3675
rect 12423 3704 12476 3755
rect 12423 3682 12430 3704
rect 12468 3682 12476 3704
rect 12423 3673 12476 3682
rect 13672 3686 13735 3755
rect 13166 3657 13310 3673
rect 13672 3663 13682 3686
rect 13717 3663 13735 3686
rect 13672 3659 13735 3663
rect 12072 3649 13476 3657
rect 12072 3643 13187 3649
rect 12072 3626 12092 3643
rect 12276 3626 12321 3643
rect 12505 3626 12550 3643
rect 12734 3626 12779 3643
rect 12963 3626 13187 3643
rect 12072 3610 13187 3626
rect 13061 3597 13187 3610
rect 13166 3590 13187 3597
rect 13291 3639 13476 3649
rect 13291 3630 14402 3639
rect 13291 3613 13500 3630
rect 13684 3613 13729 3630
rect 13913 3613 13958 3630
rect 14142 3613 14187 3630
rect 14371 3613 14402 3630
rect 13291 3597 14402 3613
rect 13291 3590 13310 3597
rect 13166 3568 13310 3590
rect 14722 3561 14763 3755
rect 15025 3750 15799 3755
rect 15025 3697 15074 3750
rect 15025 3675 15032 3697
rect 15065 3675 15074 3697
rect 15025 3668 15074 3675
rect 15920 3693 15979 3755
rect 15920 3675 15934 3693
rect 15970 3675 15979 3693
rect 12039 3552 13015 3559
rect 11351 3551 11496 3552
rect 10656 3546 11633 3551
rect 10656 3510 10680 3546
rect 10697 3544 11633 3546
rect 10697 3510 11141 3544
rect 10656 3508 11141 3510
rect 11158 3508 11598 3544
rect 11615 3508 11633 3544
rect 10656 3507 11633 3508
rect 10656 3503 11402 3507
rect 11444 3503 11633 3507
rect 12039 3547 12058 3552
rect 12076 3549 13015 3552
rect 12076 3547 12517 3549
rect 12039 3501 12054 3547
rect 12107 3508 12517 3547
rect 12535 3508 12974 3549
rect 12992 3508 13015 3549
rect 12107 3501 13015 3508
rect 12039 3494 13015 3501
rect 13449 3551 14430 3559
rect 13449 3549 14384 3551
rect 13449 3544 13468 3549
rect 13493 3547 14384 3549
rect 13449 3499 13463 3544
rect 13493 3504 13928 3547
rect 13948 3508 14384 3547
rect 14404 3508 14430 3551
rect 13948 3504 14430 3508
rect 13493 3503 14430 3504
rect 13490 3499 14430 3503
rect 13449 3493 14430 3499
rect 14720 3555 15676 3561
rect 14720 3550 15648 3555
rect 14720 3536 15194 3550
rect 14720 3505 14733 3536
rect 14751 3505 15194 3536
rect 14720 3504 15194 3505
rect 15213 3509 15648 3550
rect 15667 3509 15676 3555
rect 15213 3504 15676 3509
rect 14720 3485 15676 3504
rect 15920 3551 15979 3675
rect 17687 3704 17740 3755
rect 17687 3682 17694 3704
rect 17732 3682 17740 3704
rect 17687 3673 17740 3682
rect 18936 3686 18999 3755
rect 18430 3657 18575 3673
rect 18936 3663 18946 3686
rect 18981 3663 18999 3686
rect 18936 3659 18999 3663
rect 17336 3649 18740 3657
rect 17336 3643 18452 3649
rect 17336 3626 17356 3643
rect 17540 3626 17585 3643
rect 17769 3626 17814 3643
rect 17998 3626 18043 3643
rect 18227 3626 18452 3643
rect 17336 3610 18452 3626
rect 18325 3597 18452 3610
rect 18430 3590 18452 3597
rect 18555 3639 18740 3649
rect 18555 3630 19666 3639
rect 18555 3613 18764 3630
rect 18948 3613 18993 3630
rect 19177 3613 19222 3630
rect 19406 3613 19451 3630
rect 19635 3613 19666 3630
rect 18555 3597 19666 3613
rect 18555 3590 18575 3597
rect 18430 3568 18575 3590
rect 19986 3561 20027 3755
rect 20289 3750 21063 3755
rect 20289 3697 20338 3750
rect 20289 3675 20296 3697
rect 20329 3675 20338 3697
rect 20289 3668 20338 3675
rect 21225 3693 21284 3755
rect 21225 3675 21239 3693
rect 21275 3675 21284 3693
rect 17303 3552 18279 3559
rect 16615 3551 16760 3552
rect 15920 3546 16897 3551
rect 15920 3510 15944 3546
rect 15961 3544 16897 3546
rect 15961 3510 16405 3544
rect 15920 3508 16405 3510
rect 16422 3508 16862 3544
rect 16879 3508 16897 3544
rect 15920 3507 16897 3508
rect 15920 3503 16666 3507
rect 16708 3503 16897 3507
rect 17303 3547 17322 3552
rect 17340 3549 18279 3552
rect 17340 3547 17781 3549
rect 17303 3501 17318 3547
rect 17371 3508 17781 3547
rect 17799 3508 18238 3549
rect 18256 3508 18279 3549
rect 17371 3501 18279 3508
rect 17303 3494 18279 3501
rect 18713 3551 19694 3559
rect 18713 3549 19648 3551
rect 18713 3544 18732 3549
rect 18757 3547 19648 3549
rect 18713 3499 18727 3544
rect 18757 3504 19192 3547
rect 19212 3508 19648 3547
rect 19668 3508 19694 3551
rect 19212 3504 19694 3508
rect 18757 3503 19694 3504
rect 18754 3499 19694 3503
rect 18713 3493 19694 3499
rect 19984 3555 20940 3561
rect 19984 3550 20912 3555
rect 19984 3536 20458 3550
rect 19984 3505 19997 3536
rect 20015 3505 20458 3536
rect 19984 3504 20458 3505
rect 20477 3509 20912 3550
rect 20931 3509 20940 3555
rect 20477 3504 20940 3509
rect 19984 3485 20940 3504
rect 21225 3551 21284 3675
rect 22992 3704 23045 3755
rect 22992 3682 22999 3704
rect 23037 3682 23045 3704
rect 22992 3673 23045 3682
rect 24241 3686 24304 3755
rect 23722 3657 23866 3673
rect 24241 3663 24251 3686
rect 24286 3663 24304 3686
rect 24241 3659 24304 3663
rect 22641 3649 24045 3657
rect 22641 3643 23743 3649
rect 22641 3626 22661 3643
rect 22845 3626 22890 3643
rect 23074 3626 23119 3643
rect 23303 3626 23348 3643
rect 23532 3626 23743 3643
rect 22641 3610 23743 3626
rect 23630 3597 23743 3610
rect 23722 3590 23743 3597
rect 23847 3639 24045 3649
rect 23847 3630 24971 3639
rect 23847 3613 24069 3630
rect 24253 3613 24298 3630
rect 24482 3613 24527 3630
rect 24711 3613 24756 3630
rect 24940 3613 24971 3630
rect 23847 3597 24971 3613
rect 23847 3590 23866 3597
rect 23722 3568 23866 3590
rect 25291 3561 25332 3755
rect 25594 3750 26368 3755
rect 25594 3697 25643 3750
rect 25594 3675 25601 3697
rect 25634 3675 25643 3697
rect 25594 3668 25643 3675
rect 26489 3693 26548 3755
rect 26489 3675 26503 3693
rect 26539 3675 26548 3693
rect 22608 3552 23584 3559
rect 21920 3551 22065 3552
rect 21225 3546 22202 3551
rect 21225 3510 21249 3546
rect 21266 3544 22202 3546
rect 21266 3510 21710 3544
rect 21225 3508 21710 3510
rect 21727 3508 22167 3544
rect 22184 3508 22202 3544
rect 21225 3507 22202 3508
rect 21225 3503 21971 3507
rect 22013 3503 22202 3507
rect 22608 3547 22627 3552
rect 22645 3549 23584 3552
rect 22645 3547 23086 3549
rect 22608 3501 22623 3547
rect 22676 3508 23086 3547
rect 23104 3508 23543 3549
rect 23561 3508 23584 3549
rect 22676 3501 23584 3508
rect 22608 3494 23584 3501
rect 24018 3551 24999 3559
rect 24018 3549 24953 3551
rect 24018 3544 24037 3549
rect 24062 3547 24953 3549
rect 24018 3499 24032 3544
rect 24062 3504 24497 3547
rect 24517 3508 24953 3547
rect 24973 3508 24999 3551
rect 24517 3504 24999 3508
rect 24062 3503 24999 3504
rect 24059 3499 24999 3503
rect 24018 3493 24999 3499
rect 25289 3555 26245 3561
rect 25289 3550 26217 3555
rect 25289 3536 25763 3550
rect 25289 3505 25302 3536
rect 25320 3505 25763 3536
rect 25289 3504 25763 3505
rect 25782 3509 26217 3550
rect 26236 3509 26245 3555
rect 25782 3504 26245 3509
rect 25289 3485 26245 3504
rect 26489 3551 26548 3675
rect 28256 3704 28309 3755
rect 28256 3682 28263 3704
rect 28301 3682 28309 3704
rect 28256 3673 28309 3682
rect 29505 3686 29568 3755
rect 29007 3664 29151 3680
rect 29001 3657 29158 3664
rect 29505 3663 29515 3686
rect 29550 3663 29568 3686
rect 29505 3659 29568 3663
rect 27905 3656 29309 3657
rect 27905 3643 29028 3656
rect 27905 3626 27925 3643
rect 28109 3626 28154 3643
rect 28338 3626 28383 3643
rect 28567 3626 28612 3643
rect 28796 3626 29028 3643
rect 27905 3610 29028 3626
rect 28894 3597 29028 3610
rect 29132 3639 29309 3656
rect 29132 3630 30235 3639
rect 29132 3613 29333 3630
rect 29517 3613 29562 3630
rect 29746 3613 29791 3630
rect 29975 3613 30020 3630
rect 30204 3613 30235 3630
rect 29132 3597 30235 3613
rect 29007 3575 29151 3597
rect 30555 3561 30596 3755
rect 30858 3750 31632 3755
rect 30858 3697 30907 3750
rect 30858 3675 30865 3697
rect 30898 3675 30907 3697
rect 30858 3668 30907 3675
rect 27872 3552 28848 3559
rect 27184 3551 27329 3552
rect 26489 3546 27466 3551
rect 26489 3510 26513 3546
rect 26530 3544 27466 3546
rect 26530 3510 26974 3544
rect 26489 3508 26974 3510
rect 26991 3508 27431 3544
rect 27448 3508 27466 3544
rect 26489 3507 27466 3508
rect 26489 3503 27235 3507
rect 27277 3503 27466 3507
rect 27872 3547 27891 3552
rect 27909 3549 28848 3552
rect 27909 3547 28350 3549
rect 27872 3501 27887 3547
rect 27940 3508 28350 3547
rect 28368 3508 28807 3549
rect 28825 3508 28848 3549
rect 27940 3501 28848 3508
rect 27872 3494 28848 3501
rect 29282 3551 30263 3559
rect 29282 3549 30217 3551
rect 29282 3544 29301 3549
rect 29326 3547 30217 3549
rect 29282 3499 29296 3544
rect 29326 3504 29761 3547
rect 29781 3508 30217 3547
rect 30237 3508 30263 3551
rect 29781 3504 30263 3508
rect 29326 3503 30263 3504
rect 29323 3499 30263 3503
rect 29282 3493 30263 3499
rect 30553 3555 31509 3561
rect 30553 3550 31481 3555
rect 30553 3536 31027 3550
rect 30553 3505 30566 3536
rect 30584 3505 31027 3536
rect 30553 3504 31027 3505
rect 31046 3509 31481 3550
rect 31500 3509 31509 3555
rect 31046 3504 31509 3509
rect 30553 3485 31509 3504
rect 6976 3447 7472 3450
rect 12280 3447 12776 3450
rect 17544 3447 18040 3450
rect 22849 3447 23345 3450
rect 28113 3447 28609 3450
rect 6963 3443 7472 3447
rect 5580 3392 6098 3403
rect 5580 3389 6063 3392
rect 5580 3353 5608 3389
rect 5625 3353 6063 3389
rect 6081 3353 6098 3392
rect 5580 3342 6098 3353
rect 6963 3402 6983 3443
rect 7001 3440 7472 3443
rect 7001 3402 7447 3440
rect 6963 3399 7447 3402
rect 7465 3399 7472 3440
rect 12267 3443 12776 3447
rect 6963 3383 7472 3399
rect 8379 3403 8892 3417
rect 6029 2589 6095 3342
rect 5377 2580 6304 2589
rect 5377 2563 5407 2580
rect 5591 2563 5636 2580
rect 5820 2563 5865 2580
rect 6049 2563 6094 2580
rect 6278 2563 6304 2580
rect 5377 2545 6304 2563
rect 6029 2455 6095 2545
rect 6963 2455 7028 3383
rect 8379 3360 8395 3403
rect 8415 3360 8853 3403
rect 8873 3360 8892 3403
rect 10884 3392 11402 3403
rect 10884 3389 11367 3392
rect 9636 3380 10151 3382
rect 8379 3351 8892 3360
rect 9631 3364 10151 3380
rect 9631 3360 10107 3364
rect 8824 2457 8890 3351
rect 9631 3307 9646 3360
rect 9680 3311 10107 3360
rect 10141 3311 10151 3364
rect 10884 3353 10912 3389
rect 10929 3353 11367 3389
rect 11385 3353 11402 3392
rect 10884 3342 11402 3353
rect 12267 3402 12287 3443
rect 12305 3440 12776 3443
rect 12305 3402 12751 3440
rect 12267 3399 12751 3402
rect 12769 3399 12776 3440
rect 17531 3443 18040 3447
rect 12267 3383 12776 3399
rect 13683 3403 14196 3417
rect 9680 3307 10151 3311
rect 9631 3292 10151 3307
rect 9631 2589 9692 3292
rect 11333 2589 11399 3342
rect 9434 2577 10352 2589
rect 9434 2560 9458 2577
rect 9642 2560 9687 2577
rect 9871 2560 9916 2577
rect 10100 2560 10145 2577
rect 10329 2560 10352 2577
rect 9434 2551 10352 2560
rect 10681 2580 11608 2589
rect 10681 2563 10711 2580
rect 10895 2563 10940 2580
rect 11124 2563 11169 2580
rect 11353 2563 11398 2580
rect 11582 2563 11608 2580
rect 9631 2485 9692 2551
rect 10681 2545 11608 2563
rect 9631 2457 9691 2485
rect 6029 2439 7028 2455
rect 6029 2390 7031 2439
rect 8822 2434 9691 2457
rect 8822 2415 9238 2434
rect 6479 2318 6588 2390
rect 6479 2249 6498 2318
rect 6567 2249 6588 2318
rect 6479 2065 6588 2249
rect 5427 2045 6030 2048
rect 5427 2016 5435 2045
rect 5778 2039 6030 2045
rect 6479 2047 6492 2065
rect 6562 2047 6588 2065
rect 6479 2040 6588 2047
rect 9227 2386 9238 2415
rect 9275 2415 9691 2434
rect 11333 2455 11399 2545
rect 12267 2455 12332 3383
rect 13683 3360 13699 3403
rect 13719 3360 14157 3403
rect 14177 3360 14196 3403
rect 16148 3392 16666 3403
rect 16148 3389 16631 3392
rect 14940 3380 15455 3382
rect 13683 3351 14196 3360
rect 14935 3364 15455 3380
rect 14935 3360 15411 3364
rect 14128 2457 14194 3351
rect 14935 3307 14950 3360
rect 14984 3311 15411 3360
rect 15445 3311 15455 3364
rect 16148 3353 16176 3389
rect 16193 3353 16631 3389
rect 16649 3353 16666 3392
rect 16148 3342 16666 3353
rect 17531 3402 17551 3443
rect 17569 3440 18040 3443
rect 17569 3402 18015 3440
rect 17531 3399 18015 3402
rect 18033 3399 18040 3440
rect 22836 3443 23345 3447
rect 17531 3383 18040 3399
rect 18947 3403 19460 3417
rect 14984 3307 15455 3311
rect 14935 3292 15455 3307
rect 14935 2589 14996 3292
rect 16597 2589 16663 3342
rect 14738 2577 15656 2589
rect 14738 2560 14762 2577
rect 14946 2560 14991 2577
rect 15175 2560 15220 2577
rect 15404 2560 15449 2577
rect 15633 2560 15656 2577
rect 14738 2551 15656 2560
rect 15945 2580 16872 2589
rect 15945 2563 15975 2580
rect 16159 2563 16204 2580
rect 16388 2563 16433 2580
rect 16617 2563 16662 2580
rect 16846 2563 16872 2580
rect 14935 2485 14996 2551
rect 15945 2545 16872 2563
rect 14935 2457 14995 2485
rect 11333 2439 12332 2455
rect 14126 2444 14995 2457
rect 9275 2386 9284 2415
rect 11333 2390 12335 2439
rect 14126 2415 14542 2444
rect 14531 2411 14542 2415
rect 14575 2415 14995 2444
rect 16597 2455 16663 2545
rect 17531 2455 17596 3383
rect 18947 3360 18963 3403
rect 18983 3360 19421 3403
rect 19441 3360 19460 3403
rect 21453 3392 21971 3403
rect 21453 3389 21936 3392
rect 20204 3380 20719 3382
rect 18947 3351 19460 3360
rect 20199 3364 20719 3380
rect 20199 3360 20675 3364
rect 19392 2457 19458 3351
rect 20199 3307 20214 3360
rect 20248 3311 20675 3360
rect 20709 3311 20719 3364
rect 21453 3353 21481 3389
rect 21498 3353 21936 3389
rect 21954 3353 21971 3392
rect 21453 3342 21971 3353
rect 22836 3402 22856 3443
rect 22874 3440 23345 3443
rect 22874 3402 23320 3440
rect 22836 3399 23320 3402
rect 23338 3399 23345 3440
rect 28100 3443 28609 3447
rect 22836 3383 23345 3399
rect 24252 3403 24765 3417
rect 20248 3307 20719 3311
rect 20199 3292 20719 3307
rect 20199 2589 20260 3292
rect 21902 2589 21968 3342
rect 20002 2577 20920 2589
rect 20002 2560 20026 2577
rect 20210 2560 20255 2577
rect 20439 2560 20484 2577
rect 20668 2560 20713 2577
rect 20897 2560 20920 2577
rect 20002 2551 20920 2560
rect 21250 2580 22177 2589
rect 21250 2563 21280 2580
rect 21464 2563 21509 2580
rect 21693 2563 21738 2580
rect 21922 2563 21967 2580
rect 22151 2563 22177 2580
rect 20199 2485 20260 2551
rect 21250 2545 22177 2563
rect 20199 2457 20259 2485
rect 16597 2439 17596 2455
rect 19390 2443 20259 2457
rect 14575 2411 14588 2415
rect 9227 2071 9284 2386
rect 9227 2051 9236 2071
rect 9278 2051 9284 2071
rect 11783 2354 11892 2390
rect 11783 2274 11805 2354
rect 11874 2274 11892 2354
rect 10814 2061 10936 2068
rect 11783 2065 11892 2274
rect 9227 2044 9284 2051
rect 9775 2044 9809 2054
rect 5778 2022 6004 2039
rect 6021 2022 6030 2039
rect 5778 2016 6030 2022
rect 5427 2013 6030 2016
rect 6477 2017 6599 2025
rect 6477 1994 6509 2017
rect 6562 1994 6599 2017
rect 6477 1963 6599 1994
rect 6477 1940 6505 1963
rect 6558 1940 6599 1963
rect 6477 1885 6599 1940
rect 9223 2023 9291 2028
rect 9223 2003 9236 2023
rect 9276 2003 9291 2023
rect 9223 1970 9291 2003
rect 9223 1950 9237 1970
rect 9277 1950 9291 1970
rect 9223 1885 9291 1950
rect 9775 2027 9784 2044
rect 9801 2027 9809 2044
rect 6477 1795 9298 1885
rect 9775 1873 9809 2027
rect 10814 2051 11160 2061
rect 10814 2004 10826 2051
rect 10920 2048 11160 2051
rect 10920 2039 11334 2048
rect 11783 2047 11796 2065
rect 11866 2047 11892 2065
rect 11783 2040 11892 2047
rect 14531 2071 14588 2411
rect 16597 2390 17599 2439
rect 19390 2415 19806 2443
rect 19795 2398 19806 2415
rect 19844 2415 20259 2443
rect 21902 2455 21968 2545
rect 22836 2455 22901 3383
rect 24252 3360 24268 3403
rect 24288 3360 24726 3403
rect 24746 3360 24765 3403
rect 26717 3392 27235 3403
rect 26717 3389 27200 3392
rect 25509 3380 26024 3382
rect 24252 3351 24765 3360
rect 25504 3364 26024 3380
rect 25504 3360 25980 3364
rect 24697 2457 24763 3351
rect 25504 3307 25519 3360
rect 25553 3311 25980 3360
rect 26014 3311 26024 3364
rect 26717 3353 26745 3389
rect 26762 3353 27200 3389
rect 27218 3353 27235 3392
rect 26717 3342 27235 3353
rect 28100 3402 28120 3443
rect 28138 3440 28609 3443
rect 28138 3402 28584 3440
rect 28100 3399 28584 3402
rect 28602 3399 28609 3440
rect 28100 3383 28609 3399
rect 29516 3403 30029 3417
rect 25553 3307 26024 3311
rect 25504 3292 26024 3307
rect 25504 2589 25565 3292
rect 27166 2589 27232 3342
rect 25307 2577 26225 2589
rect 25307 2560 25331 2577
rect 25515 2560 25560 2577
rect 25744 2560 25789 2577
rect 25973 2560 26018 2577
rect 26202 2560 26225 2577
rect 25307 2551 26225 2560
rect 26514 2580 27441 2589
rect 26514 2563 26544 2580
rect 26728 2563 26773 2580
rect 26957 2563 27002 2580
rect 27186 2563 27231 2580
rect 27415 2563 27441 2580
rect 25504 2485 25565 2551
rect 26514 2545 27441 2563
rect 25504 2457 25564 2485
rect 21902 2439 22901 2455
rect 24695 2449 25564 2457
rect 19844 2398 19852 2415
rect 14531 2051 14540 2071
rect 14582 2051 14588 2071
rect 17047 2347 17156 2390
rect 17047 2266 17059 2347
rect 17145 2266 17156 2347
rect 17047 2065 17156 2266
rect 16054 2056 16399 2061
rect 14531 2044 14588 2051
rect 15079 2044 15113 2054
rect 10920 2022 11308 2039
rect 11325 2022 11334 2039
rect 10920 2013 11334 2022
rect 11781 2017 11903 2025
rect 10920 2004 11160 2013
rect 10814 1992 11160 2004
rect 11781 1994 11813 2017
rect 11866 1994 11903 2017
rect 11781 1963 11903 1994
rect 11781 1940 11809 1963
rect 11862 1940 11903 1963
rect 11781 1885 11903 1940
rect 14527 2023 14595 2028
rect 14527 2003 14540 2023
rect 14580 2003 14595 2023
rect 14527 1970 14595 2003
rect 14527 1950 14541 1970
rect 14581 1950 14595 1970
rect 14527 1885 14595 1950
rect 15079 2027 15088 2044
rect 15105 2027 15113 2044
rect 15079 1897 15113 2027
rect 16054 1998 16058 2056
rect 16162 2048 16399 2056
rect 16162 2039 16598 2048
rect 17047 2047 17060 2065
rect 17130 2047 17156 2065
rect 17047 2040 17156 2047
rect 19795 2071 19852 2398
rect 21902 2390 22904 2439
rect 24695 2415 25106 2449
rect 25100 2413 25106 2415
rect 25150 2415 25564 2449
rect 27166 2455 27232 2545
rect 28100 2455 28165 3383
rect 29516 3360 29532 3403
rect 29552 3360 29990 3403
rect 30010 3360 30029 3403
rect 30773 3380 31288 3382
rect 29516 3351 30029 3360
rect 30768 3364 31288 3380
rect 30768 3360 31244 3364
rect 29961 2457 30027 3351
rect 30768 3307 30783 3360
rect 30817 3311 31244 3360
rect 31278 3311 31288 3364
rect 30817 3307 31288 3311
rect 30768 3292 31288 3307
rect 30768 2589 30829 3292
rect 30571 2577 31489 2589
rect 30571 2560 30595 2577
rect 30779 2560 30824 2577
rect 31008 2560 31053 2577
rect 31237 2560 31282 2577
rect 31466 2560 31489 2577
rect 30571 2551 31489 2560
rect 30768 2485 30829 2551
rect 30768 2457 30828 2485
rect 27166 2439 28165 2455
rect 29959 2448 30828 2457
rect 25150 2413 25157 2415
rect 22352 2370 22461 2390
rect 22352 2281 22373 2370
rect 22444 2281 22461 2370
rect 19795 2051 19804 2071
rect 19846 2051 19852 2071
rect 21391 2089 21692 2107
rect 19795 2044 19852 2051
rect 20343 2044 20377 2055
rect 16162 2022 16572 2039
rect 16589 2022 16598 2039
rect 16162 2013 16598 2022
rect 17045 2017 17167 2025
rect 16162 1998 16399 2013
rect 16054 1993 16399 1998
rect 17045 1994 17077 2017
rect 17130 1994 17167 2017
rect 17045 1963 17167 1994
rect 17045 1940 17073 1963
rect 17126 1940 17167 1963
rect 9751 1831 9838 1873
rect 6477 1792 6599 1795
rect 8111 1488 8257 1795
rect 9751 1791 9766 1831
rect 9818 1791 9838 1831
rect 11781 1795 14602 1885
rect 15002 1848 15192 1897
rect 11781 1792 11903 1795
rect 9751 1772 9838 1791
rect 13415 1488 13561 1795
rect 15002 1779 15066 1848
rect 15136 1779 15192 1848
rect 17045 1885 17167 1940
rect 19791 2023 19859 2028
rect 19791 2003 19804 2023
rect 19844 2003 19859 2023
rect 19791 1970 19859 2003
rect 19791 1950 19805 1970
rect 19845 1950 19859 1970
rect 19791 1885 19859 1950
rect 20343 2027 20352 2044
rect 20369 2027 20377 2044
rect 17045 1795 19866 1885
rect 20343 1875 20377 2027
rect 21391 1927 21403 2089
rect 21480 2048 21692 2089
rect 22352 2065 22461 2281
rect 21480 2039 21903 2048
rect 22352 2047 22365 2065
rect 22435 2047 22461 2065
rect 22352 2040 22461 2047
rect 25100 2071 25157 2413
rect 27166 2390 28168 2439
rect 29959 2415 30372 2448
rect 30364 2402 30372 2415
rect 30410 2415 30828 2448
rect 30410 2402 30421 2415
rect 27616 2306 27725 2390
rect 27616 2196 27623 2306
rect 27712 2196 27725 2306
rect 25100 2051 25109 2071
rect 25151 2051 25157 2071
rect 26634 2092 26922 2119
rect 25100 2044 25157 2051
rect 25648 2044 25682 2054
rect 21480 2022 21877 2039
rect 21894 2022 21903 2039
rect 21480 2013 21903 2022
rect 22350 2017 22472 2025
rect 21480 1927 21692 2013
rect 21391 1915 21692 1927
rect 22350 1994 22382 2017
rect 22435 1994 22472 2017
rect 22350 1963 22472 1994
rect 22350 1940 22378 1963
rect 22431 1940 22472 1963
rect 22350 1885 22472 1940
rect 25096 2023 25164 2028
rect 25096 2003 25109 2023
rect 25149 2003 25164 2023
rect 25096 1970 25164 2003
rect 25096 1950 25110 1970
rect 25150 1950 25164 1970
rect 25096 1885 25164 1950
rect 25648 2027 25657 2044
rect 25674 2027 25682 2044
rect 25648 1891 25682 2027
rect 26634 1955 26659 2092
rect 26890 2048 26922 2092
rect 27616 2065 27725 2196
rect 26890 2039 27167 2048
rect 27616 2047 27629 2065
rect 27699 2047 27725 2065
rect 27616 2040 27725 2047
rect 30364 2071 30421 2402
rect 30364 2051 30373 2071
rect 30415 2051 30421 2071
rect 30364 2044 30421 2051
rect 30912 2044 30947 2054
rect 26890 2022 27141 2039
rect 27158 2022 27167 2039
rect 26890 2013 27167 2022
rect 27614 2017 27736 2025
rect 26890 1955 26922 2013
rect 26634 1930 26922 1955
rect 27614 1994 27646 2017
rect 27699 1994 27736 2017
rect 27614 1963 27736 1994
rect 27614 1940 27642 1963
rect 27695 1940 27736 1963
rect 20282 1821 20478 1875
rect 17045 1792 17167 1795
rect 15002 1727 15192 1779
rect 15079 1726 15113 1727
rect 18679 1488 18825 1795
rect 20282 1739 20336 1821
rect 20419 1739 20478 1821
rect 22350 1795 25171 1885
rect 25589 1861 25752 1891
rect 22350 1792 22472 1795
rect 20282 1684 20478 1739
rect 23984 1488 24130 1795
rect 25589 1730 25606 1861
rect 25734 1730 25752 1861
rect 27614 1885 27736 1940
rect 30360 2023 30428 2028
rect 30360 2003 30373 2023
rect 30413 2003 30428 2023
rect 30360 1970 30428 2003
rect 30360 1950 30374 1970
rect 30414 1950 30428 1970
rect 30360 1885 30428 1950
rect 30912 2027 30921 2044
rect 30938 2027 30947 2044
rect 30912 1895 30947 2027
rect 27614 1795 30435 1885
rect 30865 1876 31002 1895
rect 27614 1792 27736 1795
rect 25589 1713 25752 1730
rect 29248 1488 29394 1795
rect 30865 1793 30893 1876
rect 30980 1793 31002 1876
rect 30865 1649 31002 1793
rect 7183 1485 9537 1488
rect 7183 1481 8582 1485
rect 7183 1479 8128 1481
rect 7183 1431 7211 1479
rect 7235 1475 8128 1479
rect 7235 1431 7669 1475
rect 7183 1427 7669 1431
rect 7693 1433 8128 1475
rect 8152 1437 8582 1481
rect 8606 1482 9537 1485
rect 8606 1437 9035 1482
rect 8152 1434 9035 1437
rect 9059 1434 9501 1482
rect 9525 1434 9537 1482
rect 8152 1433 9537 1434
rect 7693 1427 9537 1433
rect 7183 1422 9537 1427
rect 12487 1485 14841 1488
rect 12487 1481 13886 1485
rect 12487 1479 13432 1481
rect 12487 1431 12515 1479
rect 12539 1475 13432 1479
rect 12539 1431 12973 1475
rect 12487 1427 12973 1431
rect 12997 1433 13432 1475
rect 13456 1437 13886 1481
rect 13910 1482 14841 1485
rect 13910 1437 14339 1482
rect 13456 1434 14339 1437
rect 14363 1434 14805 1482
rect 14829 1434 14841 1482
rect 13456 1433 14841 1434
rect 12997 1427 14841 1433
rect 12487 1422 14841 1427
rect 17751 1485 20105 1488
rect 17751 1481 19150 1485
rect 17751 1479 18696 1481
rect 17751 1431 17779 1479
rect 17803 1475 18696 1479
rect 17803 1431 18237 1475
rect 17751 1427 18237 1431
rect 18261 1433 18696 1475
rect 18720 1437 19150 1481
rect 19174 1482 20105 1485
rect 19174 1437 19603 1482
rect 18720 1434 19603 1437
rect 19627 1434 20069 1482
rect 20093 1434 20105 1482
rect 18720 1433 20105 1434
rect 18261 1427 20105 1433
rect 17751 1422 20105 1427
rect 23056 1485 25410 1488
rect 23056 1481 24455 1485
rect 23056 1479 24001 1481
rect 23056 1431 23084 1479
rect 23108 1475 24001 1479
rect 23108 1431 23542 1475
rect 23056 1427 23542 1431
rect 23566 1433 24001 1475
rect 24025 1437 24455 1481
rect 24479 1482 25410 1485
rect 24479 1437 24908 1482
rect 24025 1434 24908 1437
rect 24932 1434 25374 1482
rect 25398 1434 25410 1482
rect 24025 1433 25410 1434
rect 23566 1427 25410 1433
rect 23056 1422 25410 1427
rect 28320 1485 30674 1488
rect 28320 1481 29719 1485
rect 28320 1479 29265 1481
rect 28320 1431 28348 1479
rect 28372 1475 29265 1479
rect 28372 1431 28806 1475
rect 28320 1427 28806 1431
rect 28830 1433 29265 1475
rect 29289 1437 29719 1481
rect 29743 1482 30674 1485
rect 29743 1437 30172 1482
rect 29289 1434 30172 1437
rect 30196 1434 30638 1482
rect 30662 1434 30674 1482
rect 29289 1433 30674 1434
rect 28830 1427 30674 1433
rect 28320 1422 30674 1427
rect 8111 1417 8257 1422
rect 13415 1417 13561 1422
rect 18679 1417 18825 1422
rect 23984 1417 24130 1422
rect 29248 1417 29394 1422
rect 7401 1393 9778 1396
rect 7401 1390 9720 1393
rect 7401 1384 8348 1390
rect 7401 1378 7889 1384
rect 7401 1323 7427 1378
rect 7462 1329 7889 1378
rect 7924 1379 8348 1384
rect 8383 1379 8810 1390
rect 7924 1329 8342 1379
rect 8399 1335 8810 1379
rect 8845 1384 9720 1390
rect 8845 1335 9272 1384
rect 7462 1325 8342 1329
rect 8399 1329 9272 1335
rect 9307 1338 9720 1384
rect 9755 1338 9778 1393
rect 9307 1329 9778 1338
rect 8399 1325 9778 1329
rect 7462 1323 9778 1325
rect 7401 1314 9778 1323
rect 12705 1393 15082 1396
rect 12705 1390 15024 1393
rect 12705 1384 13652 1390
rect 12705 1378 13193 1384
rect 12705 1323 12731 1378
rect 12766 1329 13193 1378
rect 13228 1379 13652 1384
rect 13687 1379 14114 1390
rect 13228 1329 13646 1379
rect 13703 1335 14114 1379
rect 14149 1384 15024 1390
rect 14149 1335 14576 1384
rect 12766 1325 13646 1329
rect 13703 1329 14576 1335
rect 14611 1338 15024 1384
rect 15059 1338 15082 1393
rect 14611 1329 15082 1338
rect 13703 1325 15082 1329
rect 12766 1323 15082 1325
rect 12705 1314 15082 1323
rect 17969 1393 20346 1396
rect 17969 1390 20288 1393
rect 17969 1384 18916 1390
rect 17969 1378 18457 1384
rect 17969 1323 17995 1378
rect 18030 1329 18457 1378
rect 18492 1379 18916 1384
rect 18951 1379 19378 1390
rect 18492 1329 18910 1379
rect 18967 1335 19378 1379
rect 19413 1384 20288 1390
rect 19413 1335 19840 1384
rect 18030 1325 18910 1329
rect 18967 1329 19840 1335
rect 19875 1338 20288 1384
rect 20323 1338 20346 1393
rect 19875 1329 20346 1338
rect 18967 1325 20346 1329
rect 18030 1323 20346 1325
rect 17969 1314 20346 1323
rect 23274 1393 25651 1396
rect 23274 1390 25593 1393
rect 23274 1384 24221 1390
rect 23274 1378 23762 1384
rect 23274 1323 23300 1378
rect 23335 1329 23762 1378
rect 23797 1379 24221 1384
rect 24256 1379 24683 1390
rect 23797 1329 24215 1379
rect 24272 1335 24683 1379
rect 24718 1384 25593 1390
rect 24718 1335 25145 1384
rect 23335 1325 24215 1329
rect 24272 1329 25145 1335
rect 25180 1338 25593 1384
rect 25628 1338 25651 1393
rect 25180 1329 25651 1338
rect 24272 1325 25651 1329
rect 23335 1323 25651 1325
rect 23274 1314 25651 1323
rect 28538 1393 30915 1396
rect 28538 1390 30857 1393
rect 28538 1384 29485 1390
rect 28538 1378 29026 1384
rect 28538 1323 28564 1378
rect 28599 1329 29026 1378
rect 29061 1379 29485 1384
rect 29520 1379 29947 1390
rect 29061 1329 29479 1379
rect 29536 1335 29947 1379
rect 29982 1384 30857 1390
rect 29982 1335 30409 1384
rect 28599 1325 29479 1329
rect 29536 1329 30409 1335
rect 30444 1338 30857 1384
rect 30892 1338 30915 1393
rect 30444 1329 30915 1338
rect 29536 1325 30915 1329
rect 28599 1323 30915 1325
rect 28538 1314 30915 1323
rect 6433 307 30901 324
rect 6433 290 7245 307
rect 7429 290 7474 307
rect 7658 290 7703 307
rect 7887 290 7932 307
rect 8116 290 8161 307
rect 8345 290 8390 307
rect 8574 290 8619 307
rect 8803 290 8848 307
rect 9032 290 9077 307
rect 9261 290 9306 307
rect 9490 290 9535 307
rect 9719 290 12549 307
rect 12733 290 12778 307
rect 12962 290 13007 307
rect 13191 290 13236 307
rect 13420 290 13465 307
rect 13649 290 13694 307
rect 13878 290 13923 307
rect 14107 290 14152 307
rect 14336 290 14381 307
rect 14565 290 14610 307
rect 14794 290 14839 307
rect 15023 290 17813 307
rect 17997 290 18042 307
rect 18226 290 18271 307
rect 18455 290 18500 307
rect 18684 290 18729 307
rect 18913 290 18958 307
rect 19142 290 19187 307
rect 19371 290 19416 307
rect 19600 290 19645 307
rect 19829 290 19874 307
rect 20058 290 20103 307
rect 20287 290 23118 307
rect 23302 290 23347 307
rect 23531 290 23576 307
rect 23760 290 23805 307
rect 23989 290 24034 307
rect 24218 290 24263 307
rect 24447 290 24492 307
rect 24676 290 24721 307
rect 24905 290 24950 307
rect 25134 290 25179 307
rect 25363 290 25408 307
rect 25592 290 28382 307
rect 28566 290 28611 307
rect 28795 290 28840 307
rect 29024 290 29069 307
rect 29253 290 29298 307
rect 29482 290 29527 307
rect 29711 290 29756 307
rect 29940 290 29985 307
rect 30169 290 30214 307
rect 30398 290 30443 307
rect 30627 290 30672 307
rect 30856 290 30901 307
rect 6433 283 30901 290
rect 6433 281 7273 283
rect 12296 281 12577 283
rect 17560 281 17841 283
rect 22865 281 23146 283
rect 28129 281 28410 283
rect 9161 252 9249 266
rect 9161 235 9172 252
rect 9223 235 9249 252
rect 9161 181 9249 235
rect 14465 252 14553 266
rect 14465 235 14476 252
rect 14527 235 14553 252
rect 14465 181 14553 235
rect 19729 252 19817 266
rect 19729 235 19740 252
rect 19791 235 19817 252
rect 19729 181 19817 235
rect 25034 252 25122 266
rect 25034 235 25045 252
rect 25096 235 25122 252
rect 25034 181 25122 235
rect 30298 252 30386 266
rect 30298 235 30309 252
rect 30360 235 30386 252
rect 30298 181 30386 235
rect 5274 139 31632 181
rect 5274 136 8574 139
rect 5274 82 7186 136
rect 7243 128 8104 136
rect 7243 82 7659 128
rect 5274 74 7659 82
rect 7716 82 8104 128
rect 8161 127 8574 136
rect 8161 82 8342 127
rect 7716 74 8342 82
rect 5274 73 8342 74
rect 8399 85 8574 127
rect 8631 136 9485 139
rect 8631 85 9038 136
rect 8399 82 9038 85
rect 9095 85 9485 136
rect 9542 136 13878 139
rect 9542 85 12490 136
rect 9095 82 12490 85
rect 12547 128 13408 136
rect 12547 82 12963 128
rect 8399 74 12963 82
rect 13020 82 13408 128
rect 13465 127 13878 136
rect 13465 82 13646 127
rect 13020 74 13646 82
rect 8399 73 13646 74
rect 13703 85 13878 127
rect 13935 136 14789 139
rect 13935 85 14342 136
rect 13703 82 14342 85
rect 14399 85 14789 136
rect 14846 136 19142 139
rect 14846 85 17754 136
rect 14399 82 17754 85
rect 17811 128 18672 136
rect 17811 82 18227 128
rect 13703 74 18227 82
rect 18284 82 18672 128
rect 18729 127 19142 136
rect 18729 82 18910 127
rect 18284 74 18910 82
rect 13703 73 18910 74
rect 18967 85 19142 127
rect 19199 136 20053 139
rect 19199 85 19606 136
rect 18967 82 19606 85
rect 19663 85 20053 136
rect 20110 136 24447 139
rect 20110 85 23059 136
rect 19663 82 23059 85
rect 23116 128 23977 136
rect 23116 82 23532 128
rect 18967 74 23532 82
rect 23589 82 23977 128
rect 24034 127 24447 136
rect 24034 82 24215 127
rect 23589 74 24215 82
rect 18967 73 24215 74
rect 24272 85 24447 127
rect 24504 136 25358 139
rect 24504 85 24911 136
rect 24272 82 24911 85
rect 24968 85 25358 136
rect 25415 136 29711 139
rect 25415 85 28323 136
rect 24968 82 28323 85
rect 28380 128 29241 136
rect 28380 82 28796 128
rect 24272 74 28796 82
rect 28853 82 29241 128
rect 29298 127 29711 136
rect 29298 82 29479 127
rect 28853 74 29479 82
rect 24272 73 29479 74
rect 29536 85 29711 127
rect 29768 136 30622 139
rect 29768 85 30175 136
rect 29536 82 30175 85
rect 30232 85 30622 136
rect 30679 85 31632 139
rect 30232 82 31632 85
rect 29536 73 31632 82
rect 5274 -64 31632 73
<< via1 >>
rect 8160 3843 8187 3848
rect 6748 3790 6804 3835
rect 8160 3803 8187 3843
rect 13464 3843 13491 3848
rect 12052 3790 12108 3835
rect 13464 3803 13491 3843
rect 18728 3843 18755 3848
rect 17316 3790 17372 3835
rect 18728 3803 18755 3843
rect 24033 3843 24060 3848
rect 22621 3790 22677 3835
rect 24033 3803 24060 3843
rect 29297 3843 29324 3848
rect 27885 3790 27941 3835
rect 29297 3803 29324 3843
rect 7882 3592 7986 3652
rect 6750 3511 6754 3547
rect 6754 3511 6772 3547
rect 6772 3511 6803 3547
rect 6750 3501 6803 3511
rect 8159 3503 8164 3544
rect 8164 3503 8186 3544
rect 8159 3499 8186 3503
rect 13187 3590 13291 3649
rect 12054 3511 12058 3547
rect 12058 3511 12076 3547
rect 12076 3511 12107 3547
rect 12054 3501 12107 3511
rect 13463 3503 13468 3544
rect 13468 3503 13490 3544
rect 13463 3499 13490 3503
rect 18452 3590 18555 3649
rect 17318 3511 17322 3547
rect 17322 3511 17340 3547
rect 17340 3511 17371 3547
rect 17318 3501 17371 3511
rect 18727 3503 18732 3544
rect 18732 3503 18754 3544
rect 18727 3499 18754 3503
rect 23743 3590 23847 3649
rect 22623 3511 22627 3547
rect 22627 3511 22645 3547
rect 22645 3511 22676 3547
rect 22623 3501 22676 3511
rect 24032 3503 24037 3544
rect 24037 3503 24059 3544
rect 24032 3499 24059 3503
rect 29028 3597 29132 3656
rect 27887 3511 27891 3547
rect 27891 3511 27909 3547
rect 27909 3511 27940 3547
rect 27887 3501 27940 3511
rect 29296 3503 29301 3544
rect 29301 3503 29323 3544
rect 29296 3499 29323 3503
rect 6498 2249 6567 2318
rect 5435 2016 5778 2045
rect 9238 2386 9275 2434
rect 14542 2411 14575 2444
rect 11805 2274 11874 2354
rect 10826 2004 10920 2051
rect 19806 2398 19844 2443
rect 17059 2266 17145 2347
rect 16058 1998 16162 2056
rect 25106 2413 25150 2449
rect 22373 2281 22444 2370
rect 9766 1791 9818 1831
rect 15066 1779 15136 1848
rect 21403 1927 21480 2089
rect 30372 2402 30410 2448
rect 27623 2196 27712 2306
rect 26659 1955 26890 2092
rect 20336 1739 20419 1821
rect 25606 1730 25734 1861
rect 30893 1793 30980 1876
rect 8342 1335 8348 1379
rect 8348 1335 8383 1379
rect 8383 1335 8399 1379
rect 8342 1325 8399 1335
rect 13646 1335 13652 1379
rect 13652 1335 13687 1379
rect 13687 1335 13703 1379
rect 13646 1325 13703 1335
rect 18910 1335 18916 1379
rect 18916 1335 18951 1379
rect 18951 1335 18967 1379
rect 18910 1325 18967 1335
rect 24215 1335 24221 1379
rect 24221 1335 24256 1379
rect 24256 1335 24272 1379
rect 24215 1325 24272 1335
rect 29479 1335 29485 1379
rect 29485 1335 29520 1379
rect 29520 1335 29536 1379
rect 29479 1325 29536 1335
rect 8342 73 8399 127
rect 13646 73 13703 127
rect 18910 73 18967 127
rect 24215 73 24272 127
rect 29479 73 29536 127
<< metal2 >>
rect 2420 7135 5195 7136
rect 32007 7135 32932 7153
rect 2420 7062 32932 7135
rect 2420 6541 32338 7062
rect 32847 6541 32932 7062
rect 2420 6474 32932 6541
rect 2420 6471 32160 6474
rect 2420 1847 3283 6471
rect 5084 5574 32135 5577
rect 4369 4913 32135 5574
rect 4369 2141 5139 4913
rect 6737 3835 6823 3882
rect 6737 3790 6748 3835
rect 6804 3790 6823 3835
rect 6737 3547 6823 3790
rect 8152 3848 8195 3886
rect 8152 3803 8160 3848
rect 8187 3803 8195 3848
rect 7861 3666 8005 3675
rect 7861 3580 7870 3666
rect 7997 3580 8005 3666
rect 7861 3571 8005 3580
rect 6737 3501 6750 3547
rect 6803 3501 6823 3547
rect 6737 3481 6823 3501
rect 8152 3544 8195 3803
rect 8152 3499 8159 3544
rect 8186 3499 8195 3544
rect 8152 3483 8195 3499
rect 12041 3835 12127 3882
rect 12041 3790 12052 3835
rect 12108 3790 12127 3835
rect 12041 3547 12127 3790
rect 13456 3848 13499 3886
rect 13456 3803 13464 3848
rect 13491 3803 13499 3848
rect 13166 3663 13310 3673
rect 13166 3578 13175 3663
rect 13302 3578 13310 3663
rect 13166 3568 13310 3578
rect 12041 3501 12054 3547
rect 12107 3501 12127 3547
rect 12041 3481 12127 3501
rect 13456 3544 13499 3803
rect 13456 3499 13463 3544
rect 13490 3499 13499 3544
rect 13456 3483 13499 3499
rect 17305 3835 17391 3882
rect 17305 3790 17316 3835
rect 17372 3790 17391 3835
rect 17305 3547 17391 3790
rect 18720 3848 18763 3886
rect 18720 3803 18728 3848
rect 18755 3803 18763 3848
rect 18430 3663 18575 3673
rect 18430 3578 18440 3663
rect 18566 3578 18575 3663
rect 18430 3568 18575 3578
rect 17305 3501 17318 3547
rect 17371 3501 17391 3547
rect 17305 3481 17391 3501
rect 18720 3544 18763 3803
rect 18720 3499 18727 3544
rect 18754 3499 18763 3544
rect 18720 3483 18763 3499
rect 22610 3835 22696 3882
rect 22610 3790 22621 3835
rect 22677 3790 22696 3835
rect 22610 3547 22696 3790
rect 24025 3848 24068 3886
rect 24025 3803 24033 3848
rect 24060 3803 24068 3848
rect 23722 3663 23866 3673
rect 23722 3578 23731 3663
rect 23858 3578 23866 3663
rect 23722 3568 23866 3578
rect 22610 3501 22623 3547
rect 22676 3501 22696 3547
rect 22610 3481 22696 3501
rect 24025 3544 24068 3803
rect 24025 3499 24032 3544
rect 24059 3499 24068 3544
rect 24025 3483 24068 3499
rect 27874 3835 27960 3882
rect 27874 3790 27885 3835
rect 27941 3790 27960 3835
rect 27874 3547 27960 3790
rect 29289 3848 29332 3886
rect 29289 3803 29297 3848
rect 29324 3803 29332 3848
rect 29007 3670 29151 3680
rect 29007 3585 29016 3670
rect 29143 3585 29151 3670
rect 29007 3575 29151 3585
rect 27874 3501 27887 3547
rect 27940 3501 27960 3547
rect 27874 3481 27960 3501
rect 29289 3544 29332 3803
rect 29289 3499 29296 3544
rect 29323 3499 29332 3544
rect 29289 3483 29332 3499
rect 14529 2455 14591 2462
rect 9225 2442 9286 2455
rect 9225 2384 9234 2442
rect 9277 2384 9286 2442
rect 14529 2406 14538 2455
rect 14583 2406 14591 2455
rect 14529 2398 14591 2406
rect 19785 2449 19862 2460
rect 19785 2401 19797 2449
rect 19850 2401 19862 2449
rect 25099 2454 25160 2460
rect 25099 2412 25105 2454
rect 25153 2412 25160 2454
rect 25099 2406 25160 2412
rect 30358 2450 30432 2465
rect 19785 2398 19806 2401
rect 19844 2398 19862 2401
rect 19785 2388 19862 2398
rect 30358 2398 30369 2450
rect 30424 2398 30432 2450
rect 30358 2387 30432 2398
rect 9225 2375 9286 2384
rect 22334 2370 26782 2386
rect 16021 2362 16183 2365
rect 11763 2354 16183 2362
rect 6456 2318 10937 2331
rect 6456 2249 6498 2318
rect 6567 2249 10937 2318
rect 11763 2274 11805 2354
rect 11874 2274 16183 2354
rect 11763 2252 16183 2274
rect 6456 2225 10937 2249
rect 4369 2097 5510 2141
rect 4369 2045 6032 2097
rect 4369 2016 5435 2045
rect 5778 2016 6032 2045
rect 4369 1965 6032 2016
rect 10814 2051 10937 2225
rect 10814 2004 10826 2051
rect 10920 2004 10937 2051
rect 10814 1992 10937 2004
rect 16021 2056 16183 2252
rect 17033 2347 21498 2362
rect 17033 2266 17059 2347
rect 17145 2266 21498 2347
rect 17033 2250 21498 2266
rect 22334 2281 22373 2370
rect 22444 2281 26782 2370
rect 31843 2337 32135 4913
rect 22334 2255 26782 2281
rect 27585 2306 32135 2337
rect 16021 1998 16058 2056
rect 16162 1998 16183 2056
rect 4369 1962 5510 1965
rect 16021 1902 16183 1998
rect 21390 2089 21496 2250
rect 21390 1927 21403 2089
rect 21480 1927 21496 2089
rect 26634 2119 26780 2255
rect 27585 2196 27623 2306
rect 27712 2196 32135 2306
rect 27585 2151 32135 2196
rect 31843 2149 32135 2151
rect 26634 2092 26922 2119
rect 26634 1955 26659 2092
rect 26890 1955 26922 2092
rect 26634 1930 26922 1955
rect 21390 1917 21496 1927
rect 15002 1848 15192 1897
rect 2420 1844 4480 1847
rect 2420 1831 9838 1844
rect 2420 1791 9766 1831
rect 9818 1791 9838 1831
rect 2420 1713 9838 1791
rect 15002 1840 15066 1848
rect 15136 1840 15192 1848
rect 15002 1735 15012 1840
rect 15180 1735 15192 1840
rect 15002 1727 15192 1735
rect 20282 1821 20478 1875
rect 20282 1753 20336 1821
rect 20419 1753 20478 1821
rect 2420 1616 4480 1713
rect 20282 1698 20300 1753
rect 20457 1698 20478 1753
rect 25589 1861 25752 1891
rect 25589 1730 25606 1861
rect 25734 1822 25752 1861
rect 25737 1739 25752 1822
rect 25734 1730 25752 1739
rect 25589 1713 25752 1730
rect 30865 1876 31002 1895
rect 30865 1793 30893 1876
rect 30980 1793 31002 1876
rect 30865 1757 31002 1793
rect 20282 1684 20478 1698
rect 30865 1655 30874 1757
rect 30957 1655 31002 1757
rect 30865 1649 31002 1655
rect 2420 1604 3283 1616
rect 8331 1379 8422 1390
rect 8331 1325 8342 1379
rect 8399 1325 8422 1379
rect 8331 127 8422 1325
rect 8331 73 8342 127
rect 8399 73 8422 127
rect 8331 69 8422 73
rect 13635 1379 13726 1390
rect 13635 1325 13646 1379
rect 13703 1325 13726 1379
rect 13635 127 13726 1325
rect 13635 73 13646 127
rect 13703 73 13726 127
rect 13635 69 13726 73
rect 18899 1379 18990 1390
rect 18899 1325 18910 1379
rect 18967 1325 18990 1379
rect 18899 127 18990 1325
rect 18899 73 18910 127
rect 18967 73 18990 127
rect 18899 69 18990 73
rect 24204 1379 24295 1390
rect 24204 1325 24215 1379
rect 24272 1325 24295 1379
rect 24204 127 24295 1325
rect 24204 73 24215 127
rect 24272 73 24295 127
rect 24204 69 24295 73
rect 29468 1379 29559 1390
rect 29468 1325 29479 1379
rect 29536 1325 29559 1379
rect 29468 127 29559 1325
rect 29468 73 29479 127
rect 29536 73 29559 127
rect 29468 69 29559 73
<< via2 >>
rect 32338 6541 32847 7062
rect 7870 3652 7997 3666
rect 7870 3592 7882 3652
rect 7882 3592 7986 3652
rect 7986 3592 7997 3652
rect 7870 3580 7997 3592
rect 13175 3649 13302 3663
rect 13175 3590 13187 3649
rect 13187 3590 13291 3649
rect 13291 3590 13302 3649
rect 13175 3578 13302 3590
rect 18440 3649 18566 3663
rect 18440 3590 18452 3649
rect 18452 3590 18555 3649
rect 18555 3590 18566 3649
rect 18440 3578 18566 3590
rect 23731 3649 23858 3663
rect 23731 3590 23743 3649
rect 23743 3590 23847 3649
rect 23847 3590 23858 3649
rect 23731 3578 23858 3590
rect 29016 3656 29143 3670
rect 29016 3597 29028 3656
rect 29028 3597 29132 3656
rect 29132 3597 29143 3656
rect 29016 3585 29143 3597
rect 9234 2434 9277 2442
rect 9234 2386 9238 2434
rect 9238 2386 9275 2434
rect 9275 2386 9277 2434
rect 9234 2384 9277 2386
rect 14538 2444 14583 2455
rect 14538 2411 14542 2444
rect 14542 2411 14575 2444
rect 14575 2411 14583 2444
rect 14538 2406 14583 2411
rect 19797 2443 19850 2449
rect 19797 2401 19806 2443
rect 19806 2401 19844 2443
rect 19844 2401 19850 2443
rect 25105 2449 25153 2454
rect 25105 2413 25106 2449
rect 25106 2413 25150 2449
rect 25150 2413 25153 2449
rect 25105 2412 25153 2413
rect 30369 2448 30424 2450
rect 30369 2402 30372 2448
rect 30372 2402 30410 2448
rect 30410 2402 30424 2448
rect 30369 2398 30424 2402
rect 15012 1779 15066 1840
rect 15066 1779 15136 1840
rect 15136 1779 15180 1840
rect 15012 1735 15180 1779
rect 20300 1739 20336 1753
rect 20336 1739 20419 1753
rect 20419 1739 20457 1753
rect 20300 1698 20457 1739
rect 25608 1739 25734 1822
rect 25734 1739 25737 1822
rect 30874 1655 30957 1757
<< metal3 >>
rect 32281 7062 32939 7157
rect 32281 6541 32338 7062
rect 32847 6541 32939 7062
rect 7611 4343 29158 4375
rect 7611 4182 7641 4343
rect 7877 4182 29158 4343
rect 7611 4153 29158 4182
rect 7855 3666 8012 4153
rect 7855 3580 7870 3666
rect 7997 3580 8012 3666
rect 7855 3563 8012 3580
rect 13160 3663 13317 4153
rect 13160 3578 13175 3663
rect 13302 3578 13317 3663
rect 13160 3561 13317 3578
rect 18424 3681 18581 4153
rect 18424 3663 18582 3681
rect 18424 3578 18440 3663
rect 18566 3578 18582 3663
rect 18424 3561 18582 3578
rect 23716 3663 23873 4153
rect 23716 3578 23731 3663
rect 23858 3578 23873 3663
rect 23716 3561 23873 3578
rect 29001 3670 29158 4153
rect 29001 3585 29016 3670
rect 29143 3585 29158 3670
rect 29001 3568 29158 3585
rect 32281 2471 32939 6541
rect 9220 2442 10463 2458
rect 9220 2384 9234 2442
rect 9277 2384 10463 2442
rect 14503 2455 15839 2468
rect 14503 2406 14538 2455
rect 14583 2406 15839 2455
rect 14503 2388 15839 2406
rect 19766 2449 21167 2468
rect 19766 2401 19797 2449
rect 19850 2401 21167 2449
rect 9220 2373 10463 2384
rect 10377 2075 10463 2373
rect 10354 1854 10504 2075
rect 10354 1840 15192 1854
rect 10354 1735 15012 1840
rect 15180 1735 15192 1840
rect 10354 1727 15192 1735
rect 15684 1772 15838 2388
rect 19766 2380 21167 2401
rect 25093 2454 26528 2469
rect 25093 2412 25105 2454
rect 25153 2412 26528 2454
rect 25093 2400 26528 2412
rect 30346 2450 32939 2471
rect 21030 1837 21166 2380
rect 21030 1822 25745 1837
rect 15684 1753 20475 1772
rect 10354 1724 10504 1727
rect 15684 1698 20300 1753
rect 20457 1698 20475 1753
rect 15684 1684 20475 1698
rect 21030 1739 25608 1822
rect 25737 1739 25745 1822
rect 26414 1770 26527 2400
rect 30346 2398 30369 2450
rect 30424 2398 32939 2450
rect 30346 2378 32939 2398
rect 32281 2343 32939 2378
rect 21030 1718 25745 1739
rect 26410 1757 30965 1770
rect 21030 1571 21166 1718
rect 26410 1655 30874 1757
rect 30957 1655 30965 1757
rect 26410 1646 30965 1655
rect 26414 1535 26527 1646
<< via3 >>
rect 7641 4182 7877 4343
<< metal4 >>
rect 7609 4355 7926 4386
rect 7609 4343 7646 4355
rect 7609 4182 7641 4343
rect 7609 4175 7646 4182
rect 7901 4175 7926 4355
rect 7609 4145 7926 4175
<< via4 >>
rect 7646 4343 7901 4355
rect 7646 4182 7877 4343
rect 7877 4182 7901 4343
rect 7646 4175 7901 4182
<< metal5 >>
rect 7519 4355 7967 4450
rect 7519 4175 7646 4355
rect 7901 4175 7967 4355
rect 7519 4119 7967 4175
<< labels >>
rlabel metal1 5887 3761 5997 3875 1 Vdd
port 1 n
rlabel metal1 7925 3619 7990 3644 1 Vctrl
port 3 n
rlabel metal1 7001 287 7047 322 1 vbn
port 8 n
rlabel metal1 8229 65 8308 123 1 Gnd
port 9 n
rlabel metal1 16455 3761 16565 3875 1 Vdd
port 1 n
rlabel metal1 18493 3619 18558 3644 1 Vctrl
port 3 n
rlabel metal1 17569 287 17615 322 1 vbn
port 8 n
rlabel metal1 18797 65 18876 123 1 Gnd
port 9 n
rlabel metal1 11191 3761 11301 3875 1 Vdd
port 1 n
rlabel metal1 13229 3619 13294 3644 1 Vctrl
port 3 n
rlabel metal1 12305 287 12351 322 1 vbn
port 8 n
rlabel metal1 13533 65 13612 123 1 Gnd
port 9 n
rlabel metal1 27024 3761 27134 3875 1 Vdd
port 1 n
rlabel via1 29062 3619 29127 3644 1 Vctrl
port 3 n
rlabel metal1 28138 287 28184 322 1 vbn
port 8 n
rlabel metal1 29366 65 29445 123 1 Gnd
port 9 n
rlabel metal1 21760 3761 21870 3875 1 Vdd
port 1 n
rlabel metal1 23798 3619 23863 3644 1 Vctrl
port 3 n
rlabel metal1 22874 287 22920 322 1 vbn
port 8 n
rlabel metal1 24102 65 24181 123 1 Gnd
port 9 n
rlabel metal1 29083 3626 29148 3651 1 Vctrl
port 3 n
rlabel metal2 4485 2055 5051 2373 1 inp
port 10 n
rlabel metal2 2574 2059 3140 2377 1 inn
port 11 n
<< end >>
