magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect -296 -1219 296 1219
<< pmoslvt >>
rect -100 -1000 100 1000
<< pdiff >>
rect -158 969 -100 1000
rect -158 935 -146 969
rect -112 935 -100 969
rect -158 901 -100 935
rect -158 867 -146 901
rect -112 867 -100 901
rect -158 833 -100 867
rect -158 799 -146 833
rect -112 799 -100 833
rect -158 765 -100 799
rect -158 731 -146 765
rect -112 731 -100 765
rect -158 697 -100 731
rect -158 663 -146 697
rect -112 663 -100 697
rect -158 629 -100 663
rect -158 595 -146 629
rect -112 595 -100 629
rect -158 561 -100 595
rect -158 527 -146 561
rect -112 527 -100 561
rect -158 493 -100 527
rect -158 459 -146 493
rect -112 459 -100 493
rect -158 425 -100 459
rect -158 391 -146 425
rect -112 391 -100 425
rect -158 357 -100 391
rect -158 323 -146 357
rect -112 323 -100 357
rect -158 289 -100 323
rect -158 255 -146 289
rect -112 255 -100 289
rect -158 221 -100 255
rect -158 187 -146 221
rect -112 187 -100 221
rect -158 153 -100 187
rect -158 119 -146 153
rect -112 119 -100 153
rect -158 85 -100 119
rect -158 51 -146 85
rect -112 51 -100 85
rect -158 17 -100 51
rect -158 -17 -146 17
rect -112 -17 -100 17
rect -158 -51 -100 -17
rect -158 -85 -146 -51
rect -112 -85 -100 -51
rect -158 -119 -100 -85
rect -158 -153 -146 -119
rect -112 -153 -100 -119
rect -158 -187 -100 -153
rect -158 -221 -146 -187
rect -112 -221 -100 -187
rect -158 -255 -100 -221
rect -158 -289 -146 -255
rect -112 -289 -100 -255
rect -158 -323 -100 -289
rect -158 -357 -146 -323
rect -112 -357 -100 -323
rect -158 -391 -100 -357
rect -158 -425 -146 -391
rect -112 -425 -100 -391
rect -158 -459 -100 -425
rect -158 -493 -146 -459
rect -112 -493 -100 -459
rect -158 -527 -100 -493
rect -158 -561 -146 -527
rect -112 -561 -100 -527
rect -158 -595 -100 -561
rect -158 -629 -146 -595
rect -112 -629 -100 -595
rect -158 -663 -100 -629
rect -158 -697 -146 -663
rect -112 -697 -100 -663
rect -158 -731 -100 -697
rect -158 -765 -146 -731
rect -112 -765 -100 -731
rect -158 -799 -100 -765
rect -158 -833 -146 -799
rect -112 -833 -100 -799
rect -158 -867 -100 -833
rect -158 -901 -146 -867
rect -112 -901 -100 -867
rect -158 -935 -100 -901
rect -158 -969 -146 -935
rect -112 -969 -100 -935
rect -158 -1000 -100 -969
rect 100 969 158 1000
rect 100 935 112 969
rect 146 935 158 969
rect 100 901 158 935
rect 100 867 112 901
rect 146 867 158 901
rect 100 833 158 867
rect 100 799 112 833
rect 146 799 158 833
rect 100 765 158 799
rect 100 731 112 765
rect 146 731 158 765
rect 100 697 158 731
rect 100 663 112 697
rect 146 663 158 697
rect 100 629 158 663
rect 100 595 112 629
rect 146 595 158 629
rect 100 561 158 595
rect 100 527 112 561
rect 146 527 158 561
rect 100 493 158 527
rect 100 459 112 493
rect 146 459 158 493
rect 100 425 158 459
rect 100 391 112 425
rect 146 391 158 425
rect 100 357 158 391
rect 100 323 112 357
rect 146 323 158 357
rect 100 289 158 323
rect 100 255 112 289
rect 146 255 158 289
rect 100 221 158 255
rect 100 187 112 221
rect 146 187 158 221
rect 100 153 158 187
rect 100 119 112 153
rect 146 119 158 153
rect 100 85 158 119
rect 100 51 112 85
rect 146 51 158 85
rect 100 17 158 51
rect 100 -17 112 17
rect 146 -17 158 17
rect 100 -51 158 -17
rect 100 -85 112 -51
rect 146 -85 158 -51
rect 100 -119 158 -85
rect 100 -153 112 -119
rect 146 -153 158 -119
rect 100 -187 158 -153
rect 100 -221 112 -187
rect 146 -221 158 -187
rect 100 -255 158 -221
rect 100 -289 112 -255
rect 146 -289 158 -255
rect 100 -323 158 -289
rect 100 -357 112 -323
rect 146 -357 158 -323
rect 100 -391 158 -357
rect 100 -425 112 -391
rect 146 -425 158 -391
rect 100 -459 158 -425
rect 100 -493 112 -459
rect 146 -493 158 -459
rect 100 -527 158 -493
rect 100 -561 112 -527
rect 146 -561 158 -527
rect 100 -595 158 -561
rect 100 -629 112 -595
rect 146 -629 158 -595
rect 100 -663 158 -629
rect 100 -697 112 -663
rect 146 -697 158 -663
rect 100 -731 158 -697
rect 100 -765 112 -731
rect 146 -765 158 -731
rect 100 -799 158 -765
rect 100 -833 112 -799
rect 146 -833 158 -799
rect 100 -867 158 -833
rect 100 -901 112 -867
rect 146 -901 158 -867
rect 100 -935 158 -901
rect 100 -969 112 -935
rect 146 -969 158 -935
rect 100 -1000 158 -969
<< pdiffc >>
rect -146 935 -112 969
rect -146 867 -112 901
rect -146 799 -112 833
rect -146 731 -112 765
rect -146 663 -112 697
rect -146 595 -112 629
rect -146 527 -112 561
rect -146 459 -112 493
rect -146 391 -112 425
rect -146 323 -112 357
rect -146 255 -112 289
rect -146 187 -112 221
rect -146 119 -112 153
rect -146 51 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -51
rect -146 -153 -112 -119
rect -146 -221 -112 -187
rect -146 -289 -112 -255
rect -146 -357 -112 -323
rect -146 -425 -112 -391
rect -146 -493 -112 -459
rect -146 -561 -112 -527
rect -146 -629 -112 -595
rect -146 -697 -112 -663
rect -146 -765 -112 -731
rect -146 -833 -112 -799
rect -146 -901 -112 -867
rect -146 -969 -112 -935
rect 112 935 146 969
rect 112 867 146 901
rect 112 799 146 833
rect 112 731 146 765
rect 112 663 146 697
rect 112 595 146 629
rect 112 527 146 561
rect 112 459 146 493
rect 112 391 146 425
rect 112 323 146 357
rect 112 255 146 289
rect 112 187 146 221
rect 112 119 146 153
rect 112 51 146 85
rect 112 -17 146 17
rect 112 -85 146 -51
rect 112 -153 146 -119
rect 112 -221 146 -187
rect 112 -289 146 -255
rect 112 -357 146 -323
rect 112 -425 146 -391
rect 112 -493 146 -459
rect 112 -561 146 -527
rect 112 -629 146 -595
rect 112 -697 146 -663
rect 112 -765 146 -731
rect 112 -833 146 -799
rect 112 -901 146 -867
rect 112 -969 146 -935
<< nsubdiff >>
rect -260 1149 -153 1183
rect -119 1149 -85 1183
rect -51 1149 -17 1183
rect 17 1149 51 1183
rect 85 1149 119 1183
rect 153 1149 260 1183
rect -260 1071 -226 1149
rect -260 1003 -226 1037
rect 226 1071 260 1149
rect 226 1003 260 1037
rect -260 935 -226 969
rect -260 867 -226 901
rect -260 799 -226 833
rect -260 731 -226 765
rect -260 663 -226 697
rect -260 595 -226 629
rect -260 527 -226 561
rect -260 459 -226 493
rect -260 391 -226 425
rect -260 323 -226 357
rect -260 255 -226 289
rect -260 187 -226 221
rect -260 119 -226 153
rect -260 51 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect -260 -153 -226 -119
rect -260 -221 -226 -187
rect -260 -289 -226 -255
rect -260 -357 -226 -323
rect -260 -425 -226 -391
rect -260 -493 -226 -459
rect -260 -561 -226 -527
rect -260 -629 -226 -595
rect -260 -697 -226 -663
rect -260 -765 -226 -731
rect -260 -833 -226 -799
rect -260 -901 -226 -867
rect -260 -969 -226 -935
rect 226 935 260 969
rect 226 867 260 901
rect 226 799 260 833
rect 226 731 260 765
rect 226 663 260 697
rect 226 595 260 629
rect 226 527 260 561
rect 226 459 260 493
rect 226 391 260 425
rect 226 323 260 357
rect 226 255 260 289
rect 226 187 260 221
rect 226 119 260 153
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -153 260 -119
rect 226 -221 260 -187
rect 226 -289 260 -255
rect 226 -357 260 -323
rect 226 -425 260 -391
rect 226 -493 260 -459
rect 226 -561 260 -527
rect 226 -629 260 -595
rect 226 -697 260 -663
rect 226 -765 260 -731
rect 226 -833 260 -799
rect 226 -901 260 -867
rect 226 -969 260 -935
rect -260 -1037 -226 -1003
rect -260 -1149 -226 -1071
rect 226 -1037 260 -1003
rect 226 -1149 260 -1071
rect -260 -1183 -153 -1149
rect -119 -1183 -85 -1149
rect -51 -1183 -17 -1149
rect 17 -1183 51 -1149
rect 85 -1183 119 -1149
rect 153 -1183 260 -1149
<< nsubdiffcont >>
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect -260 1037 -226 1071
rect -260 969 -226 1003
rect 226 1037 260 1071
rect -260 901 -226 935
rect -260 833 -226 867
rect -260 765 -226 799
rect -260 697 -226 731
rect -260 629 -226 663
rect -260 561 -226 595
rect -260 493 -226 527
rect -260 425 -226 459
rect -260 357 -226 391
rect -260 289 -226 323
rect -260 221 -226 255
rect -260 153 -226 187
rect -260 85 -226 119
rect -260 17 -226 51
rect -260 -51 -226 -17
rect -260 -119 -226 -85
rect -260 -187 -226 -153
rect -260 -255 -226 -221
rect -260 -323 -226 -289
rect -260 -391 -226 -357
rect -260 -459 -226 -425
rect -260 -527 -226 -493
rect -260 -595 -226 -561
rect -260 -663 -226 -629
rect -260 -731 -226 -697
rect -260 -799 -226 -765
rect -260 -867 -226 -833
rect -260 -935 -226 -901
rect -260 -1003 -226 -969
rect 226 969 260 1003
rect 226 901 260 935
rect 226 833 260 867
rect 226 765 260 799
rect 226 697 260 731
rect 226 629 260 663
rect 226 561 260 595
rect 226 493 260 527
rect 226 425 260 459
rect 226 357 260 391
rect 226 289 260 323
rect 226 221 260 255
rect 226 153 260 187
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect 226 -119 260 -85
rect 226 -187 260 -153
rect 226 -255 260 -221
rect 226 -323 260 -289
rect 226 -391 260 -357
rect 226 -459 260 -425
rect 226 -527 260 -493
rect 226 -595 260 -561
rect 226 -663 260 -629
rect 226 -731 260 -697
rect 226 -799 260 -765
rect 226 -867 260 -833
rect 226 -935 260 -901
rect -260 -1071 -226 -1037
rect 226 -1003 260 -969
rect 226 -1071 260 -1037
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
<< poly >>
rect -100 1081 100 1097
rect -100 1047 -51 1081
rect -17 1047 17 1081
rect 51 1047 100 1081
rect -100 1000 100 1047
rect -100 -1047 100 -1000
rect -100 -1081 -51 -1047
rect -17 -1081 17 -1047
rect 51 -1081 100 -1047
rect -100 -1097 100 -1081
<< polycont >>
rect -51 1047 -17 1081
rect 17 1047 51 1081
rect -51 -1081 -17 -1047
rect 17 -1081 51 -1047
<< locali >>
rect -260 1149 -153 1183
rect -119 1149 -85 1183
rect -51 1149 -17 1183
rect 17 1149 51 1183
rect 85 1149 119 1183
rect 153 1149 260 1183
rect -260 1071 -226 1149
rect -100 1047 -51 1081
rect -17 1047 17 1081
rect 51 1047 100 1081
rect 226 1071 260 1149
rect -260 1003 -226 1037
rect -260 935 -226 969
rect -260 867 -226 901
rect -260 799 -226 833
rect -260 731 -226 765
rect -260 663 -226 697
rect -260 595 -226 629
rect -260 527 -226 561
rect -260 459 -226 493
rect -260 391 -226 425
rect -260 323 -226 357
rect -260 255 -226 289
rect -260 187 -226 221
rect -260 119 -226 153
rect -260 51 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect -260 -153 -226 -119
rect -260 -221 -226 -187
rect -260 -289 -226 -255
rect -260 -357 -226 -323
rect -260 -425 -226 -391
rect -260 -493 -226 -459
rect -260 -561 -226 -527
rect -260 -629 -226 -595
rect -260 -697 -226 -663
rect -260 -765 -226 -731
rect -260 -833 -226 -799
rect -260 -901 -226 -867
rect -260 -969 -226 -935
rect -260 -1037 -226 -1003
rect -146 969 -112 1004
rect -146 901 -112 935
rect -146 833 -112 867
rect -146 765 -112 799
rect -146 697 -112 731
rect -146 629 -112 663
rect -146 561 -112 595
rect -146 493 -112 527
rect -146 425 -112 459
rect -146 357 -112 391
rect -146 289 -112 323
rect -146 221 -112 255
rect -146 153 -112 187
rect -146 85 -112 119
rect -146 17 -112 51
rect -146 -51 -112 -17
rect -146 -119 -112 -85
rect -146 -187 -112 -153
rect -146 -255 -112 -221
rect -146 -323 -112 -289
rect -146 -391 -112 -357
rect -146 -459 -112 -425
rect -146 -527 -112 -493
rect -146 -595 -112 -561
rect -146 -663 -112 -629
rect -146 -731 -112 -697
rect -146 -799 -112 -765
rect -146 -867 -112 -833
rect -146 -935 -112 -901
rect -146 -1004 -112 -969
rect 112 969 146 1004
rect 112 901 146 935
rect 112 833 146 867
rect 112 765 146 799
rect 112 697 146 731
rect 112 629 146 663
rect 112 561 146 595
rect 112 493 146 527
rect 112 425 146 459
rect 112 357 146 391
rect 112 289 146 323
rect 112 221 146 255
rect 112 153 146 187
rect 112 85 146 119
rect 112 17 146 51
rect 112 -51 146 -17
rect 112 -119 146 -85
rect 112 -187 146 -153
rect 112 -255 146 -221
rect 112 -323 146 -289
rect 112 -391 146 -357
rect 112 -459 146 -425
rect 112 -527 146 -493
rect 112 -595 146 -561
rect 112 -663 146 -629
rect 112 -731 146 -697
rect 112 -799 146 -765
rect 112 -867 146 -833
rect 112 -935 146 -901
rect 112 -1004 146 -969
rect 226 1003 260 1037
rect 226 935 260 969
rect 226 867 260 901
rect 226 799 260 833
rect 226 731 260 765
rect 226 663 260 697
rect 226 595 260 629
rect 226 527 260 561
rect 226 459 260 493
rect 226 391 260 425
rect 226 323 260 357
rect 226 255 260 289
rect 226 187 260 221
rect 226 119 260 153
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -153 260 -119
rect 226 -221 260 -187
rect 226 -289 260 -255
rect 226 -357 260 -323
rect 226 -425 260 -391
rect 226 -493 260 -459
rect 226 -561 260 -527
rect 226 -629 260 -595
rect 226 -697 260 -663
rect 226 -765 260 -731
rect 226 -833 260 -799
rect 226 -901 260 -867
rect 226 -969 260 -935
rect 226 -1037 260 -1003
rect -260 -1149 -226 -1071
rect -100 -1081 -51 -1047
rect -17 -1081 17 -1047
rect 51 -1081 100 -1047
rect 226 -1149 260 -1071
rect -260 -1183 -153 -1149
rect -119 -1183 -85 -1149
rect -51 -1183 -17 -1149
rect 17 -1183 51 -1149
rect 85 -1183 119 -1149
rect 153 -1183 260 -1149
<< properties >>
string FIXED_BBOX -243 -1166 243 1166
<< end >>
