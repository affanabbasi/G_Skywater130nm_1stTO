magic
tech sky130A
magscale 1 2
timestamp 1608071797
<< nwell >>
rect -1770 -919 1770 919
<< pmos >>
rect -1574 -700 -1174 700
rect -1116 -700 -716 700
rect -658 -700 -258 700
rect -200 -700 200 700
rect 258 -700 658 700
rect 716 -700 1116 700
rect 1174 -700 1574 700
<< pdiff >>
rect -1632 688 -1574 700
rect -1632 -688 -1620 688
rect -1586 -688 -1574 688
rect -1632 -700 -1574 -688
rect -1174 688 -1116 700
rect -1174 -688 -1162 688
rect -1128 -688 -1116 688
rect -1174 -700 -1116 -688
rect -716 688 -658 700
rect -716 -688 -704 688
rect -670 -688 -658 688
rect -716 -700 -658 -688
rect -258 688 -200 700
rect -258 -688 -246 688
rect -212 -688 -200 688
rect -258 -700 -200 -688
rect 200 688 258 700
rect 200 -688 212 688
rect 246 -688 258 688
rect 200 -700 258 -688
rect 658 688 716 700
rect 658 -688 670 688
rect 704 -688 716 688
rect 658 -700 716 -688
rect 1116 688 1174 700
rect 1116 -688 1128 688
rect 1162 -688 1174 688
rect 1116 -700 1174 -688
rect 1574 688 1632 700
rect 1574 -688 1586 688
rect 1620 -688 1632 688
rect 1574 -700 1632 -688
<< pdiffc >>
rect -1620 -688 -1586 688
rect -1162 -688 -1128 688
rect -704 -688 -670 688
rect -246 -688 -212 688
rect 212 -688 246 688
rect 670 -688 704 688
rect 1128 -688 1162 688
rect 1586 -688 1620 688
<< nsubdiff >>
rect -1734 849 -1638 883
rect 1638 849 1734 883
rect -1734 787 -1700 849
rect 1700 787 1734 849
rect -1734 -849 -1700 -787
rect 1700 -849 1734 -787
rect -1734 -883 -1638 -849
rect 1638 -883 1734 -849
<< nsubdiffcont >>
rect -1638 849 1638 883
rect -1734 -787 -1700 787
rect 1700 -787 1734 787
rect -1638 -883 1638 -849
<< poly >>
rect -1574 781 -1174 797
rect -1574 747 -1558 781
rect -1190 747 -1174 781
rect -1574 700 -1174 747
rect -1116 781 -716 797
rect -1116 747 -1100 781
rect -732 747 -716 781
rect -1116 700 -716 747
rect -658 781 -258 797
rect -658 747 -642 781
rect -274 747 -258 781
rect -658 700 -258 747
rect -200 781 200 797
rect -200 747 -184 781
rect 184 747 200 781
rect -200 700 200 747
rect 258 781 658 797
rect 258 747 274 781
rect 642 747 658 781
rect 258 700 658 747
rect 716 781 1116 797
rect 716 747 732 781
rect 1100 747 1116 781
rect 716 700 1116 747
rect 1174 781 1574 797
rect 1174 747 1190 781
rect 1558 747 1574 781
rect 1174 700 1574 747
rect -1574 -747 -1174 -700
rect -1574 -781 -1558 -747
rect -1190 -781 -1174 -747
rect -1574 -797 -1174 -781
rect -1116 -747 -716 -700
rect -1116 -781 -1100 -747
rect -732 -781 -716 -747
rect -1116 -797 -716 -781
rect -658 -747 -258 -700
rect -658 -781 -642 -747
rect -274 -781 -258 -747
rect -658 -797 -258 -781
rect -200 -747 200 -700
rect -200 -781 -184 -747
rect 184 -781 200 -747
rect -200 -797 200 -781
rect 258 -747 658 -700
rect 258 -781 274 -747
rect 642 -781 658 -747
rect 258 -797 658 -781
rect 716 -747 1116 -700
rect 716 -781 732 -747
rect 1100 -781 1116 -747
rect 716 -797 1116 -781
rect 1174 -747 1574 -700
rect 1174 -781 1190 -747
rect 1558 -781 1574 -747
rect 1174 -797 1574 -781
<< polycont >>
rect -1558 747 -1190 781
rect -1100 747 -732 781
rect -642 747 -274 781
rect -184 747 184 781
rect 274 747 642 781
rect 732 747 1100 781
rect 1190 747 1558 781
rect -1558 -781 -1190 -747
rect -1100 -781 -732 -747
rect -642 -781 -274 -747
rect -184 -781 184 -747
rect 274 -781 642 -747
rect 732 -781 1100 -747
rect 1190 -781 1558 -747
<< locali >>
rect -1734 849 -1638 883
rect 1638 849 1734 883
rect -1734 787 -1700 849
rect 1700 787 1734 849
rect -1574 747 -1558 781
rect -1190 747 -1174 781
rect -1116 747 -1100 781
rect -732 747 -716 781
rect -658 747 -642 781
rect -274 747 -258 781
rect -200 747 -184 781
rect 184 747 200 781
rect 258 747 274 781
rect 642 747 658 781
rect 716 747 732 781
rect 1100 747 1116 781
rect 1174 747 1190 781
rect 1558 747 1574 781
rect -1620 688 -1586 704
rect -1620 -704 -1586 -688
rect -1162 688 -1128 704
rect -1162 -704 -1128 -688
rect -704 688 -670 704
rect -704 -704 -670 -688
rect -246 688 -212 704
rect -246 -704 -212 -688
rect 212 688 246 704
rect 212 -704 246 -688
rect 670 688 704 704
rect 670 -704 704 -688
rect 1128 688 1162 704
rect 1128 -704 1162 -688
rect 1586 688 1620 704
rect 1586 -704 1620 -688
rect -1574 -781 -1558 -747
rect -1190 -781 -1174 -747
rect -1116 -781 -1100 -747
rect -732 -781 -716 -747
rect -658 -781 -642 -747
rect -274 -781 -258 -747
rect -200 -781 -184 -747
rect 184 -781 200 -747
rect 258 -781 274 -747
rect 642 -781 658 -747
rect 716 -781 732 -747
rect 1100 -781 1116 -747
rect 1174 -781 1190 -747
rect 1558 -781 1574 -747
rect -1734 -849 -1700 -787
rect 1700 -849 1734 -787
rect -1734 -883 -1638 -849
rect 1638 -883 1734 -849
<< viali >>
rect -1558 747 -1190 781
rect -1100 747 -732 781
rect -642 747 -274 781
rect -184 747 184 781
rect 274 747 642 781
rect 732 747 1100 781
rect 1190 747 1558 781
rect -1558 -781 -1190 -747
rect -1100 -781 -732 -747
rect -642 -781 -274 -747
rect -184 -781 184 -747
rect 274 -781 642 -747
rect 732 -781 1100 -747
rect 1190 -781 1558 -747
<< metal1 >>
rect -1570 781 -1178 787
rect -1570 747 -1558 781
rect -1190 747 -1178 781
rect -1570 741 -1178 747
rect -1112 781 -720 787
rect -1112 747 -1100 781
rect -732 747 -720 781
rect -1112 741 -720 747
rect -654 781 -262 787
rect -654 747 -642 781
rect -274 747 -262 781
rect -654 741 -262 747
rect -196 781 196 787
rect -196 747 -184 781
rect 184 747 196 781
rect -196 741 196 747
rect 262 781 654 787
rect 262 747 274 781
rect 642 747 654 781
rect 262 741 654 747
rect 720 781 1112 787
rect 720 747 732 781
rect 1100 747 1112 781
rect 720 741 1112 747
rect 1178 781 1570 787
rect 1178 747 1190 781
rect 1558 747 1570 781
rect 1178 741 1570 747
rect -1570 -747 -1178 -741
rect -1570 -781 -1558 -747
rect -1190 -781 -1178 -747
rect -1570 -787 -1178 -781
rect -1112 -747 -720 -741
rect -1112 -781 -1100 -747
rect -732 -781 -720 -747
rect -1112 -787 -720 -781
rect -654 -747 -262 -741
rect -654 -781 -642 -747
rect -274 -781 -262 -747
rect -654 -787 -262 -781
rect -196 -747 196 -741
rect -196 -781 -184 -747
rect 184 -781 196 -747
rect -196 -787 196 -781
rect 262 -747 654 -741
rect 262 -781 274 -747
rect 642 -781 654 -747
rect 262 -787 654 -781
rect 720 -747 1112 -741
rect 720 -781 732 -747
rect 1100 -781 1112 -747
rect 720 -787 1112 -781
rect 1178 -747 1570 -741
rect 1178 -781 1190 -747
rect 1558 -781 1570 -747
rect 1178 -787 1570 -781
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1717 -866 1717 866
string parameters w 7 l 2 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 0 viasrc 0
string library sky130
<< end >>
