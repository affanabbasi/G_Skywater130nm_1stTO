magic
tech sky130A
magscale 1 2
timestamp 1607564249
<< error_s >>
rect 38804 378341 38805 378386
rect 38833 378375 38834 378386
rect 38844 378341 38845 378375
rect 38804 378273 38805 378318
rect 38833 378307 38834 378318
rect 38844 378273 38845 378307
rect 38804 378205 38805 378250
rect 38833 378239 38834 378250
rect 38844 378205 38845 378239
rect 7892 378104 7960 378105
rect 8050 378104 8118 378105
rect 8208 378104 8276 378105
rect 8366 378104 8434 378105
rect 8524 378104 8592 378105
rect 8682 378104 8750 378105
rect 8840 378104 8908 378105
rect 8998 378104 9066 378105
rect 9156 378104 9224 378105
rect 9314 378104 9382 378105
rect 9472 378104 9540 378105
rect 39390 378034 39424 378049
rect 39389 378033 39424 378034
rect 39470 378033 39471 378043
rect 39669 378033 39670 378043
rect 39716 378033 39750 378049
rect 40027 378035 40061 378050
rect 40026 378034 40061 378035
rect 40107 378034 40108 378044
rect 40306 378034 40307 378044
rect 39389 378001 39390 378033
rect 39440 378031 39700 378033
rect 39470 378001 39471 378031
rect 39389 378000 39423 378001
rect 39716 378000 39717 378033
rect 40026 378002 40027 378034
rect 40077 378032 40337 378034
rect 40107 378002 40108 378032
rect 40026 378001 40060 378002
rect 39390 377985 39424 378000
rect 39716 377985 39750 378000
rect 40027 377986 40061 378001
rect 40353 377986 40387 378050
rect 38684 377907 38748 377909
rect 38794 377907 38960 377909
rect 36342 377163 36343 377164
rect 37461 377163 37462 377164
rect 36341 377162 36342 377163
rect 37462 377162 37463 377163
rect 38981 376333 38983 377597
rect 40907 376337 40909 377601
rect 5303 375993 5305 376109
rect 5867 376008 5869 376042
rect 5901 376015 5903 376115
rect 7876 376058 7976 376059
rect 8034 376058 8134 376059
rect 8192 376058 8292 376059
rect 8350 376058 8450 376059
rect 8508 376058 8608 376059
rect 8666 376058 8766 376059
rect 8824 376058 8924 376059
rect 8982 376058 9082 376059
rect 9140 376058 9240 376059
rect 9298 376058 9398 376059
rect 9456 376058 9556 376059
rect 36341 376043 36342 376044
rect 37462 376043 37463 376044
rect 36342 376042 36343 376043
rect 37461 376042 37462 376043
rect 5901 375999 5903 376008
rect 36460 375611 36461 375612
rect 37579 375611 37580 375612
rect 36459 375610 36460 375611
rect 37580 375610 37581 375611
rect 6072 375534 6110 375588
rect 6076 375532 6130 375534
rect 6110 375530 6130 375532
rect 60922 375242 60924 375358
rect 61486 375257 61488 375291
rect 61520 375264 61522 375364
rect 61520 375248 61522 375257
rect 39003 375138 39037 375202
rect 39241 375186 39275 375188
rect 39053 375184 39225 375186
rect 61691 374783 61729 374837
rect 61695 374781 61749 374783
rect 61729 374779 61749 374781
rect 36459 374491 36460 374492
rect 37580 374491 37581 374492
rect 36460 374490 36461 374491
rect 37579 374490 37580 374491
<< nwell >>
rect 39886 377808 39894 378228
<< metal1 >>
rect 226738 -32043 357511 -31948
rect 226738 -32400 354392 -32043
rect 357432 -32400 357511 -32043
rect 226738 -32479 357511 -32400
rect 320307 -32733 322284 -32479
rect 234229 -43727 286945 -40124
rect 234229 -45211 234764 -43727
rect 286475 -45211 286945 -43727
rect 234229 -45806 286945 -45211
<< via1 >>
rect 354392 -32400 357432 -32043
rect 236556 -39428 236637 -39363
rect 234764 -45211 286475 -43727
<< metal2 >>
rect 54068 382528 95797 384682
rect 54068 375428 55689 382528
rect 54068 374841 58946 375428
rect 63466 374856 64082 375443
rect 73283 375165 74904 382528
rect 94176 376752 95797 382528
rect 94176 376165 99689 376752
rect 73283 374578 78161 375165
rect 5151 369751 6242 373268
rect 63369 369751 64414 374079
rect 77713 369751 78139 374217
rect 5151 368243 78139 369751
rect -19560 -21048 173239 -20510
rect -19560 -29114 -19099 -21048
rect -11205 -29114 173239 -21048
rect -19560 -29621 173239 -29114
rect 354300 -32043 357511 -31920
rect 354300 -32400 354392 -32043
rect 357432 -32400 357511 -32043
rect 354300 -33958 357511 -32400
rect 234261 -39363 236666 -38413
rect 234261 -39428 236556 -39363
rect 236637 -39428 236666 -39363
rect 234261 -39463 236666 -39428
rect 234229 -43637 286945 -43222
rect 234229 -45351 234646 -43637
rect 286559 -45351 286945 -43637
rect 234229 -45806 286945 -45351
<< via2 >>
rect -19099 -29114 -11205 -21048
rect 234646 -43727 286559 -43637
rect 234646 -45211 234764 -43727
rect 234764 -45211 286475 -43727
rect 286475 -45211 286559 -43727
rect 234646 -45351 286559 -45211
<< metal3 >>
rect -19560 380290 38105 381411
rect -19560 -21048 -10715 380290
rect -3560 378399 -2469 380290
rect 37014 378002 38105 380290
rect 67277 381251 91037 383003
rect 67277 375443 68898 381251
rect 63466 374856 68898 375443
rect 89478 375901 91037 381251
rect 100799 375901 101451 376667
rect 89478 375314 101451 375901
rect 89478 375217 91037 375314
rect 83993 374610 91037 375217
rect -19560 -29114 -19099 -21048
rect -11205 -29114 -10715 -21048
rect -19560 -29621 -10715 -29114
rect 234229 -43530 286945 -43222
rect 234229 -45474 234540 -43530
rect 286648 -45474 286945 -43530
rect 234229 -45806 286945 -45474
<< via3 >>
rect 234540 -43637 286648 -43530
rect 234540 -45351 234646 -43637
rect 234646 -45351 286559 -43637
rect 286559 -45351 286648 -43637
rect 234540 -45474 286648 -45351
<< metal4 >>
rect 95894 360081 97123 373638
rect -34915 349108 97123 360081
rect -34915 -51999 -25820 349108
rect 185527 -36496 196607 -33773
rect 192914 -51999 196607 -36496
rect 234229 -43417 286945 -43222
rect 234229 -45623 234401 -43417
rect 286756 -45623 286945 -43417
rect 234229 -45806 286945 -45623
rect -34915 -57298 196607 -51999
<< via4 >>
rect 234401 -43530 286756 -43417
rect 234401 -45474 234540 -43530
rect 234540 -45474 286648 -43530
rect 286648 -45474 286756 -43530
rect 234401 -45623 286756 -45474
<< metal5 >>
rect 14438 385214 112146 389734
rect 14438 377432 16116 385214
rect 39590 378351 40052 385214
rect 59233 379762 63127 385214
rect 80138 380492 82041 385214
rect 96486 381115 97126 385214
rect 14470 364767 15874 374282
rect 39447 364767 40212 373690
rect 59219 364767 63111 372295
rect 80247 364767 82311 372084
rect 97955 364767 98612 372645
rect -52977 360247 112178 364767
rect -52977 -43222 -47130 360247
rect 178831 -29552 354135 -24375
rect 238719 -31764 239616 -29552
rect 317049 -34344 317515 -29552
rect 353386 -34766 354135 -29552
rect 184807 -43222 187145 -38239
rect 317046 -43222 317512 -37088
rect 354350 -43222 357843 -36038
rect -52977 -43417 358077 -43222
rect -52977 -45623 234401 -43417
rect 286756 -45623 358077 -43417
rect -52977 -46201 358077 -45623
use LVDS2_Top  LVDS2_Top_0
timestamp 1607564249
transform 1 0 78399 0 1 375538
box -694 -3510 6019 4973
use LVDSBias_Top  LVDSBias_Top_0
timestamp 1607564249
transform 1 0 39318 0 1 377835
box -3702 -5224 3568 842
use LVDStop  LVDStop_0
timestamp 1607564249
transform 1 0 -2045 0 1 373048
box -1515 0 20087 5918
use PA_1  PA_1_0
timestamp 1606531739
transform 1 0 15084 0 1 -7863
box 0 -31847 352952 379374
use BiasVCO  BiasVCO_0 
timestamp 1607564249
transform 1 0 317789 0 1 -35727
box -743 -1581 14424 3042
use foldedcascode1  foldedcascode1_0
timestamp 1607564249
transform 1 0 100046 0 1 376620
box -3600 -4460 11100 4600
use LVDS1_Top  LVDS1_Top_0
timestamp 1607564249
transform 1 0 59453 0 1 375677
box -1992 -3503 5464 4095
use Delay_Top  Delay_Top_0
timestamp 1607293554
transform 1 0 223681 0 1 -40002
box 3056 -128 65878 14314
use RO  RO_0 
timestamp 1606670916
transform 1 0 354350 0 1 -35359
box -918 -686 4384 1644
<< labels >>
rlabel metal5 350574 -28978 353470 -25117 1 p_vgate
port 1 n
rlabel space 355778 341564 365860 351484 1 pa_vdd
port 2 n
rlabel metal5 15373 386177 18490 389054 1 p_vdd
port 3 n
rlabel metal5 354549 -46011 357666 -43134 1 p_vss
port 4 n
rlabel metal4 -33179 350269 -26691 358785 1 p_isrc
port 5 n
rlabel space 358217 -35355 358690 -34477 1 ro_out
port 6 n
rlabel space 320328 -37256 320662 -36917 1 selfb_vinit
port 7 n
rlabel space 317084 -36228 317493 -35818 1 selfb_vbn
port 8 n
rlabel space 317085 -35318 317474 -34934 1 inv1in
port 9 n
rlabel space 232970 -35488 233359 -35104 1 dvco_outn
port 10 n
rlabel space 229038 -36503 229427 -36119 1 dvco_outp
port 11 n
rlabel metal2 234466 -39151 234911 -38685 1 dvco_vbn
port 12 n
rlabel space 183113 -31067 183558 -30601 1 pa_rnode
port 13 n
rlabel space 164633 -17763 168822 -12003 1 pa_out
port 14 n
rlabel space 17146 375540 17814 376244 1 lvdstop_out
port 15 n
rlabel space -3189 376859 -2851 377183 1 lvdstop_inp
port 16 n
rlabel space -3154 375288 -2816 375612 1 lvdstop_inn
port 17 n
rlabel metal2 5345 368405 6973 369580 1 lvds_vbiasn
port 18 n
rlabel space 35734 376337 35891 376501 1 lvdsbias_inp
port 19 n
rlabel space 35734 374811 35891 374975 1 lvdsbias_inn
port 20 n
rlabel space 42549 376929 42755 377132 1 lvdsbias_vp
port 21 n
rlabel space 42549 375903 42755 376106 1 lvdsbias_vn
port 22 n
rlabel space 57700 376413 58664 377615 1 lvds1_on1a
port 23 n
rlabel space 63680 376312 64644 377514 1 lvds1_on2a
port 24 n
rlabel metal2 54419 382763 57012 384413 1 lvds_vp
port 25 n
rlabel metal3 67486 381298 70113 382427 1 lvds_vn
port 26 n
rlabel space 77777 375393 78027 375661 1 lvds2_on2b
port 27 n
rlabel space 84072 375393 84322 375661 1 lvds2_on1b
port 28 n
rlabel space 108574 377846 109032 378241 1 fc_out
port 29 n
rlabel metal2 354618 -33602 357246 -32661 1 ocs_vdd
port 30 n
<< end >>
