magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect 1370 1334 1460 1460
<< locali >>
rect 186 2022 3244 2060
rect 186 1988 261 2022
rect 295 2020 2477 2022
rect 295 2016 2037 2020
rect 295 1988 571 2016
rect 186 1982 571 1988
rect 605 2010 1363 2016
rect 605 1982 887 2010
rect 186 1976 887 1982
rect 921 1982 1363 2010
rect 1397 1986 2037 2016
rect 2071 1988 2477 2020
rect 2511 1988 2771 2022
rect 2805 1988 3073 2022
rect 3107 1988 3244 2022
rect 2071 1986 3244 1988
rect 1397 1982 3244 1986
rect 921 1976 3244 1982
rect 186 1936 3244 1976
rect 2316 1573 2386 1592
rect 2316 1539 2334 1573
rect 2368 1539 2386 1573
rect 2316 1501 2386 1539
rect 2316 1467 2334 1501
rect 2368 1467 2386 1501
rect 2316 1429 2386 1467
rect 2316 1395 2334 1429
rect 2368 1395 2386 1429
rect 2316 1357 2386 1395
rect 2316 1323 2334 1357
rect 2368 1323 2386 1357
rect 2316 1285 2386 1323
rect 2316 1251 2334 1285
rect 2368 1251 2386 1285
rect 2316 1213 2386 1251
rect 2316 1179 2334 1213
rect 2368 1179 2386 1213
rect 2316 1160 2386 1179
rect 2634 1573 2704 1592
rect 2634 1539 2652 1573
rect 2686 1539 2704 1573
rect 2634 1501 2704 1539
rect 2634 1467 2652 1501
rect 2686 1467 2704 1501
rect 2634 1429 2704 1467
rect 2634 1395 2652 1429
rect 2686 1395 2704 1429
rect 2634 1357 2704 1395
rect 2634 1323 2652 1357
rect 2686 1323 2704 1357
rect 2634 1285 2704 1323
rect 2634 1251 2652 1285
rect 2686 1251 2704 1285
rect 2634 1213 2704 1251
rect 2634 1179 2652 1213
rect 2686 1179 2704 1213
rect 2634 1160 2704 1179
rect 2952 1573 3022 1592
rect 2952 1539 2970 1573
rect 3004 1539 3022 1573
rect 2952 1501 3022 1539
rect 2952 1467 2970 1501
rect 3004 1467 3022 1501
rect 2952 1429 3022 1467
rect 2952 1395 2970 1429
rect 3004 1395 3022 1429
rect 2952 1357 3022 1395
rect 2952 1323 2970 1357
rect 3004 1323 3022 1357
rect 2952 1285 3022 1323
rect 2952 1251 2970 1285
rect 3004 1251 3022 1285
rect 2952 1213 3022 1251
rect 2952 1179 2970 1213
rect 3004 1179 3022 1213
rect 2952 1160 3022 1179
rect 3270 1573 3340 1592
rect 3270 1539 3288 1573
rect 3322 1539 3340 1573
rect 3270 1501 3340 1539
rect 3270 1467 3288 1501
rect 3322 1467 3340 1501
rect 3270 1429 3340 1467
rect 3270 1395 3288 1429
rect 3322 1395 3340 1429
rect 3270 1357 3340 1395
rect 3270 1323 3288 1357
rect 3322 1323 3340 1357
rect 3270 1285 3340 1323
rect 3270 1251 3288 1285
rect 3322 1251 3340 1285
rect 3270 1213 3340 1251
rect 3270 1179 3288 1213
rect 3322 1179 3340 1213
rect 3270 1160 3340 1179
rect 490 -908 493 -874
rect 527 -908 565 -874
rect 599 -908 637 -874
rect 671 -908 709 -874
rect 743 -908 781 -874
rect 815 -908 853 -874
rect 887 -908 925 -874
rect 959 -908 997 -874
rect 1031 -908 1069 -874
rect 1103 -908 1141 -874
rect 1175 -908 1213 -874
rect 1247 -908 1285 -874
rect 1319 -908 1357 -874
rect 1391 -908 1429 -874
rect 1463 -908 1466 -874
rect 406 -959 440 -936
rect 406 -1031 440 -993
rect 406 -1103 440 -1065
rect 406 -1175 440 -1137
rect 406 -1247 440 -1209
rect 406 -1304 440 -1281
rect 1516 -959 1550 -936
rect 1516 -1031 1550 -993
rect 1516 -1103 1550 -1065
rect 1516 -1175 1550 -1137
rect 1516 -1247 1550 -1209
rect 1516 -1304 1550 -1281
rect 1968 -947 2002 -924
rect 1968 -1019 2002 -981
rect 1968 -1091 2002 -1053
rect 1968 -1163 2002 -1125
rect 1968 -1235 2002 -1197
rect 1968 -1292 2002 -1269
rect 934 -1366 949 -1332
rect 983 -1366 1021 -1332
rect 1055 -1366 1070 -1332
rect 2494 -1354 2507 -1320
rect 2541 -1354 2579 -1320
rect 2613 -1354 2626 -1320
rect 400 -1480 421 -1446
rect 455 -1480 493 -1446
rect 527 -1480 565 -1446
rect 599 -1480 637 -1446
rect 671 -1480 709 -1446
rect 743 -1480 781 -1446
rect 815 -1480 853 -1446
rect 887 -1480 925 -1446
rect 959 -1480 997 -1446
rect 1031 -1480 1069 -1446
rect 1103 -1480 1141 -1446
rect 1175 -1480 1213 -1446
rect 1247 -1480 1285 -1446
rect 1319 -1480 1357 -1446
rect 1391 -1480 1429 -1446
rect 1463 -1480 1501 -1446
rect 1535 -1480 1556 -1446
rect 1962 -1468 1983 -1434
rect 2017 -1468 2055 -1434
rect 2089 -1468 2127 -1434
rect 2161 -1468 2199 -1434
rect 2233 -1468 2271 -1434
rect 2305 -1468 2343 -1434
rect 2377 -1468 2415 -1434
rect 2449 -1468 2487 -1434
rect 2521 -1468 2559 -1434
rect 2593 -1468 2631 -1434
rect 2665 -1468 2703 -1434
rect 2737 -1468 2775 -1434
rect 2809 -1468 2847 -1434
rect 2881 -1468 2919 -1434
rect 2953 -1468 2991 -1434
rect 3025 -1468 3063 -1434
rect 3097 -1468 3118 -1434
<< viali >>
rect 261 1988 295 2022
rect 571 1982 605 2016
rect 887 1976 921 2010
rect 1363 1982 1397 2016
rect 2037 1986 2071 2020
rect 2477 1988 2511 2022
rect 2771 1988 2805 2022
rect 3073 1988 3107 2022
rect 2334 1539 2368 1573
rect 2334 1467 2368 1501
rect 2334 1395 2368 1429
rect 2334 1323 2368 1357
rect 2334 1251 2368 1285
rect 2334 1179 2368 1213
rect 2652 1539 2686 1573
rect 2652 1467 2686 1501
rect 2652 1395 2686 1429
rect 2652 1323 2686 1357
rect 2652 1251 2686 1285
rect 2652 1179 2686 1213
rect 2970 1539 3004 1573
rect 2970 1467 3004 1501
rect 2970 1395 3004 1429
rect 2970 1323 3004 1357
rect 2970 1251 3004 1285
rect 2970 1179 3004 1213
rect 3288 1539 3322 1573
rect 3288 1467 3322 1501
rect 3288 1395 3322 1429
rect 3288 1323 3322 1357
rect 3288 1251 3322 1285
rect 3288 1179 3322 1213
rect 493 -908 527 -874
rect 565 -908 599 -874
rect 637 -908 671 -874
rect 709 -908 743 -874
rect 781 -908 815 -874
rect 853 -908 887 -874
rect 925 -908 959 -874
rect 997 -908 1031 -874
rect 1069 -908 1103 -874
rect 1141 -908 1175 -874
rect 1213 -908 1247 -874
rect 1285 -908 1319 -874
rect 1357 -908 1391 -874
rect 1429 -908 1463 -874
rect 406 -993 440 -959
rect 406 -1065 440 -1031
rect 406 -1137 440 -1103
rect 406 -1209 440 -1175
rect 406 -1281 440 -1247
rect 1516 -993 1550 -959
rect 1516 -1065 1550 -1031
rect 1516 -1137 1550 -1103
rect 1516 -1209 1550 -1175
rect 1516 -1281 1550 -1247
rect 1968 -981 2002 -947
rect 1968 -1053 2002 -1019
rect 1968 -1125 2002 -1091
rect 1968 -1197 2002 -1163
rect 1968 -1269 2002 -1235
rect 949 -1366 983 -1332
rect 1021 -1366 1055 -1332
rect 2507 -1354 2541 -1320
rect 2579 -1354 2613 -1320
rect 421 -1480 455 -1446
rect 493 -1480 527 -1446
rect 565 -1480 599 -1446
rect 637 -1480 671 -1446
rect 709 -1480 743 -1446
rect 781 -1480 815 -1446
rect 853 -1480 887 -1446
rect 925 -1480 959 -1446
rect 997 -1480 1031 -1446
rect 1069 -1480 1103 -1446
rect 1141 -1480 1175 -1446
rect 1213 -1480 1247 -1446
rect 1285 -1480 1319 -1446
rect 1357 -1480 1391 -1446
rect 1429 -1480 1463 -1446
rect 1501 -1480 1535 -1446
rect 1983 -1468 2017 -1434
rect 2055 -1468 2089 -1434
rect 2127 -1468 2161 -1434
rect 2199 -1468 2233 -1434
rect 2271 -1468 2305 -1434
rect 2343 -1468 2377 -1434
rect 2415 -1468 2449 -1434
rect 2487 -1468 2521 -1434
rect 2559 -1468 2593 -1434
rect 2631 -1468 2665 -1434
rect 2703 -1468 2737 -1434
rect 2775 -1468 2809 -1434
rect 2847 -1468 2881 -1434
rect 2919 -1468 2953 -1434
rect 2991 -1468 3025 -1434
rect 3063 -1468 3097 -1434
<< metal1 >>
rect 94 2106 3230 2114
rect 94 2047 3360 2106
rect 94 1931 156 2047
rect 3280 1931 3360 2047
rect 94 1921 3360 1931
rect 206 1888 3360 1921
rect 2004 1573 2414 1610
rect 2004 1539 2334 1573
rect 2368 1539 2414 1573
rect 1196 1521 1428 1538
rect 1196 1213 1204 1521
rect 1384 1213 1428 1521
rect 2004 1523 2414 1539
rect 2004 1221 2062 1523
rect 1196 1148 1428 1213
rect 2002 1215 2062 1221
rect 2242 1501 2414 1523
rect 2242 1467 2334 1501
rect 2368 1467 2414 1501
rect 2242 1429 2414 1467
rect 2242 1395 2334 1429
rect 2368 1395 2414 1429
rect 2242 1357 2414 1395
rect 2242 1323 2334 1357
rect 2368 1323 2414 1357
rect 2242 1285 2414 1323
rect 2242 1251 2334 1285
rect 2368 1251 2414 1285
rect 2242 1215 2414 1251
rect 2002 1213 2414 1215
rect 2002 1193 2334 1213
rect 2004 1142 2032 1193
rect 2076 1179 2334 1193
rect 2368 1179 2414 1213
rect 2076 1142 2414 1179
rect 2616 1573 3040 1616
rect 2616 1539 2652 1573
rect 2686 1539 2970 1573
rect 3004 1539 3040 1573
rect 2616 1501 3040 1539
rect 2616 1467 2652 1501
rect 2686 1467 2970 1501
rect 3004 1467 3040 1501
rect 2616 1429 3040 1467
rect 2616 1395 2652 1429
rect 2686 1395 2970 1429
rect 3004 1395 3040 1429
rect 2616 1357 3040 1395
rect 2616 1323 2652 1357
rect 2686 1323 2970 1357
rect 3004 1323 3040 1357
rect 2616 1285 3040 1323
rect 2616 1251 2652 1285
rect 2686 1251 2970 1285
rect 3004 1251 3040 1285
rect 2616 1213 3040 1251
rect 2616 1179 2652 1213
rect 2686 1179 2970 1213
rect 3004 1179 3040 1213
rect 2616 1142 3040 1179
rect 3254 1573 3360 1888
rect 3254 1539 3288 1573
rect 3322 1539 3360 1573
rect 3254 1501 3360 1539
rect 3254 1467 3288 1501
rect 3322 1467 3360 1501
rect 3254 1429 3360 1467
rect 3254 1395 3288 1429
rect 3322 1395 3360 1429
rect 3254 1357 3360 1395
rect 3254 1323 3288 1357
rect 3322 1323 3360 1357
rect 3254 1285 3360 1323
rect 3254 1251 3288 1285
rect 3322 1251 3360 1285
rect 3254 1213 3360 1251
rect 3254 1179 3288 1213
rect 3322 1179 3360 1213
rect 3254 1144 3360 1179
rect 1372 -470 1440 -466
rect 1372 -522 1381 -470
rect 1433 -522 1440 -470
rect 1372 -526 1440 -522
rect 1972 -487 2034 -474
rect 1972 -539 1978 -487
rect 2030 -539 2034 -487
rect 1972 -554 2034 -539
rect 384 -874 1566 -858
rect 384 -908 493 -874
rect 527 -908 565 -874
rect 599 -908 637 -874
rect 671 -908 709 -874
rect 743 -908 781 -874
rect 815 -908 853 -874
rect 887 -908 925 -874
rect 959 -908 997 -874
rect 1031 -908 1069 -874
rect 1103 -908 1141 -874
rect 1175 -908 1213 -874
rect 1247 -908 1285 -874
rect 1319 -908 1357 -874
rect 1391 -908 1429 -874
rect 1463 -902 1566 -874
rect 1463 -908 2012 -902
rect 384 -922 2012 -908
rect 384 -959 470 -922
rect 384 -993 406 -959
rect 440 -993 470 -959
rect 384 -1031 470 -993
rect 384 -1065 406 -1031
rect 440 -1065 470 -1031
rect 384 -1103 470 -1065
rect 384 -1137 406 -1103
rect 440 -1137 470 -1103
rect 384 -1175 470 -1137
rect 384 -1209 406 -1175
rect 440 -1209 470 -1175
rect 384 -1247 470 -1209
rect 384 -1281 406 -1247
rect 440 -1281 470 -1247
rect 384 -1320 470 -1281
rect 1510 -947 2012 -922
rect 1510 -959 1968 -947
rect 1510 -993 1516 -959
rect 1550 -981 1968 -959
rect 2002 -981 2012 -947
rect 1550 -993 2012 -981
rect 1510 -1001 2012 -993
rect 1510 -1031 1724 -1001
rect 1510 -1065 1516 -1031
rect 1550 -1053 1724 -1031
rect 1776 -1019 2012 -1001
rect 1776 -1053 1968 -1019
rect 2002 -1053 2012 -1019
rect 1550 -1065 2012 -1053
rect 1510 -1103 1724 -1065
rect 1510 -1137 1516 -1103
rect 1550 -1117 1724 -1103
rect 1776 -1091 2012 -1065
rect 1776 -1117 1968 -1091
rect 1550 -1125 1968 -1117
rect 2002 -1125 2012 -1091
rect 1550 -1129 2012 -1125
rect 1550 -1137 1724 -1129
rect 1510 -1175 1724 -1137
rect 1510 -1209 1516 -1175
rect 1550 -1181 1724 -1175
rect 1776 -1163 2012 -1129
rect 1776 -1181 1968 -1163
rect 1550 -1193 1968 -1181
rect 1550 -1209 1724 -1193
rect 1510 -1245 1724 -1209
rect 1776 -1197 1968 -1193
rect 2002 -1197 2012 -1163
rect 1776 -1235 2012 -1197
rect 1776 -1245 1968 -1235
rect 1510 -1247 1968 -1245
rect 1510 -1281 1516 -1247
rect 1550 -1269 1968 -1247
rect 2002 -1269 2012 -1235
rect 1550 -1281 2012 -1269
rect 1510 -1326 2012 -1281
rect 2436 -1320 2714 -1312
rect 884 -1332 1132 -1326
rect 884 -1366 949 -1332
rect 983 -1366 1021 -1332
rect 1055 -1366 1132 -1332
rect 884 -1402 1132 -1366
rect 2436 -1354 2507 -1320
rect 2541 -1354 2579 -1320
rect 2613 -1354 2714 -1320
rect 350 -1404 1668 -1402
rect 2436 -1404 2714 -1354
rect 3030 -1404 3146 -1402
rect 350 -1434 3146 -1404
rect 350 -1446 1983 -1434
rect 350 -1480 421 -1446
rect 455 -1480 493 -1446
rect 527 -1480 565 -1446
rect 599 -1480 637 -1446
rect 671 -1480 709 -1446
rect 743 -1480 781 -1446
rect 815 -1480 853 -1446
rect 887 -1480 925 -1446
rect 959 -1480 997 -1446
rect 1031 -1480 1069 -1446
rect 1103 -1480 1141 -1446
rect 1175 -1480 1213 -1446
rect 1247 -1480 1285 -1446
rect 1319 -1480 1357 -1446
rect 1391 -1480 1429 -1446
rect 1463 -1480 1501 -1446
rect 1535 -1468 1983 -1446
rect 2017 -1468 2055 -1434
rect 2089 -1468 2127 -1434
rect 2161 -1468 2199 -1434
rect 2233 -1468 2271 -1434
rect 2305 -1468 2343 -1434
rect 2377 -1468 2415 -1434
rect 2449 -1468 2487 -1434
rect 2521 -1468 2559 -1434
rect 2593 -1468 2631 -1434
rect 2665 -1468 2703 -1434
rect 2737 -1468 2775 -1434
rect 2809 -1468 2847 -1434
rect 2881 -1468 2919 -1434
rect 2953 -1468 2991 -1434
rect 3025 -1468 3063 -1434
rect 3097 -1468 3146 -1434
rect 1535 -1480 3146 -1468
rect 350 -2573 3146 -1480
rect 224 -2596 3228 -2573
rect 224 -2712 328 -2596
rect 3132 -2712 3228 -2596
rect 224 -2837 3228 -2712
<< via1 >>
rect 156 2022 3280 2047
rect 156 1988 261 2022
rect 261 1988 295 2022
rect 295 2020 2477 2022
rect 295 2016 2037 2020
rect 295 1988 571 2016
rect 156 1982 571 1988
rect 571 1982 605 2016
rect 605 2010 1363 2016
rect 605 1982 887 2010
rect 156 1976 887 1982
rect 887 1976 921 2010
rect 921 1982 1363 2010
rect 1363 1982 1397 2016
rect 1397 1986 2037 2016
rect 2037 1986 2071 2020
rect 2071 1988 2477 2020
rect 2477 1988 2511 2022
rect 2511 1988 2771 2022
rect 2771 1988 2805 2022
rect 2805 1988 3073 2022
rect 3073 1988 3107 2022
rect 3107 1988 3280 2022
rect 2071 1986 3280 1988
rect 1397 1982 3280 1986
rect 921 1976 3280 1982
rect 156 1931 3280 1976
rect 1204 1213 1384 1521
rect 2062 1215 2242 1523
rect 1381 -522 1433 -470
rect 1978 -539 2030 -487
rect 1724 -1053 1776 -1001
rect 1724 -1117 1776 -1065
rect 1724 -1181 1776 -1129
rect 1724 -1245 1776 -1193
rect 328 -2712 3132 -2596
<< metal2 >>
rect 36 2818 3394 2927
rect 36 2682 117 2818
rect 3293 2682 3394 2818
rect 36 2047 3394 2682
rect 36 1931 156 2047
rect 3280 1931 3394 2047
rect 36 1870 3394 1931
rect -922 1534 1484 1626
rect -922 1238 -834 1534
rect -618 1521 1484 1534
rect -618 1238 1204 1521
rect -922 1213 1204 1238
rect 1384 1213 1484 1521
rect -922 1137 1484 1213
rect 1992 1523 4464 1615
rect 1992 1215 2062 1523
rect 2242 1500 4464 1523
rect 2242 1215 4158 1500
rect 1992 1204 4158 1215
rect 4374 1204 4464 1500
rect 1992 1125 4464 1204
rect -1024 -467 -731 -375
rect 4118 -462 4411 -375
rect 1098 -467 1440 -466
rect -1024 -470 1440 -467
rect -1024 -480 1381 -470
rect -1024 -616 -986 -480
rect -850 -522 1381 -480
rect 1433 -522 1440 -470
rect -850 -526 1440 -522
rect 1966 -480 4411 -462
rect 1966 -487 4156 -480
rect -850 -527 1122 -526
rect -850 -616 -731 -527
rect 1966 -539 1978 -487
rect 2030 -539 4156 -487
rect 1966 -554 4156 -539
rect -1024 -709 -731 -616
rect 4118 -616 4156 -554
rect 4292 -616 4411 -480
rect 4118 -709 4411 -616
rect 1632 -1001 1891 -892
rect 1632 -1053 1724 -1001
rect 1776 -1053 1891 -1001
rect 1632 -1065 1891 -1053
rect 1632 -1117 1724 -1065
rect 1776 -1117 1891 -1065
rect 1632 -1129 1891 -1117
rect 1632 -1181 1724 -1129
rect 1776 -1181 1891 -1129
rect 1632 -1193 1891 -1181
rect 1632 -1245 1724 -1193
rect 1776 -1245 1891 -1193
rect 1632 -1636 1891 -1245
rect 1632 -1754 4391 -1636
rect 1632 -1890 4112 -1754
rect 4248 -1890 4391 -1754
rect 1632 -1999 4391 -1890
rect 151 -2596 3297 -2515
rect 151 -2712 328 -2596
rect 3132 -2712 3297 -2596
rect 151 -2810 333 -2712
rect 3109 -2810 3297 -2712
rect 151 -2900 3297 -2810
<< via2 >>
rect 117 2682 3293 2818
rect -834 1238 -618 1534
rect 4158 1204 4374 1500
rect -986 -616 -850 -480
rect 4156 -616 4292 -480
rect 4112 -1890 4248 -1754
rect 333 -2712 3109 -2674
rect 333 -2810 3109 -2712
<< metal3 >>
rect 36 3024 3394 3193
rect 36 2880 114 3024
rect 3298 2880 3394 3024
rect 36 2818 3394 2880
rect 36 2682 117 2818
rect 3293 2682 3394 2818
rect 36 2592 3394 2682
rect -1334 1582 -555 1768
rect -1334 1198 -1209 1582
rect -745 1534 -555 1582
rect -618 1238 -555 1534
rect -745 1198 -555 1238
rect -1334 1000 -555 1198
rect 4073 1550 4681 1711
rect 4073 1500 4227 1550
rect 4073 1204 4158 1500
rect 4073 1166 4227 1204
rect 4531 1166 4681 1550
rect 4073 1006 4681 1166
rect -1059 -439 -618 -341
rect -1059 -480 -946 -439
rect -1059 -616 -986 -480
rect -1059 -663 -946 -616
rect -722 -663 -618 -439
rect -1059 -750 -618 -663
rect 4083 -439 4524 -341
rect 4083 -480 4196 -439
rect 4083 -616 4156 -480
rect 4083 -663 4196 -616
rect 4420 -663 4524 -439
rect 4083 -750 4524 -663
rect 4003 -1711 4406 -1618
rect 4003 -1935 4095 -1711
rect 4319 -1935 4406 -1711
rect 4003 -2015 4406 -1935
rect 93 -2622 3309 -2475
rect 93 -2846 226 -2622
rect 3170 -2846 3309 -2622
rect 93 -2958 3309 -2846
<< via3 >>
rect 114 2880 3298 3024
rect -1209 1534 -745 1582
rect -1209 1238 -834 1534
rect -834 1238 -745 1534
rect -1209 1198 -745 1238
rect 4227 1500 4531 1550
rect 4227 1204 4374 1500
rect 4374 1204 4531 1500
rect 4227 1166 4531 1204
rect -946 -480 -722 -439
rect -946 -616 -850 -480
rect -850 -616 -722 -480
rect -946 -663 -722 -616
rect 4196 -480 4420 -439
rect 4196 -616 4292 -480
rect 4292 -616 4420 -480
rect 4196 -663 4420 -616
rect 4095 -1754 4319 -1711
rect 4095 -1890 4112 -1754
rect 4112 -1890 4248 -1754
rect 4248 -1890 4319 -1754
rect 4095 -1935 4319 -1890
rect 226 -2674 3170 -2622
rect 226 -2810 333 -2674
rect 333 -2810 3109 -2674
rect 3109 -2810 3170 -2674
rect 226 -2846 3170 -2810
<< metal4 >>
rect 36 3591 3405 3794
rect 36 3355 321 3591
rect 557 3355 641 3591
rect 877 3355 961 3591
rect 1197 3355 1281 3591
rect 1517 3355 1601 3591
rect 1837 3355 1921 3591
rect 2157 3355 2241 3591
rect 2477 3355 2561 3591
rect 2797 3355 2881 3591
rect 3117 3355 3405 3591
rect 36 3024 3405 3355
rect 36 2880 114 3024
rect 3298 2880 3405 3024
rect 36 2750 3405 2880
rect -1611 1650 -555 1941
rect -1611 1094 -1373 1650
rect -817 1582 -555 1650
rect -745 1198 -555 1582
rect -817 1094 -555 1198
rect -1611 804 -555 1094
rect 4033 1752 4785 1804
rect 4033 1662 5000 1752
rect 4033 971 4109 1662
rect 4095 786 4109 971
rect 4985 786 5000 1662
rect 4095 697 5000 786
rect -1073 -438 -598 -321
rect -1073 -674 -961 -438
rect -725 -439 -598 -438
rect -722 -663 -598 -439
rect -725 -674 -598 -663
rect -1073 -761 -598 -674
rect 4069 -438 4544 -321
rect 4069 -674 4181 -438
rect 4417 -439 4544 -438
rect 4420 -663 4544 -439
rect 4417 -674 4544 -663
rect 4069 -761 4544 -674
rect 3977 -1697 4475 -1589
rect 3977 -1711 4105 -1697
rect 3977 -1935 4095 -1711
rect 4341 -1933 4475 -1697
rect 4319 -1935 4475 -1933
rect 3977 -2041 4475 -1935
rect 42 -2621 3389 -2395
rect 42 -2622 320 -2621
rect 556 -2622 640 -2621
rect 876 -2622 960 -2621
rect 1196 -2622 1280 -2621
rect 1516 -2622 1600 -2621
rect 1836 -2622 1920 -2621
rect 2156 -2622 2240 -2621
rect 2476 -2622 2560 -2621
rect 2796 -2622 2880 -2621
rect 3116 -2622 3389 -2621
rect 42 -2846 226 -2622
rect 3170 -2846 3389 -2622
rect 42 -2857 320 -2846
rect 556 -2857 640 -2846
rect 876 -2857 960 -2846
rect 1196 -2857 1280 -2846
rect 1516 -2857 1600 -2846
rect 1836 -2857 1920 -2846
rect 2156 -2857 2240 -2846
rect 2476 -2857 2560 -2846
rect 2796 -2857 2880 -2846
rect 3116 -2857 3389 -2846
rect 42 -3090 3389 -2857
<< via4 >>
rect 321 3355 557 3591
rect 641 3355 877 3591
rect 961 3355 1197 3591
rect 1281 3355 1517 3591
rect 1601 3355 1837 3591
rect 1921 3355 2157 3591
rect 2241 3355 2477 3591
rect 2561 3355 2797 3591
rect 2881 3355 3117 3591
rect -1373 1582 -817 1650
rect -1373 1198 -1209 1582
rect -1209 1198 -817 1582
rect -1373 1094 -817 1198
rect 4109 1550 4985 1662
rect 4109 1166 4227 1550
rect 4227 1166 4531 1550
rect 4531 1166 4985 1550
rect 4109 786 4985 1166
rect -961 -439 -725 -438
rect -961 -663 -946 -439
rect -946 -663 -725 -439
rect -961 -674 -725 -663
rect 4181 -439 4417 -438
rect 4181 -663 4196 -439
rect 4196 -663 4417 -439
rect 4181 -674 4417 -663
rect 4105 -1711 4341 -1697
rect 4105 -1933 4319 -1711
rect 4319 -1933 4341 -1711
rect 320 -2622 556 -2621
rect 640 -2622 876 -2621
rect 960 -2622 1196 -2621
rect 1280 -2622 1516 -2621
rect 1600 -2622 1836 -2621
rect 1920 -2622 2156 -2621
rect 2240 -2622 2476 -2621
rect 2560 -2622 2796 -2621
rect 2880 -2622 3116 -2621
rect 320 -2846 556 -2622
rect 640 -2846 876 -2622
rect 960 -2846 1196 -2622
rect 1280 -2846 1516 -2622
rect 1600 -2846 1836 -2622
rect 1920 -2846 2156 -2622
rect 2240 -2846 2476 -2622
rect 2560 -2846 2796 -2622
rect 2880 -2846 3116 -2622
rect 320 -2857 556 -2846
rect 640 -2857 876 -2846
rect 960 -2857 1196 -2846
rect 1280 -2857 1516 -2846
rect 1600 -2857 1836 -2846
rect 1920 -2857 2156 -2846
rect 2240 -2857 2476 -2846
rect 2560 -2857 2796 -2846
rect 2880 -2857 3116 -2846
<< metal5 >>
rect -220 3591 3674 4095
rect -220 3355 321 3591
rect 557 3355 641 3591
rect 877 3355 961 3591
rect 1197 3355 1281 3591
rect 1517 3355 1601 3591
rect 1837 3355 1921 3591
rect 2157 3355 2241 3591
rect 2477 3355 2561 3591
rect 2797 3355 2881 3591
rect 3117 3355 3674 3591
rect -220 2777 3674 3355
rect -1992 1650 -532 2143
rect -1992 1094 -1373 1650
rect -817 1094 -532 1650
rect -1992 556 -532 1094
rect 3968 1662 5464 2135
rect 3968 786 4109 1662
rect 4985 786 5464 1662
rect 3968 419 5464 786
rect -1122 -438 -508 -257
rect -1122 -674 -961 -438
rect -725 -674 -508 -438
rect -1122 -819 -508 -674
rect 4020 -438 4634 -257
rect 4020 -674 4181 -438
rect 4417 -674 4634 -438
rect 4020 -819 4634 -674
rect 3922 -1697 4565 -1505
rect 3922 -1933 4105 -1697
rect 4341 -1933 4565 -1697
rect 3922 -2087 4565 -1933
rect -136 -2621 3561 -2263
rect -136 -2857 320 -2621
rect 556 -2857 640 -2621
rect 876 -2857 960 -2621
rect 1196 -2857 1280 -2621
rect 1516 -2857 1600 -2621
rect 1836 -2857 1920 -2621
rect 2156 -2857 2240 -2621
rect 2476 -2857 2560 -2621
rect 2796 -2857 2880 -2621
rect 3116 -2857 3561 -2621
rect -136 -3503 3561 -2857
use LVDS1  LVDS1_0
timestamp 1611881054
transform 1 0 0 0 1 0
box -17 -1584 3470 2114
<< labels >>
rlabel metal2 s 1676 1966 1770 2038 4 Vdd
port 1 nsew
rlabel metal1 s 2018 1326 2108 1452 4 ON2a
port 2 nsew
rlabel pwell s 1370 1334 1460 1460 4 ON1a
port 3 nsew
rlabel metal1 s 1720 -1526 1794 -1482 4 Gnd
port 4 nsew
rlabel metal2 s 1720 -1144 1792 -1080 4 vbiasn
port 5 nsew
<< end >>
