magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect -2760 4240 11100 4600
<< pwell >>
rect -2720 -3840 10560 -3680
<< psubdiff >>
rect -2720 -3709 10560 -3680
rect -2720 -3743 -1603 -3709
rect -2720 -3777 -2650 -3743
rect -2616 -3777 -2582 -3743
rect -2548 -3777 -2514 -3743
rect -2480 -3777 -2446 -3743
rect -2412 -3777 -2378 -3743
rect -2344 -3777 -2310 -3743
rect -2276 -3777 -2242 -3743
rect -2208 -3777 -2174 -3743
rect -2140 -3777 -2106 -3743
rect -2072 -3777 -2038 -3743
rect -2004 -3777 -1970 -3743
rect -1936 -3777 -1902 -3743
rect -1868 -3777 -1834 -3743
rect -1800 -3777 -1766 -3743
rect -1732 -3777 -1698 -3743
rect -1664 -3777 -1603 -3743
rect -2720 -3811 -1603 -3777
rect 2783 -3743 10560 -3709
rect 2783 -3777 2852 -3743
rect 2886 -3777 2920 -3743
rect 2954 -3777 2988 -3743
rect 3022 -3777 3056 -3743
rect 3090 -3777 3124 -3743
rect 3158 -3777 3192 -3743
rect 3226 -3777 3260 -3743
rect 3294 -3777 3328 -3743
rect 3362 -3777 3396 -3743
rect 3430 -3777 3464 -3743
rect 3498 -3777 3532 -3743
rect 3566 -3777 3600 -3743
rect 3634 -3777 3668 -3743
rect 3702 -3777 3736 -3743
rect 3770 -3777 3804 -3743
rect 3838 -3777 3872 -3743
rect 3906 -3777 3940 -3743
rect 3974 -3777 4008 -3743
rect 4042 -3777 4076 -3743
rect 4110 -3777 4144 -3743
rect 4178 -3777 4212 -3743
rect 4246 -3777 4280 -3743
rect 4314 -3777 4348 -3743
rect 4382 -3777 4416 -3743
rect 4450 -3777 4484 -3743
rect 4518 -3777 4552 -3743
rect 4586 -3777 4620 -3743
rect 4654 -3777 4688 -3743
rect 4722 -3777 4756 -3743
rect 4790 -3777 4824 -3743
rect 4858 -3777 4892 -3743
rect 4926 -3777 4960 -3743
rect 4994 -3777 5028 -3743
rect 5062 -3777 5096 -3743
rect 5130 -3777 5164 -3743
rect 5198 -3777 5232 -3743
rect 5266 -3777 5300 -3743
rect 5334 -3777 5368 -3743
rect 5402 -3777 5436 -3743
rect 5470 -3777 5504 -3743
rect 5538 -3777 5572 -3743
rect 5606 -3777 5640 -3743
rect 5674 -3777 5708 -3743
rect 5742 -3777 5776 -3743
rect 5810 -3777 5844 -3743
rect 5878 -3777 5912 -3743
rect 5946 -3777 5980 -3743
rect 6014 -3777 6048 -3743
rect 6082 -3777 6116 -3743
rect 6150 -3777 6184 -3743
rect 6218 -3777 6252 -3743
rect 6286 -3777 6320 -3743
rect 6354 -3777 6388 -3743
rect 6422 -3777 6456 -3743
rect 6490 -3777 6524 -3743
rect 6558 -3777 6592 -3743
rect 6626 -3777 6660 -3743
rect 6694 -3777 6728 -3743
rect 6762 -3777 6796 -3743
rect 6830 -3777 6864 -3743
rect 6898 -3777 6932 -3743
rect 6966 -3777 7000 -3743
rect 7034 -3777 7068 -3743
rect 7102 -3777 7136 -3743
rect 7170 -3777 7204 -3743
rect 7238 -3777 7272 -3743
rect 7306 -3777 7340 -3743
rect 7374 -3777 7408 -3743
rect 7442 -3777 7476 -3743
rect 7510 -3777 7544 -3743
rect 7578 -3777 7612 -3743
rect 7646 -3777 7680 -3743
rect 7714 -3777 7748 -3743
rect 7782 -3777 7816 -3743
rect 7850 -3777 7884 -3743
rect 7918 -3777 7952 -3743
rect 7986 -3777 8020 -3743
rect 8054 -3777 8088 -3743
rect 8122 -3777 8156 -3743
rect 8190 -3777 8224 -3743
rect 8258 -3777 8292 -3743
rect 8326 -3777 8360 -3743
rect 8394 -3777 8428 -3743
rect 8462 -3777 8496 -3743
rect 8530 -3777 8564 -3743
rect 8598 -3777 8632 -3743
rect 8666 -3777 8700 -3743
rect 8734 -3777 8768 -3743
rect 8802 -3777 8836 -3743
rect 8870 -3777 8904 -3743
rect 8938 -3777 8972 -3743
rect 9006 -3777 9040 -3743
rect 9074 -3777 9108 -3743
rect 9142 -3777 9176 -3743
rect 9210 -3777 9244 -3743
rect 9278 -3777 9312 -3743
rect 9346 -3777 9380 -3743
rect 9414 -3777 9448 -3743
rect 9482 -3777 9516 -3743
rect 9550 -3777 9584 -3743
rect 9618 -3777 9652 -3743
rect 9686 -3777 9720 -3743
rect 9754 -3777 9788 -3743
rect 9822 -3777 9856 -3743
rect 9890 -3777 9924 -3743
rect 9958 -3777 9992 -3743
rect 10026 -3777 10060 -3743
rect 10094 -3777 10128 -3743
rect 10162 -3777 10196 -3743
rect 10230 -3777 10264 -3743
rect 10298 -3777 10332 -3743
rect 10366 -3777 10400 -3743
rect 10434 -3777 10468 -3743
rect 10502 -3777 10560 -3743
rect 2783 -3811 10560 -3777
rect -2720 -3840 10560 -3811
<< nsubdiff >>
rect -2620 4437 10980 4480
rect -2620 4403 -2579 4437
rect -2545 4403 -2511 4437
rect -2477 4403 -2443 4437
rect -2409 4403 -2375 4437
rect -2341 4403 -2307 4437
rect -2273 4403 -2239 4437
rect -2205 4403 -2171 4437
rect -2137 4403 -2103 4437
rect -2069 4403 -2035 4437
rect -2001 4403 -1967 4437
rect -1933 4403 -1899 4437
rect -1865 4403 -1831 4437
rect -1797 4403 -1763 4437
rect -1729 4403 -1695 4437
rect -1661 4403 -1627 4437
rect -1593 4403 -1559 4437
rect -1525 4403 -1491 4437
rect -1457 4403 -1423 4437
rect -1389 4403 -1355 4437
rect -1321 4403 -1287 4437
rect -1253 4403 -1219 4437
rect -1185 4403 -1151 4437
rect -1117 4403 -1083 4437
rect -1049 4403 -1015 4437
rect -981 4403 -947 4437
rect -913 4403 -879 4437
rect -845 4403 -811 4437
rect -777 4403 -743 4437
rect -709 4403 -675 4437
rect -641 4403 -607 4437
rect -573 4403 -539 4437
rect -505 4403 -471 4437
rect -437 4403 -403 4437
rect -369 4403 -335 4437
rect -301 4403 -267 4437
rect -233 4403 -199 4437
rect -165 4403 -131 4437
rect -97 4403 -63 4437
rect -29 4403 5 4437
rect 39 4403 73 4437
rect 107 4403 141 4437
rect 175 4403 209 4437
rect 243 4403 277 4437
rect 311 4403 345 4437
rect 379 4403 413 4437
rect 447 4403 481 4437
rect 515 4403 549 4437
rect 583 4403 617 4437
rect 651 4403 685 4437
rect 719 4403 753 4437
rect 787 4403 821 4437
rect 855 4403 889 4437
rect 923 4403 957 4437
rect 991 4403 1025 4437
rect 1059 4403 1093 4437
rect 1127 4403 1161 4437
rect 1195 4403 1229 4437
rect 1263 4403 1297 4437
rect 1331 4403 1365 4437
rect 1399 4403 1433 4437
rect 1467 4403 1501 4437
rect 1535 4403 1569 4437
rect 1603 4403 1637 4437
rect 1671 4403 1705 4437
rect 1739 4403 1773 4437
rect 1807 4403 1841 4437
rect 1875 4403 1909 4437
rect 1943 4403 1977 4437
rect 2011 4403 2045 4437
rect 2079 4403 2113 4437
rect 2147 4403 2181 4437
rect 2215 4403 2249 4437
rect 2283 4403 2317 4437
rect 2351 4403 2385 4437
rect 2419 4403 2453 4437
rect 2487 4403 2521 4437
rect 2555 4403 2589 4437
rect 2623 4403 2657 4437
rect 2691 4403 2725 4437
rect 2759 4403 2793 4437
rect 2827 4403 2861 4437
rect 2895 4403 2929 4437
rect 2963 4403 2997 4437
rect 3031 4403 3065 4437
rect 3099 4403 3133 4437
rect 3167 4403 3201 4437
rect 3235 4403 3269 4437
rect 3303 4403 3337 4437
rect 3371 4403 3405 4437
rect 3439 4403 3473 4437
rect 3507 4403 3541 4437
rect 3575 4403 3609 4437
rect 3643 4403 3677 4437
rect 3711 4403 3745 4437
rect 3779 4403 3813 4437
rect 3847 4403 3881 4437
rect 3915 4403 3949 4437
rect 3983 4403 4017 4437
rect 4051 4403 4085 4437
rect 4119 4403 4153 4437
rect 4187 4403 4221 4437
rect 4255 4403 4289 4437
rect 4323 4403 4357 4437
rect 4391 4403 4425 4437
rect 4459 4403 4493 4437
rect 4527 4403 4561 4437
rect 4595 4403 4629 4437
rect 4663 4403 4697 4437
rect 4731 4403 4765 4437
rect 4799 4403 4833 4437
rect 4867 4403 4901 4437
rect 4935 4403 4969 4437
rect 5003 4403 5037 4437
rect 5071 4403 5105 4437
rect 5139 4403 5173 4437
rect 5207 4403 5241 4437
rect 5275 4403 5309 4437
rect 5343 4403 5377 4437
rect 5411 4403 5445 4437
rect 5479 4403 5513 4437
rect 5547 4403 5581 4437
rect 5615 4403 5649 4437
rect 5683 4403 5717 4437
rect 5751 4403 5785 4437
rect 5819 4403 5853 4437
rect 5887 4403 5921 4437
rect 5955 4403 5989 4437
rect 6023 4403 6057 4437
rect 6091 4403 6125 4437
rect 6159 4403 6193 4437
rect 6227 4403 6261 4437
rect 6295 4403 6329 4437
rect 6363 4403 6397 4437
rect 6431 4403 6465 4437
rect 6499 4403 6533 4437
rect 6567 4403 6601 4437
rect 6635 4403 6669 4437
rect 6703 4403 6737 4437
rect 6771 4403 6805 4437
rect 6839 4403 6873 4437
rect 6907 4403 6941 4437
rect 6975 4403 7009 4437
rect 7043 4403 7077 4437
rect 7111 4403 7145 4437
rect 7179 4403 7213 4437
rect 7247 4403 7281 4437
rect 7315 4403 7349 4437
rect 7383 4403 7417 4437
rect 7451 4403 7485 4437
rect 7519 4403 7553 4437
rect 7587 4403 7621 4437
rect 7655 4403 7689 4437
rect 7723 4403 7757 4437
rect 7791 4403 7825 4437
rect 7859 4403 7893 4437
rect 7927 4403 7961 4437
rect 7995 4403 8029 4437
rect 8063 4403 8097 4437
rect 8131 4403 8165 4437
rect 8199 4403 8233 4437
rect 8267 4403 8301 4437
rect 8335 4403 8369 4437
rect 8403 4403 8437 4437
rect 8471 4403 8505 4437
rect 8539 4403 8573 4437
rect 8607 4403 8641 4437
rect 8675 4403 8709 4437
rect 8743 4403 8777 4437
rect 8811 4403 8845 4437
rect 8879 4403 8913 4437
rect 8947 4403 8981 4437
rect 9015 4403 9049 4437
rect 9083 4403 9117 4437
rect 9151 4403 9185 4437
rect 9219 4403 9253 4437
rect 9287 4403 9321 4437
rect 9355 4403 9389 4437
rect 9423 4403 9457 4437
rect 9491 4403 9525 4437
rect 9559 4403 9593 4437
rect 9627 4403 9661 4437
rect 9695 4403 9729 4437
rect 9763 4403 9797 4437
rect 9831 4403 9865 4437
rect 9899 4403 9933 4437
rect 9967 4403 10001 4437
rect 10035 4403 10069 4437
rect 10103 4403 10137 4437
rect 10171 4403 10205 4437
rect 10239 4403 10273 4437
rect 10307 4403 10341 4437
rect 10375 4403 10409 4437
rect 10443 4403 10477 4437
rect 10511 4403 10545 4437
rect 10579 4403 10613 4437
rect 10647 4403 10681 4437
rect 10715 4403 10749 4437
rect 10783 4403 10817 4437
rect 10851 4403 10885 4437
rect 10919 4403 10980 4437
rect -2620 4360 10980 4403
<< psubdiffcont >>
rect -2650 -3777 -2616 -3743
rect -2582 -3777 -2548 -3743
rect -2514 -3777 -2480 -3743
rect -2446 -3777 -2412 -3743
rect -2378 -3777 -2344 -3743
rect -2310 -3777 -2276 -3743
rect -2242 -3777 -2208 -3743
rect -2174 -3777 -2140 -3743
rect -2106 -3777 -2072 -3743
rect -2038 -3777 -2004 -3743
rect -1970 -3777 -1936 -3743
rect -1902 -3777 -1868 -3743
rect -1834 -3777 -1800 -3743
rect -1766 -3777 -1732 -3743
rect -1698 -3777 -1664 -3743
rect -1603 -3811 2783 -3709
rect 2852 -3777 2886 -3743
rect 2920 -3777 2954 -3743
rect 2988 -3777 3022 -3743
rect 3056 -3777 3090 -3743
rect 3124 -3777 3158 -3743
rect 3192 -3777 3226 -3743
rect 3260 -3777 3294 -3743
rect 3328 -3777 3362 -3743
rect 3396 -3777 3430 -3743
rect 3464 -3777 3498 -3743
rect 3532 -3777 3566 -3743
rect 3600 -3777 3634 -3743
rect 3668 -3777 3702 -3743
rect 3736 -3777 3770 -3743
rect 3804 -3777 3838 -3743
rect 3872 -3777 3906 -3743
rect 3940 -3777 3974 -3743
rect 4008 -3777 4042 -3743
rect 4076 -3777 4110 -3743
rect 4144 -3777 4178 -3743
rect 4212 -3777 4246 -3743
rect 4280 -3777 4314 -3743
rect 4348 -3777 4382 -3743
rect 4416 -3777 4450 -3743
rect 4484 -3777 4518 -3743
rect 4552 -3777 4586 -3743
rect 4620 -3777 4654 -3743
rect 4688 -3777 4722 -3743
rect 4756 -3777 4790 -3743
rect 4824 -3777 4858 -3743
rect 4892 -3777 4926 -3743
rect 4960 -3777 4994 -3743
rect 5028 -3777 5062 -3743
rect 5096 -3777 5130 -3743
rect 5164 -3777 5198 -3743
rect 5232 -3777 5266 -3743
rect 5300 -3777 5334 -3743
rect 5368 -3777 5402 -3743
rect 5436 -3777 5470 -3743
rect 5504 -3777 5538 -3743
rect 5572 -3777 5606 -3743
rect 5640 -3777 5674 -3743
rect 5708 -3777 5742 -3743
rect 5776 -3777 5810 -3743
rect 5844 -3777 5878 -3743
rect 5912 -3777 5946 -3743
rect 5980 -3777 6014 -3743
rect 6048 -3777 6082 -3743
rect 6116 -3777 6150 -3743
rect 6184 -3777 6218 -3743
rect 6252 -3777 6286 -3743
rect 6320 -3777 6354 -3743
rect 6388 -3777 6422 -3743
rect 6456 -3777 6490 -3743
rect 6524 -3777 6558 -3743
rect 6592 -3777 6626 -3743
rect 6660 -3777 6694 -3743
rect 6728 -3777 6762 -3743
rect 6796 -3777 6830 -3743
rect 6864 -3777 6898 -3743
rect 6932 -3777 6966 -3743
rect 7000 -3777 7034 -3743
rect 7068 -3777 7102 -3743
rect 7136 -3777 7170 -3743
rect 7204 -3777 7238 -3743
rect 7272 -3777 7306 -3743
rect 7340 -3777 7374 -3743
rect 7408 -3777 7442 -3743
rect 7476 -3777 7510 -3743
rect 7544 -3777 7578 -3743
rect 7612 -3777 7646 -3743
rect 7680 -3777 7714 -3743
rect 7748 -3777 7782 -3743
rect 7816 -3777 7850 -3743
rect 7884 -3777 7918 -3743
rect 7952 -3777 7986 -3743
rect 8020 -3777 8054 -3743
rect 8088 -3777 8122 -3743
rect 8156 -3777 8190 -3743
rect 8224 -3777 8258 -3743
rect 8292 -3777 8326 -3743
rect 8360 -3777 8394 -3743
rect 8428 -3777 8462 -3743
rect 8496 -3777 8530 -3743
rect 8564 -3777 8598 -3743
rect 8632 -3777 8666 -3743
rect 8700 -3777 8734 -3743
rect 8768 -3777 8802 -3743
rect 8836 -3777 8870 -3743
rect 8904 -3777 8938 -3743
rect 8972 -3777 9006 -3743
rect 9040 -3777 9074 -3743
rect 9108 -3777 9142 -3743
rect 9176 -3777 9210 -3743
rect 9244 -3777 9278 -3743
rect 9312 -3777 9346 -3743
rect 9380 -3777 9414 -3743
rect 9448 -3777 9482 -3743
rect 9516 -3777 9550 -3743
rect 9584 -3777 9618 -3743
rect 9652 -3777 9686 -3743
rect 9720 -3777 9754 -3743
rect 9788 -3777 9822 -3743
rect 9856 -3777 9890 -3743
rect 9924 -3777 9958 -3743
rect 9992 -3777 10026 -3743
rect 10060 -3777 10094 -3743
rect 10128 -3777 10162 -3743
rect 10196 -3777 10230 -3743
rect 10264 -3777 10298 -3743
rect 10332 -3777 10366 -3743
rect 10400 -3777 10434 -3743
rect 10468 -3777 10502 -3743
<< nsubdiffcont >>
rect -2579 4403 -2545 4437
rect -2511 4403 -2477 4437
rect -2443 4403 -2409 4437
rect -2375 4403 -2341 4437
rect -2307 4403 -2273 4437
rect -2239 4403 -2205 4437
rect -2171 4403 -2137 4437
rect -2103 4403 -2069 4437
rect -2035 4403 -2001 4437
rect -1967 4403 -1933 4437
rect -1899 4403 -1865 4437
rect -1831 4403 -1797 4437
rect -1763 4403 -1729 4437
rect -1695 4403 -1661 4437
rect -1627 4403 -1593 4437
rect -1559 4403 -1525 4437
rect -1491 4403 -1457 4437
rect -1423 4403 -1389 4437
rect -1355 4403 -1321 4437
rect -1287 4403 -1253 4437
rect -1219 4403 -1185 4437
rect -1151 4403 -1117 4437
rect -1083 4403 -1049 4437
rect -1015 4403 -981 4437
rect -947 4403 -913 4437
rect -879 4403 -845 4437
rect -811 4403 -777 4437
rect -743 4403 -709 4437
rect -675 4403 -641 4437
rect -607 4403 -573 4437
rect -539 4403 -505 4437
rect -471 4403 -437 4437
rect -403 4403 -369 4437
rect -335 4403 -301 4437
rect -267 4403 -233 4437
rect -199 4403 -165 4437
rect -131 4403 -97 4437
rect -63 4403 -29 4437
rect 5 4403 39 4437
rect 73 4403 107 4437
rect 141 4403 175 4437
rect 209 4403 243 4437
rect 277 4403 311 4437
rect 345 4403 379 4437
rect 413 4403 447 4437
rect 481 4403 515 4437
rect 549 4403 583 4437
rect 617 4403 651 4437
rect 685 4403 719 4437
rect 753 4403 787 4437
rect 821 4403 855 4437
rect 889 4403 923 4437
rect 957 4403 991 4437
rect 1025 4403 1059 4437
rect 1093 4403 1127 4437
rect 1161 4403 1195 4437
rect 1229 4403 1263 4437
rect 1297 4403 1331 4437
rect 1365 4403 1399 4437
rect 1433 4403 1467 4437
rect 1501 4403 1535 4437
rect 1569 4403 1603 4437
rect 1637 4403 1671 4437
rect 1705 4403 1739 4437
rect 1773 4403 1807 4437
rect 1841 4403 1875 4437
rect 1909 4403 1943 4437
rect 1977 4403 2011 4437
rect 2045 4403 2079 4437
rect 2113 4403 2147 4437
rect 2181 4403 2215 4437
rect 2249 4403 2283 4437
rect 2317 4403 2351 4437
rect 2385 4403 2419 4437
rect 2453 4403 2487 4437
rect 2521 4403 2555 4437
rect 2589 4403 2623 4437
rect 2657 4403 2691 4437
rect 2725 4403 2759 4437
rect 2793 4403 2827 4437
rect 2861 4403 2895 4437
rect 2929 4403 2963 4437
rect 2997 4403 3031 4437
rect 3065 4403 3099 4437
rect 3133 4403 3167 4437
rect 3201 4403 3235 4437
rect 3269 4403 3303 4437
rect 3337 4403 3371 4437
rect 3405 4403 3439 4437
rect 3473 4403 3507 4437
rect 3541 4403 3575 4437
rect 3609 4403 3643 4437
rect 3677 4403 3711 4437
rect 3745 4403 3779 4437
rect 3813 4403 3847 4437
rect 3881 4403 3915 4437
rect 3949 4403 3983 4437
rect 4017 4403 4051 4437
rect 4085 4403 4119 4437
rect 4153 4403 4187 4437
rect 4221 4403 4255 4437
rect 4289 4403 4323 4437
rect 4357 4403 4391 4437
rect 4425 4403 4459 4437
rect 4493 4403 4527 4437
rect 4561 4403 4595 4437
rect 4629 4403 4663 4437
rect 4697 4403 4731 4437
rect 4765 4403 4799 4437
rect 4833 4403 4867 4437
rect 4901 4403 4935 4437
rect 4969 4403 5003 4437
rect 5037 4403 5071 4437
rect 5105 4403 5139 4437
rect 5173 4403 5207 4437
rect 5241 4403 5275 4437
rect 5309 4403 5343 4437
rect 5377 4403 5411 4437
rect 5445 4403 5479 4437
rect 5513 4403 5547 4437
rect 5581 4403 5615 4437
rect 5649 4403 5683 4437
rect 5717 4403 5751 4437
rect 5785 4403 5819 4437
rect 5853 4403 5887 4437
rect 5921 4403 5955 4437
rect 5989 4403 6023 4437
rect 6057 4403 6091 4437
rect 6125 4403 6159 4437
rect 6193 4403 6227 4437
rect 6261 4403 6295 4437
rect 6329 4403 6363 4437
rect 6397 4403 6431 4437
rect 6465 4403 6499 4437
rect 6533 4403 6567 4437
rect 6601 4403 6635 4437
rect 6669 4403 6703 4437
rect 6737 4403 6771 4437
rect 6805 4403 6839 4437
rect 6873 4403 6907 4437
rect 6941 4403 6975 4437
rect 7009 4403 7043 4437
rect 7077 4403 7111 4437
rect 7145 4403 7179 4437
rect 7213 4403 7247 4437
rect 7281 4403 7315 4437
rect 7349 4403 7383 4437
rect 7417 4403 7451 4437
rect 7485 4403 7519 4437
rect 7553 4403 7587 4437
rect 7621 4403 7655 4437
rect 7689 4403 7723 4437
rect 7757 4403 7791 4437
rect 7825 4403 7859 4437
rect 7893 4403 7927 4437
rect 7961 4403 7995 4437
rect 8029 4403 8063 4437
rect 8097 4403 8131 4437
rect 8165 4403 8199 4437
rect 8233 4403 8267 4437
rect 8301 4403 8335 4437
rect 8369 4403 8403 4437
rect 8437 4403 8471 4437
rect 8505 4403 8539 4437
rect 8573 4403 8607 4437
rect 8641 4403 8675 4437
rect 8709 4403 8743 4437
rect 8777 4403 8811 4437
rect 8845 4403 8879 4437
rect 8913 4403 8947 4437
rect 8981 4403 9015 4437
rect 9049 4403 9083 4437
rect 9117 4403 9151 4437
rect 9185 4403 9219 4437
rect 9253 4403 9287 4437
rect 9321 4403 9355 4437
rect 9389 4403 9423 4437
rect 9457 4403 9491 4437
rect 9525 4403 9559 4437
rect 9593 4403 9627 4437
rect 9661 4403 9695 4437
rect 9729 4403 9763 4437
rect 9797 4403 9831 4437
rect 9865 4403 9899 4437
rect 9933 4403 9967 4437
rect 10001 4403 10035 4437
rect 10069 4403 10103 4437
rect 10137 4403 10171 4437
rect 10205 4403 10239 4437
rect 10273 4403 10307 4437
rect 10341 4403 10375 4437
rect 10409 4403 10443 4437
rect 10477 4403 10511 4437
rect 10545 4403 10579 4437
rect 10613 4403 10647 4437
rect 10681 4403 10715 4437
rect 10749 4403 10783 4437
rect 10817 4403 10851 4437
rect 10885 4403 10919 4437
<< locali >>
rect -2620 4480 781 4488
rect -2620 4437 10980 4480
rect -2620 4403 -2579 4437
rect -2545 4403 -2511 4437
rect -2473 4403 -2443 4437
rect -2401 4403 -2375 4437
rect -2329 4403 -2307 4437
rect -2257 4403 -2239 4437
rect -2185 4403 -2171 4437
rect -2113 4403 -2103 4437
rect -2041 4403 -2035 4437
rect -1969 4403 -1967 4437
rect -1933 4403 -1931 4437
rect -1865 4403 -1859 4437
rect -1797 4403 -1787 4437
rect -1729 4403 -1715 4437
rect -1661 4403 -1643 4437
rect -1593 4403 -1571 4437
rect -1525 4403 -1499 4437
rect -1457 4403 -1427 4437
rect -1389 4403 -1355 4437
rect -1321 4403 -1287 4437
rect -1249 4403 -1219 4437
rect -1177 4403 -1151 4437
rect -1105 4403 -1083 4437
rect -1033 4403 -1015 4437
rect -961 4403 -947 4437
rect -889 4403 -879 4437
rect -817 4403 -811 4437
rect -745 4403 -743 4437
rect -709 4403 -707 4437
rect -641 4403 -635 4437
rect -573 4403 -563 4437
rect -505 4403 -491 4437
rect -437 4403 -419 4437
rect -369 4403 -347 4437
rect -301 4403 -275 4437
rect -233 4403 -203 4437
rect -165 4403 -131 4437
rect -97 4403 -63 4437
rect -25 4403 5 4437
rect 47 4403 73 4437
rect 119 4403 141 4437
rect 191 4403 209 4437
rect 263 4403 277 4437
rect 335 4403 345 4437
rect 407 4403 413 4437
rect 479 4403 481 4437
rect 515 4403 517 4437
rect 583 4403 589 4437
rect 651 4403 661 4437
rect 719 4403 733 4437
rect 787 4403 805 4437
rect 855 4403 877 4437
rect 923 4403 949 4437
rect 991 4403 1021 4437
rect 1059 4403 1093 4437
rect 1127 4403 1161 4437
rect 1199 4403 1229 4437
rect 1271 4403 1297 4437
rect 1343 4403 1365 4437
rect 1415 4403 1433 4437
rect 1487 4403 1501 4437
rect 1559 4403 1569 4437
rect 1631 4403 1637 4437
rect 1703 4403 1705 4437
rect 1739 4403 1741 4437
rect 1807 4403 1813 4437
rect 1875 4403 1885 4437
rect 1943 4403 1957 4437
rect 2011 4403 2029 4437
rect 2079 4403 2101 4437
rect 2147 4403 2173 4437
rect 2215 4403 2245 4437
rect 2283 4403 2317 4437
rect 2351 4403 2385 4437
rect 2423 4403 2453 4437
rect 2495 4403 2521 4437
rect 2567 4403 2589 4437
rect 2639 4403 2657 4437
rect 2711 4403 2725 4437
rect 2783 4403 2793 4437
rect 2855 4403 2861 4437
rect 2927 4403 2929 4437
rect 2963 4403 2965 4437
rect 3031 4403 3037 4437
rect 3099 4403 3109 4437
rect 3167 4403 3181 4437
rect 3235 4403 3253 4437
rect 3303 4403 3325 4437
rect 3371 4403 3397 4437
rect 3439 4403 3469 4437
rect 3507 4403 3541 4437
rect 3575 4403 3609 4437
rect 3647 4403 3677 4437
rect 3719 4403 3745 4437
rect 3791 4403 3813 4437
rect 3863 4403 3881 4437
rect 3935 4403 3949 4437
rect 4007 4403 4017 4437
rect 4079 4403 4085 4437
rect 4151 4403 4153 4437
rect 4187 4403 4189 4437
rect 4255 4403 4261 4437
rect 4323 4403 4333 4437
rect 4391 4403 4405 4437
rect 4459 4403 4477 4437
rect 4527 4403 4549 4437
rect 4595 4403 4621 4437
rect 4663 4403 4693 4437
rect 4731 4403 4765 4437
rect 4799 4403 4833 4437
rect 4871 4403 4901 4437
rect 4943 4403 4969 4437
rect 5015 4403 5037 4437
rect 5087 4403 5105 4437
rect 5159 4403 5173 4437
rect 5231 4403 5241 4437
rect 5303 4403 5309 4437
rect 5375 4403 5377 4437
rect 5411 4403 5413 4437
rect 5479 4403 5485 4437
rect 5547 4403 5557 4437
rect 5615 4403 5629 4437
rect 5683 4403 5701 4437
rect 5751 4403 5773 4437
rect 5819 4403 5845 4437
rect 5887 4403 5917 4437
rect 5955 4403 5989 4437
rect 6023 4403 6057 4437
rect 6095 4403 6125 4437
rect 6167 4403 6193 4437
rect 6239 4403 6261 4437
rect 6311 4403 6329 4437
rect 6383 4403 6397 4437
rect 6455 4403 6465 4437
rect 6527 4403 6533 4437
rect 6599 4403 6601 4437
rect 6635 4403 6637 4437
rect 6703 4403 6709 4437
rect 6771 4403 6781 4437
rect 6839 4403 6853 4437
rect 6907 4403 6925 4437
rect 6975 4403 6997 4437
rect 7043 4403 7069 4437
rect 7111 4403 7141 4437
rect 7179 4403 7213 4437
rect 7247 4403 7281 4437
rect 7319 4403 7349 4437
rect 7391 4403 7417 4437
rect 7463 4403 7485 4437
rect 7535 4403 7553 4437
rect 7607 4403 7621 4437
rect 7679 4403 7689 4437
rect 7751 4403 7757 4437
rect 7823 4403 7825 4437
rect 7859 4403 7861 4437
rect 7927 4403 7933 4437
rect 7995 4403 8005 4437
rect 8063 4403 8077 4437
rect 8131 4403 8149 4437
rect 8199 4403 8221 4437
rect 8267 4403 8293 4437
rect 8335 4403 8365 4437
rect 8403 4403 8437 4437
rect 8471 4403 8505 4437
rect 8543 4403 8573 4437
rect 8615 4403 8641 4437
rect 8687 4403 8709 4437
rect 8759 4403 8777 4437
rect 8831 4403 8845 4437
rect 8903 4403 8913 4437
rect 8975 4403 8981 4437
rect 9047 4403 9049 4437
rect 9083 4403 9085 4437
rect 9151 4403 9157 4437
rect 9219 4403 9229 4437
rect 9287 4403 9301 4437
rect 9355 4403 9373 4437
rect 9423 4403 9445 4437
rect 9491 4403 9517 4437
rect 9559 4403 9589 4437
rect 9627 4403 9661 4437
rect 9695 4403 9729 4437
rect 9767 4403 9797 4437
rect 9839 4403 9865 4437
rect 9911 4403 9933 4437
rect 9983 4403 10001 4437
rect 10055 4403 10069 4437
rect 10127 4403 10137 4437
rect 10199 4403 10205 4437
rect 10271 4403 10273 4437
rect 10307 4403 10309 4437
rect 10375 4403 10381 4437
rect 10443 4403 10453 4437
rect 10511 4403 10525 4437
rect 10579 4403 10597 4437
rect 10647 4403 10669 4437
rect 10715 4403 10741 4437
rect 10783 4403 10813 4437
rect 10851 4403 10885 4437
rect 10919 4403 10980 4437
rect -2620 4360 10980 4403
rect -2620 4197 781 4360
rect 2632 4213 6008 4360
rect 7681 4215 10942 4360
rect -2654 4195 781 4197
rect -2654 4194 -2620 4195
rect -2380 4137 -2280 4140
rect -2380 4103 -2347 4137
rect -2313 4103 -2280 4137
rect -2380 4100 -2280 4103
rect -1900 4137 -1800 4140
rect -1900 4103 -1867 4137
rect -1833 4103 -1800 4137
rect -1900 4100 -1800 4103
rect -1460 4137 -1360 4140
rect -1460 4103 -1427 4137
rect -1393 4103 -1360 4137
rect -1460 4100 -1360 4103
rect -1000 4137 -900 4140
rect -1000 4103 -967 4137
rect -933 4103 -900 4137
rect -1000 4100 -900 4103
rect -540 4137 -440 4140
rect -540 4103 -507 4137
rect -473 4103 -440 4137
rect -540 4100 -440 4103
rect -80 4137 20 4140
rect -80 4103 -47 4137
rect -13 4103 20 4137
rect -80 4100 20 4103
rect 380 4137 480 4140
rect 380 4103 413 4137
rect 447 4103 480 4137
rect 380 4100 480 4103
rect 2900 4137 3000 4140
rect 2900 4103 2933 4137
rect 2967 4103 3000 4137
rect 2900 4100 3000 4103
rect 3360 4137 3460 4140
rect 3360 4103 3393 4137
rect 3427 4103 3460 4137
rect 3360 4100 3460 4103
rect 3820 4137 3920 4140
rect 3820 4103 3853 4137
rect 3887 4103 3920 4137
rect 3820 4100 3920 4103
rect 4280 4137 4380 4140
rect 4280 4103 4313 4137
rect 4347 4103 4380 4137
rect 4280 4100 4380 4103
rect 4720 4137 4820 4140
rect 4720 4103 4753 4137
rect 4787 4103 4820 4137
rect 4720 4100 4820 4103
rect 5200 4137 5300 4140
rect 5200 4103 5233 4137
rect 5267 4103 5300 4137
rect 5200 4100 5300 4103
rect 5680 4137 5780 4140
rect 5680 4103 5713 4137
rect 5747 4103 5780 4137
rect 5680 4100 5780 4103
rect 7920 4137 8020 4140
rect 7920 4103 7953 4137
rect 7987 4103 8020 4137
rect 7920 4100 8020 4103
rect 8360 4137 8460 4140
rect 8360 4103 8393 4137
rect 8427 4103 8460 4137
rect 8360 4100 8460 4103
rect 8820 4137 8920 4140
rect 8820 4103 8853 4137
rect 8887 4103 8920 4137
rect 8820 4100 8920 4103
rect 9280 4137 9380 4140
rect 9280 4103 9313 4137
rect 9347 4103 9380 4137
rect 9280 4100 9380 4103
rect 9740 4137 9840 4140
rect 9740 4103 9773 4137
rect 9807 4103 9840 4137
rect 9740 4100 9840 4103
rect 10200 4137 10300 4140
rect 10200 4103 10233 4137
rect 10267 4103 10300 4137
rect 10200 4100 10300 4103
rect 10660 4137 10760 4140
rect 10660 4103 10693 4137
rect 10727 4103 10760 4137
rect 10660 4100 10760 4103
rect -2580 3753 -2540 3780
rect -2580 3719 -2577 3753
rect -2543 3719 -2540 3753
rect -2580 3681 -2540 3719
rect -2580 3647 -2577 3681
rect -2543 3647 -2540 3681
rect -2580 3620 -2540 3647
rect -1660 3753 -1620 3780
rect -1660 3719 -1657 3753
rect -1623 3719 -1620 3753
rect -1660 3681 -1620 3719
rect -1660 3647 -1657 3681
rect -1623 3647 -1620 3681
rect -1660 3620 -1620 3647
rect -740 3733 -700 3760
rect -740 3699 -737 3733
rect -703 3699 -700 3733
rect -740 3661 -700 3699
rect -740 3627 -737 3661
rect -703 3627 -700 3661
rect -740 3600 -700 3627
rect 160 3753 200 3780
rect 160 3719 163 3753
rect 197 3719 200 3753
rect 160 3681 200 3719
rect 160 3647 163 3681
rect 197 3647 200 3681
rect 160 3620 200 3647
rect 740 3743 780 3760
rect 740 3709 743 3743
rect 777 3709 780 3743
rect 740 3671 780 3709
rect 740 3637 743 3671
rect 777 3637 780 3671
rect 740 3620 780 3637
rect 2700 3733 2740 3760
rect 2700 3699 2703 3733
rect 2737 3699 2740 3733
rect 2700 3661 2740 3699
rect 2700 3627 2703 3661
rect 2737 3627 2740 3661
rect 2700 3600 2740 3627
rect 3620 3759 3660 3760
rect 3620 3725 3623 3759
rect 3657 3725 3660 3759
rect 3620 3687 3660 3725
rect 3620 3653 3623 3687
rect 3657 3653 3660 3687
rect 3620 3615 3660 3653
rect 3620 3581 3623 3615
rect 3657 3581 3660 3615
rect 3620 3580 3660 3581
rect 4540 3759 4580 3760
rect 4540 3725 4543 3759
rect 4577 3725 4580 3759
rect 4540 3687 4580 3725
rect 4540 3653 4543 3687
rect 4577 3653 4580 3687
rect 4540 3615 4580 3653
rect 4540 3581 4543 3615
rect 4577 3581 4580 3615
rect 4540 3580 4580 3581
rect 5460 3759 5500 3760
rect 5460 3725 5463 3759
rect 5497 3725 5500 3759
rect 5460 3687 5500 3725
rect 5460 3653 5463 3687
rect 5497 3653 5500 3687
rect 5460 3615 5500 3653
rect 6020 3743 6060 3760
rect 6020 3709 6023 3743
rect 6057 3709 6060 3743
rect 6020 3671 6060 3709
rect 6020 3637 6023 3671
rect 6057 3637 6060 3671
rect 6020 3620 6060 3637
rect 7600 3723 7640 3740
rect 7600 3689 7603 3723
rect 7637 3689 7640 3723
rect 7600 3651 7640 3689
rect 5460 3581 5463 3615
rect 5497 3581 5500 3615
rect 7600 3617 7603 3651
rect 7637 3617 7640 3651
rect 7600 3600 7640 3617
rect 7720 3713 7760 3720
rect 7720 3679 7723 3713
rect 7757 3679 7760 3713
rect 7720 3641 7760 3679
rect 7720 3607 7723 3641
rect 7757 3607 7760 3641
rect 7720 3600 7760 3607
rect 8640 3713 8680 3720
rect 8640 3679 8643 3713
rect 8677 3679 8680 3713
rect 8640 3641 8680 3679
rect 8640 3607 8643 3641
rect 8677 3607 8680 3641
rect 8640 3600 8680 3607
rect 9560 3713 9600 3720
rect 9560 3679 9563 3713
rect 9597 3679 9600 3713
rect 9560 3641 9600 3679
rect 9560 3607 9563 3641
rect 9597 3607 9600 3641
rect 9560 3600 9600 3607
rect 10480 3713 10520 3720
rect 10480 3679 10483 3713
rect 10517 3679 10520 3713
rect 10480 3641 10520 3679
rect 10480 3607 10483 3641
rect 10517 3607 10520 3641
rect 10480 3600 10520 3607
rect 5460 3580 5500 3581
rect -2100 3027 -2060 3060
rect -2100 2993 -2097 3027
rect -2063 2993 -2060 3027
rect -2100 2960 -2060 2993
rect -1200 3027 -1160 3060
rect -1200 2993 -1197 3027
rect -1163 2993 -1160 3027
rect -1200 2960 -1160 2993
rect -280 3027 -240 3060
rect -280 2993 -277 3027
rect -243 2993 -240 3027
rect -280 2960 -240 2993
rect 640 3027 680 3060
rect 640 2993 643 3027
rect 677 2993 680 3027
rect 640 2960 680 2993
rect 3160 3013 3200 3040
rect 3160 2979 3163 3013
rect 3197 2979 3200 3013
rect 3160 2941 3200 2979
rect 3160 2907 3163 2941
rect 3197 2907 3200 2941
rect 3160 2880 3200 2907
rect 4080 3013 4120 3040
rect 4080 2979 4083 3013
rect 4117 2979 4120 3013
rect 4080 2941 4120 2979
rect 4080 2907 4083 2941
rect 4117 2907 4120 2941
rect 4080 2880 4120 2907
rect 5000 3013 5040 3040
rect 5000 2979 5003 3013
rect 5037 2979 5040 3013
rect 5000 2941 5040 2979
rect 5000 2907 5003 2941
rect 5037 2907 5040 2941
rect 5000 2880 5040 2907
rect 5900 3013 5940 3040
rect 5900 2979 5903 3013
rect 5937 2979 5940 3013
rect 5900 2941 5940 2979
rect 5900 2907 5903 2941
rect 5937 2907 5940 2941
rect 5900 2880 5940 2907
rect 8160 2867 8200 2900
rect 8160 2833 8163 2867
rect 8197 2833 8200 2867
rect 8160 2800 8200 2833
rect 9080 2867 9120 2900
rect 9080 2833 9083 2867
rect 9117 2833 9120 2867
rect 9080 2800 9120 2833
rect 10000 2867 10040 2900
rect 10000 2833 10003 2867
rect 10037 2833 10040 2867
rect 10000 2800 10040 2833
rect 10900 2867 10940 2900
rect 10900 2833 10903 2867
rect 10937 2833 10940 2867
rect 10900 2800 10940 2833
rect -513 2607 -402 2614
rect -513 2573 -511 2607
rect -477 2573 -439 2607
rect -405 2573 -402 2607
rect -513 2566 -402 2573
rect -1300 2337 -1220 2340
rect -1300 2303 -1277 2337
rect -1243 2303 -1220 2337
rect -1300 2300 -1220 2303
rect 4020 2337 4140 2340
rect 4020 2303 4027 2337
rect 4061 2303 4099 2337
rect 4133 2303 4140 2337
rect 4020 2300 4140 2303
rect 6900 2297 6960 2320
rect 6900 2263 6913 2297
rect 6947 2263 6960 2297
rect 6900 2240 6960 2263
rect 1284 2135 1410 2139
rect 1284 2101 1294 2135
rect 1328 2101 1366 2135
rect 1400 2101 1410 2135
rect 1284 2097 1410 2101
rect 4040 2137 4160 2140
rect 4040 2103 4047 2137
rect 4081 2103 4119 2137
rect 4153 2103 4160 2137
rect 4040 2100 4160 2103
rect 6880 2137 7000 2140
rect 6880 2103 6887 2137
rect 6921 2103 6959 2137
rect 6993 2103 7000 2137
rect 6880 2100 7000 2103
rect 4040 2037 4140 2040
rect 1284 2014 1410 2018
rect 1284 1980 1294 2014
rect 1328 1980 1366 2014
rect 1400 1980 1410 2014
rect 4040 2003 4073 2037
rect 4107 2003 4140 2037
rect 4040 2000 4140 2003
rect 6880 2037 7020 2040
rect 6880 2003 6897 2037
rect 6931 2003 6969 2037
rect 7003 2003 7020 2037
rect 6880 2000 7020 2003
rect 1284 1976 1410 1980
rect 2301 1886 2345 1912
rect 2301 1852 2306 1886
rect 2340 1852 2345 1886
rect 2301 1827 2345 1852
rect 3360 1887 3400 1920
rect 3360 1853 3363 1887
rect 3397 1853 3400 1887
rect 3360 1820 3400 1853
rect 4671 1912 4735 1918
rect 4671 1878 4686 1912
rect 4720 1878 4735 1912
rect 4671 1840 4735 1878
rect 4671 1806 4686 1840
rect 4720 1806 4735 1840
rect 6160 1887 6200 1920
rect 6160 1853 6163 1887
rect 6197 1853 6200 1887
rect 6160 1820 6200 1853
rect 4671 1801 4735 1806
rect 3540 1757 3700 1760
rect 2043 1748 2169 1753
rect 2043 1714 2053 1748
rect 2087 1714 2125 1748
rect 2159 1714 2169 1748
rect 3540 1723 3567 1757
rect 3601 1723 3639 1757
rect 3673 1723 3700 1757
rect 3540 1720 3700 1723
rect 6880 1757 7020 1760
rect 6880 1723 6897 1757
rect 6931 1723 6969 1757
rect 7003 1723 7020 1757
rect 6880 1720 7020 1723
rect 2043 1710 2169 1714
rect 6880 1197 7020 1200
rect 2060 1165 2140 1180
rect 2060 1131 2083 1165
rect 2117 1131 2140 1165
rect 6880 1163 6897 1197
rect 6931 1163 6969 1197
rect 7003 1163 7020 1197
rect 6880 1160 7020 1163
rect 2060 1093 2140 1131
rect 2060 1059 2083 1093
rect 2117 1059 2140 1093
rect 2060 1021 2140 1059
rect 2060 987 2083 1021
rect 2117 987 2140 1021
rect 6140 1057 6180 1060
rect 6140 1023 6143 1057
rect 6177 1023 6180 1057
rect 6140 1020 6180 1023
rect 2060 949 2140 987
rect 2060 915 2083 949
rect 2117 915 2140 949
rect 2060 900 2140 915
rect 6580 937 6740 940
rect 6580 903 6607 937
rect 6641 903 6679 937
rect 6713 903 6740 937
rect 6580 900 6740 903
rect 7500 937 7660 940
rect 7500 903 7527 937
rect 7561 903 7599 937
rect 7633 903 7660 937
rect 7500 900 7660 903
rect 4940 857 5100 860
rect 1060 833 1100 840
rect 1060 799 1063 833
rect 1097 799 1100 833
rect 4940 823 4967 857
rect 5001 823 5039 857
rect 5073 823 5100 857
rect 4940 820 5100 823
rect 1060 761 1100 799
rect 6620 817 6700 820
rect 6620 783 6643 817
rect 6677 783 6700 817
rect 6620 780 6700 783
rect 1060 727 1063 761
rect 1097 727 1100 761
rect 1060 720 1100 727
rect 2872 720 2913 747
rect 2872 686 2875 720
rect 2909 686 2913 720
rect 2872 660 2913 686
rect 5380 717 5420 740
rect 5380 683 5383 717
rect 5417 683 5420 717
rect 5380 660 5420 683
rect 3700 577 3740 580
rect 3700 543 3703 577
rect 3737 543 3740 577
rect 3700 540 3740 543
rect 2060 471 2140 500
rect 2060 437 2083 471
rect 2117 437 2140 471
rect 3660 477 3760 480
rect 3660 443 3693 477
rect 3727 443 3760 477
rect 3660 440 3760 443
rect -1900 383 -1860 400
rect -1900 349 -1897 383
rect -1863 349 -1860 383
rect -1900 311 -1860 349
rect -1900 277 -1897 311
rect -1863 277 -1860 311
rect -1900 260 -1860 277
rect -1800 383 -1760 400
rect -1800 349 -1797 383
rect -1763 349 -1760 383
rect -1800 311 -1760 349
rect -1800 277 -1797 311
rect -1763 277 -1760 311
rect -1800 260 -1760 277
rect -1338 386 -1301 398
rect -1338 352 -1337 386
rect -1303 352 -1301 386
rect -1338 314 -1301 352
rect -1338 280 -1337 314
rect -1303 280 -1301 314
rect -1338 269 -1301 280
rect -20 363 20 380
rect -20 329 -17 363
rect 17 329 20 363
rect -20 291 20 329
rect -20 257 -17 291
rect 17 257 20 291
rect -20 240 20 257
rect 80 373 120 400
rect 2060 399 2140 437
rect 80 339 83 373
rect 117 339 120 373
rect 80 301 120 339
rect 80 267 83 301
rect 117 267 120 301
rect 80 240 120 267
rect 540 372 589 383
rect 540 338 547 372
rect 581 338 589 372
rect 540 300 589 338
rect 540 266 547 300
rect 581 266 589 300
rect 540 255 589 266
rect 2060 365 2083 399
rect 2117 365 2140 399
rect 2060 327 2140 365
rect 2060 293 2083 327
rect 2117 293 2140 327
rect 2060 255 2140 293
rect 2060 221 2083 255
rect 2117 221 2140 255
rect 2060 183 2140 221
rect 298 131 311 165
rect 345 131 358 165
rect 2060 149 2083 183
rect 2117 149 2140 183
rect 5740 217 5820 220
rect 5740 183 5763 217
rect 5797 183 5820 217
rect 5740 180 5820 183
rect 2060 120 2140 149
rect -1620 87 -1460 100
rect -1620 53 -1593 87
rect -1559 53 -1521 87
rect -1487 53 -1460 87
rect -1620 40 -1460 53
rect 4620 -577 4660 -560
rect 2780 -597 2820 -580
rect 2780 -631 2783 -597
rect 2817 -631 2820 -597
rect 2780 -669 2820 -631
rect 2780 -703 2783 -669
rect 2817 -703 2820 -669
rect 2780 -720 2820 -703
rect 3700 -597 3740 -580
rect 3700 -631 3703 -597
rect 3737 -631 3740 -597
rect 3700 -669 3740 -631
rect 3700 -703 3703 -669
rect 3737 -703 3740 -669
rect 4620 -611 4623 -577
rect 4657 -611 4660 -577
rect 4620 -649 4660 -611
rect 4620 -683 4623 -649
rect 4657 -683 4660 -649
rect 4620 -700 4660 -683
rect 5540 -577 5580 -560
rect 5540 -611 5543 -577
rect 5577 -611 5580 -577
rect 5540 -649 5580 -611
rect 5540 -683 5543 -649
rect 5577 -683 5580 -649
rect 5540 -700 5580 -683
rect 6640 -587 6680 -560
rect 6640 -621 6643 -587
rect 6677 -621 6680 -587
rect 6640 -659 6680 -621
rect 6640 -693 6643 -659
rect 6677 -693 6680 -659
rect 3700 -720 3740 -703
rect 6640 -720 6680 -693
rect 7560 -587 7600 -560
rect 7560 -621 7563 -587
rect 7597 -621 7600 -587
rect 7560 -659 7600 -621
rect 7560 -693 7563 -659
rect 7597 -693 7600 -659
rect 7560 -720 7600 -693
rect 8480 -567 8520 -540
rect 8480 -601 8483 -567
rect 8517 -601 8520 -567
rect 8480 -639 8520 -601
rect 8480 -673 8483 -639
rect 8517 -673 8520 -639
rect 8480 -700 8520 -673
rect 9400 -567 9440 -540
rect 9400 -601 9403 -567
rect 9437 -601 9440 -567
rect 9400 -639 9440 -601
rect 9400 -673 9403 -639
rect 9437 -673 9440 -639
rect 9400 -700 9440 -673
rect 3240 -1093 3280 -1060
rect 3240 -1127 3243 -1093
rect 3277 -1127 3280 -1093
rect 3240 -1160 3280 -1127
rect 4160 -1093 4200 -1060
rect 4160 -1127 4163 -1093
rect 4197 -1127 4200 -1093
rect 4160 -1160 4200 -1127
rect 5080 -1093 5120 -1060
rect 5080 -1127 5083 -1093
rect 5117 -1127 5120 -1093
rect 5080 -1160 5120 -1127
rect 6000 -1093 6040 -1060
rect 6000 -1127 6003 -1093
rect 6037 -1127 6040 -1093
rect 6000 -1160 6040 -1127
rect 6100 -1103 6140 -1080
rect 6100 -1137 6103 -1103
rect 6137 -1137 6140 -1103
rect 6100 -1160 6140 -1137
rect 7100 -1093 7140 -1060
rect 7100 -1127 7103 -1093
rect 7137 -1127 7140 -1093
rect 7100 -1160 7140 -1127
rect 8020 -1093 8060 -1060
rect 8020 -1127 8023 -1093
rect 8057 -1127 8060 -1093
rect 8020 -1160 8060 -1127
rect 8940 -1093 8980 -1060
rect 8940 -1127 8943 -1093
rect 8977 -1127 8980 -1093
rect 8940 -1160 8980 -1127
rect 9860 -1093 9900 -1060
rect 9860 -1127 9863 -1093
rect 9897 -1127 9900 -1093
rect 9860 -1160 9900 -1127
rect 9960 -1083 10000 -1060
rect 9960 -1117 9963 -1083
rect 9997 -1117 10000 -1083
rect 9960 -1140 10000 -1117
rect 2980 -1303 3100 -1300
rect 2980 -1337 2987 -1303
rect 3021 -1337 3059 -1303
rect 3093 -1337 3100 -1303
rect 2980 -1340 3100 -1337
rect 3460 -1303 3580 -1300
rect 3460 -1337 3467 -1303
rect 3501 -1337 3539 -1303
rect 3573 -1337 3580 -1303
rect 3460 -1340 3580 -1337
rect 3900 -1303 4020 -1300
rect 3900 -1337 3907 -1303
rect 3941 -1337 3979 -1303
rect 4013 -1337 4020 -1303
rect 3900 -1340 4020 -1337
rect 4360 -1303 4480 -1300
rect 4360 -1337 4367 -1303
rect 4401 -1337 4439 -1303
rect 4473 -1337 4480 -1303
rect 4360 -1340 4480 -1337
rect 4840 -1303 4960 -1300
rect 4840 -1337 4847 -1303
rect 4881 -1337 4919 -1303
rect 4953 -1337 4960 -1303
rect 4840 -1340 4960 -1337
rect 5280 -1303 5400 -1300
rect 5280 -1337 5287 -1303
rect 5321 -1337 5359 -1303
rect 5393 -1337 5400 -1303
rect 5280 -1340 5400 -1337
rect 5740 -1303 5860 -1300
rect 5740 -1337 5747 -1303
rect 5781 -1337 5819 -1303
rect 5853 -1337 5860 -1303
rect 5740 -1340 5860 -1337
rect 6840 -1303 6960 -1300
rect 6840 -1337 6847 -1303
rect 6881 -1337 6919 -1303
rect 6953 -1337 6960 -1303
rect 6840 -1340 6960 -1337
rect 7320 -1303 7440 -1300
rect 7320 -1337 7327 -1303
rect 7361 -1337 7399 -1303
rect 7433 -1337 7440 -1303
rect 7320 -1340 7440 -1337
rect 7760 -1303 7880 -1300
rect 7760 -1337 7767 -1303
rect 7801 -1337 7839 -1303
rect 7873 -1337 7880 -1303
rect 7760 -1340 7880 -1337
rect 8220 -1303 8340 -1300
rect 8220 -1337 8227 -1303
rect 8261 -1337 8299 -1303
rect 8333 -1337 8340 -1303
rect 8220 -1340 8340 -1337
rect 8680 -1303 8800 -1300
rect 8680 -1337 8687 -1303
rect 8721 -1337 8759 -1303
rect 8793 -1337 8800 -1303
rect 8680 -1340 8800 -1337
rect 9160 -1303 9280 -1300
rect 9160 -1337 9167 -1303
rect 9201 -1337 9239 -1303
rect 9273 -1337 9280 -1303
rect 9160 -1340 9280 -1337
rect 9620 -1303 9740 -1300
rect 9620 -1337 9627 -1303
rect 9661 -1337 9699 -1303
rect 9733 -1337 9740 -1303
rect 9620 -1340 9740 -1337
rect -1780 -2263 -1740 -2240
rect -1780 -2297 -1777 -2263
rect -1743 -2297 -1740 -2263
rect -1780 -2320 -1740 -2297
rect -860 -2263 -820 -2240
rect -860 -2297 -857 -2263
rect -823 -2297 -820 -2263
rect -860 -2320 -820 -2297
rect 60 -2263 100 -2240
rect 60 -2297 63 -2263
rect 97 -2297 100 -2263
rect 60 -2320 100 -2297
rect 980 -2263 1020 -2240
rect 980 -2297 983 -2263
rect 1017 -2297 1020 -2263
rect 980 -2320 1020 -2297
rect 1900 -2263 1940 -2240
rect 1900 -2297 1903 -2263
rect 1937 -2297 1940 -2263
rect 1900 -2320 1940 -2297
rect 2800 -2263 2840 -2240
rect 2800 -2297 2803 -2263
rect 2837 -2297 2840 -2263
rect 2800 -2320 2840 -2297
rect 4960 -2293 5000 -2260
rect 4960 -2327 4963 -2293
rect 4997 -2327 5000 -2293
rect 4960 -2360 5000 -2327
rect 5880 -2293 5920 -2260
rect 5880 -2327 5883 -2293
rect 5917 -2327 5920 -2293
rect 5880 -2360 5920 -2327
rect 6800 -2293 6840 -2260
rect 6800 -2327 6803 -2293
rect 6837 -2327 6840 -2293
rect 6800 -2360 6840 -2327
rect 7720 -2293 7760 -2260
rect 7720 -2327 7723 -2293
rect 7757 -2327 7760 -2293
rect 7720 -2360 7760 -2327
rect 8640 -2293 8680 -2260
rect 8640 -2327 8643 -2293
rect 8677 -2327 8680 -2293
rect 8640 -2360 8680 -2327
rect 9540 -2313 9580 -2280
rect 9540 -2347 9543 -2313
rect 9577 -2347 9580 -2313
rect 9540 -2380 9580 -2347
rect 10460 -2313 10500 -2280
rect 10460 -2347 10463 -2313
rect 10497 -2347 10500 -2313
rect 10460 -2380 10500 -2347
rect -2060 -3107 -2020 -3100
rect -2180 -3143 -2140 -3120
rect -2180 -3177 -2177 -3143
rect -2143 -3177 -2140 -3143
rect -2180 -3200 -2140 -3177
rect -2060 -3141 -2057 -3107
rect -2023 -3141 -2020 -3107
rect -2060 -3179 -2020 -3141
rect -2060 -3213 -2057 -3179
rect -2023 -3213 -2020 -3179
rect -2060 -3220 -2020 -3213
rect -1880 -3153 -1840 -3120
rect -1880 -3187 -1877 -3153
rect -1843 -3187 -1840 -3153
rect -1880 -3220 -1840 -3187
rect -1320 -3143 -1280 -3120
rect -1320 -3177 -1317 -3143
rect -1283 -3177 -1280 -3143
rect -1320 -3200 -1280 -3177
rect -400 -3143 -360 -3120
rect -400 -3177 -397 -3143
rect -363 -3177 -360 -3143
rect -400 -3200 -360 -3177
rect 520 -3143 560 -3120
rect 520 -3177 523 -3143
rect 557 -3177 560 -3143
rect 520 -3200 560 -3177
rect 1440 -3143 1480 -3120
rect 1440 -3177 1443 -3143
rect 1477 -3177 1480 -3143
rect 1440 -3200 1480 -3177
rect 2340 -3143 2380 -3120
rect 2340 -3177 2343 -3143
rect 2377 -3177 2380 -3143
rect 2340 -3200 2380 -3177
rect 3880 -3143 3940 -3140
rect 3880 -3177 3893 -3143
rect 3927 -3177 3940 -3143
rect 3880 -3180 3940 -3177
rect 4860 -3143 4900 -3120
rect 4860 -3177 4863 -3143
rect 4897 -3177 4900 -3143
rect 4860 -3200 4900 -3177
rect 5420 -3143 5460 -3120
rect 5420 -3177 5423 -3143
rect 5457 -3177 5460 -3143
rect 5420 -3200 5460 -3177
rect 6340 -3143 6380 -3120
rect 6340 -3177 6343 -3143
rect 6377 -3177 6380 -3143
rect 6340 -3200 6380 -3177
rect 7260 -3143 7300 -3120
rect 7260 -3177 7263 -3143
rect 7297 -3177 7300 -3143
rect 7260 -3200 7300 -3177
rect 8160 -3143 8200 -3120
rect 8160 -3177 8163 -3143
rect 8197 -3177 8200 -3143
rect 8160 -3200 8200 -3177
rect 9080 -3143 9120 -3120
rect 9080 -3177 9083 -3143
rect 9117 -3177 9120 -3143
rect 9080 -3200 9120 -3177
rect 10000 -3143 10040 -3120
rect 10000 -3177 10003 -3143
rect 10037 -3177 10040 -3143
rect 10000 -3200 10040 -3177
rect -2640 -3333 -2600 -3300
rect -2640 -3367 -2637 -3333
rect -2603 -3367 -2600 -3333
rect -2640 -3400 -2600 -3367
rect -2480 -3443 -2340 -3440
rect -2480 -3477 -2463 -3443
rect -2429 -3477 -2391 -3443
rect -2357 -3477 -2340 -3443
rect -2480 -3480 -2340 -3477
rect -1600 -3443 -1460 -3440
rect -1600 -3477 -1583 -3443
rect -1549 -3477 -1511 -3443
rect -1477 -3477 -1460 -3443
rect -1600 -3480 -1460 -3477
rect -1140 -3443 -1000 -3440
rect -1140 -3477 -1123 -3443
rect -1089 -3477 -1051 -3443
rect -1017 -3477 -1000 -3443
rect -1140 -3480 -1000 -3477
rect -680 -3443 -540 -3440
rect -680 -3477 -663 -3443
rect -629 -3477 -591 -3443
rect -557 -3477 -540 -3443
rect -680 -3480 -540 -3477
rect -260 -3443 -120 -3440
rect -260 -3477 -243 -3443
rect -209 -3477 -171 -3443
rect -137 -3477 -120 -3443
rect -260 -3480 -120 -3477
rect 220 -3443 360 -3440
rect 220 -3477 237 -3443
rect 271 -3477 309 -3443
rect 343 -3477 360 -3443
rect 220 -3480 360 -3477
rect 680 -3443 820 -3440
rect 680 -3477 697 -3443
rect 731 -3477 769 -3443
rect 803 -3477 820 -3443
rect 680 -3480 820 -3477
rect 1140 -3443 1280 -3440
rect 1140 -3477 1157 -3443
rect 1191 -3477 1229 -3443
rect 1263 -3477 1280 -3443
rect 1140 -3480 1280 -3477
rect 1600 -3443 1740 -3440
rect 1600 -3477 1617 -3443
rect 1651 -3477 1689 -3443
rect 1723 -3477 1740 -3443
rect 1600 -3480 1740 -3477
rect 2060 -3443 2200 -3440
rect 2060 -3477 2077 -3443
rect 2111 -3477 2149 -3443
rect 2183 -3477 2200 -3443
rect 2060 -3480 2200 -3477
rect 2540 -3443 2680 -3440
rect 2540 -3477 2557 -3443
rect 2591 -3477 2629 -3443
rect 2663 -3477 2680 -3443
rect 2540 -3480 2680 -3477
rect 5160 -3443 5280 -3440
rect 5160 -3477 5167 -3443
rect 5201 -3477 5239 -3443
rect 5273 -3477 5280 -3443
rect 5160 -3480 5280 -3477
rect 5620 -3443 5740 -3440
rect 5620 -3477 5627 -3443
rect 5661 -3477 5699 -3443
rect 5733 -3477 5740 -3443
rect 5620 -3480 5740 -3477
rect 6080 -3443 6200 -3440
rect 6080 -3477 6087 -3443
rect 6121 -3477 6159 -3443
rect 6193 -3477 6200 -3443
rect 6080 -3480 6200 -3477
rect 6540 -3443 6660 -3440
rect 6540 -3477 6547 -3443
rect 6581 -3477 6619 -3443
rect 6653 -3477 6660 -3443
rect 6540 -3480 6660 -3477
rect 7000 -3443 7120 -3440
rect 7000 -3477 7007 -3443
rect 7041 -3477 7079 -3443
rect 7113 -3477 7120 -3443
rect 7000 -3480 7120 -3477
rect 7440 -3443 7560 -3440
rect 7440 -3477 7447 -3443
rect 7481 -3477 7519 -3443
rect 7553 -3477 7560 -3443
rect 7440 -3480 7560 -3477
rect 7900 -3443 8020 -3440
rect 7900 -3477 7907 -3443
rect 7941 -3477 7979 -3443
rect 8013 -3477 8020 -3443
rect 7900 -3480 8020 -3477
rect 8360 -3443 8480 -3440
rect 8360 -3477 8367 -3443
rect 8401 -3477 8439 -3443
rect 8473 -3477 8480 -3443
rect 8360 -3480 8480 -3477
rect 8840 -3443 8960 -3440
rect 8840 -3477 8847 -3443
rect 8881 -3477 8919 -3443
rect 8953 -3477 8960 -3443
rect 8840 -3480 8960 -3477
rect 9280 -3443 9400 -3440
rect 9280 -3477 9287 -3443
rect 9321 -3477 9359 -3443
rect 9393 -3477 9400 -3443
rect 9280 -3480 9400 -3477
rect 9740 -3443 9860 -3440
rect 9740 -3477 9747 -3443
rect 9781 -3477 9819 -3443
rect 9853 -3477 9860 -3443
rect 9740 -3480 9860 -3477
rect 10200 -3443 10320 -3440
rect 10200 -3477 10207 -3443
rect 10241 -3477 10279 -3443
rect 10313 -3477 10320 -3443
rect 10200 -3480 10320 -3477
rect -2720 -3709 10560 -3680
rect -2720 -3743 -1603 -3709
rect 2783 -3743 10560 -3709
rect -2720 -3777 -2650 -3743
rect -2605 -3777 -2582 -3743
rect -2533 -3777 -2514 -3743
rect -2461 -3777 -2446 -3743
rect -2389 -3777 -2378 -3743
rect -2317 -3777 -2310 -3743
rect -2245 -3777 -2242 -3743
rect -2208 -3777 -2207 -3743
rect -2140 -3777 -2135 -3743
rect -2072 -3777 -2063 -3743
rect -2004 -3777 -1991 -3743
rect -1936 -3777 -1919 -3743
rect -1868 -3777 -1847 -3743
rect -1800 -3777 -1775 -3743
rect -1732 -3777 -1703 -3743
rect -1664 -3777 -1631 -3743
rect 2795 -3777 2833 -3743
rect 2886 -3777 2905 -3743
rect 2954 -3777 2977 -3743
rect 3022 -3777 3049 -3743
rect 3090 -3777 3121 -3743
rect 3158 -3777 3192 -3743
rect 3227 -3777 3260 -3743
rect 3299 -3777 3328 -3743
rect 3371 -3777 3396 -3743
rect 3443 -3777 3464 -3743
rect 3515 -3777 3532 -3743
rect 3587 -3777 3600 -3743
rect 3659 -3777 3668 -3743
rect 3731 -3777 3736 -3743
rect 3803 -3777 3804 -3743
rect 3838 -3777 3841 -3743
rect 3906 -3777 3913 -3743
rect 3974 -3777 3985 -3743
rect 4042 -3777 4057 -3743
rect 4110 -3777 4129 -3743
rect 4178 -3777 4201 -3743
rect 4246 -3777 4273 -3743
rect 4314 -3777 4345 -3743
rect 4382 -3777 4416 -3743
rect 4451 -3777 4484 -3743
rect 4523 -3777 4552 -3743
rect 4595 -3777 4620 -3743
rect 4667 -3777 4688 -3743
rect 4739 -3777 4756 -3743
rect 4811 -3777 4824 -3743
rect 4883 -3777 4892 -3743
rect 4955 -3777 4960 -3743
rect 5027 -3777 5028 -3743
rect 5062 -3777 5065 -3743
rect 5130 -3777 5137 -3743
rect 5198 -3777 5209 -3743
rect 5266 -3777 5281 -3743
rect 5334 -3777 5353 -3743
rect 5402 -3777 5425 -3743
rect 5470 -3777 5497 -3743
rect 5538 -3777 5569 -3743
rect 5606 -3777 5640 -3743
rect 5675 -3777 5708 -3743
rect 5747 -3777 5776 -3743
rect 5819 -3777 5844 -3743
rect 5891 -3777 5912 -3743
rect 5963 -3777 5980 -3743
rect 6035 -3777 6048 -3743
rect 6107 -3777 6116 -3743
rect 6179 -3777 6184 -3743
rect 6251 -3777 6252 -3743
rect 6286 -3777 6289 -3743
rect 6354 -3777 6361 -3743
rect 6422 -3777 6433 -3743
rect 6490 -3777 6505 -3743
rect 6558 -3777 6577 -3743
rect 6626 -3777 6649 -3743
rect 6694 -3777 6721 -3743
rect 6762 -3777 6793 -3743
rect 6830 -3777 6864 -3743
rect 6899 -3777 6932 -3743
rect 6971 -3777 7000 -3743
rect 7043 -3777 7068 -3743
rect 7115 -3777 7136 -3743
rect 7187 -3777 7204 -3743
rect 7259 -3777 7272 -3743
rect 7331 -3777 7340 -3743
rect 7403 -3777 7408 -3743
rect 7475 -3777 7476 -3743
rect 7510 -3777 7513 -3743
rect 7578 -3777 7585 -3743
rect 7646 -3777 7657 -3743
rect 7714 -3777 7729 -3743
rect 7782 -3777 7801 -3743
rect 7850 -3777 7873 -3743
rect 7918 -3777 7945 -3743
rect 7986 -3777 8017 -3743
rect 8054 -3777 8088 -3743
rect 8123 -3777 8156 -3743
rect 8195 -3777 8224 -3743
rect 8267 -3777 8292 -3743
rect 8339 -3777 8360 -3743
rect 8411 -3777 8428 -3743
rect 8483 -3777 8496 -3743
rect 8555 -3777 8564 -3743
rect 8627 -3777 8632 -3743
rect 8699 -3777 8700 -3743
rect 8734 -3777 8737 -3743
rect 8802 -3777 8809 -3743
rect 8870 -3777 8881 -3743
rect 8938 -3777 8953 -3743
rect 9006 -3777 9025 -3743
rect 9074 -3777 9097 -3743
rect 9142 -3777 9169 -3743
rect 9210 -3777 9241 -3743
rect 9278 -3777 9312 -3743
rect 9347 -3777 9380 -3743
rect 9419 -3777 9448 -3743
rect 9491 -3777 9516 -3743
rect 9563 -3777 9584 -3743
rect 9635 -3777 9652 -3743
rect 9707 -3777 9720 -3743
rect 9779 -3777 9788 -3743
rect 9851 -3777 9856 -3743
rect 9923 -3777 9924 -3743
rect 9958 -3777 9961 -3743
rect 10026 -3777 10033 -3743
rect 10094 -3777 10105 -3743
rect 10162 -3777 10177 -3743
rect 10230 -3777 10249 -3743
rect 10298 -3777 10321 -3743
rect 10366 -3777 10393 -3743
rect 10434 -3777 10465 -3743
rect 10502 -3777 10560 -3743
rect -2720 -3811 -1603 -3777
rect 2783 -3811 10560 -3777
rect -2720 -3840 10560 -3811
<< viali >>
rect -2579 4403 -2545 4437
rect -2507 4403 -2477 4437
rect -2477 4403 -2473 4437
rect -2435 4403 -2409 4437
rect -2409 4403 -2401 4437
rect -2363 4403 -2341 4437
rect -2341 4403 -2329 4437
rect -2291 4403 -2273 4437
rect -2273 4403 -2257 4437
rect -2219 4403 -2205 4437
rect -2205 4403 -2185 4437
rect -2147 4403 -2137 4437
rect -2137 4403 -2113 4437
rect -2075 4403 -2069 4437
rect -2069 4403 -2041 4437
rect -2003 4403 -2001 4437
rect -2001 4403 -1969 4437
rect -1931 4403 -1899 4437
rect -1899 4403 -1897 4437
rect -1859 4403 -1831 4437
rect -1831 4403 -1825 4437
rect -1787 4403 -1763 4437
rect -1763 4403 -1753 4437
rect -1715 4403 -1695 4437
rect -1695 4403 -1681 4437
rect -1643 4403 -1627 4437
rect -1627 4403 -1609 4437
rect -1571 4403 -1559 4437
rect -1559 4403 -1537 4437
rect -1499 4403 -1491 4437
rect -1491 4403 -1465 4437
rect -1427 4403 -1423 4437
rect -1423 4403 -1393 4437
rect -1355 4403 -1321 4437
rect -1283 4403 -1253 4437
rect -1253 4403 -1249 4437
rect -1211 4403 -1185 4437
rect -1185 4403 -1177 4437
rect -1139 4403 -1117 4437
rect -1117 4403 -1105 4437
rect -1067 4403 -1049 4437
rect -1049 4403 -1033 4437
rect -995 4403 -981 4437
rect -981 4403 -961 4437
rect -923 4403 -913 4437
rect -913 4403 -889 4437
rect -851 4403 -845 4437
rect -845 4403 -817 4437
rect -779 4403 -777 4437
rect -777 4403 -745 4437
rect -707 4403 -675 4437
rect -675 4403 -673 4437
rect -635 4403 -607 4437
rect -607 4403 -601 4437
rect -563 4403 -539 4437
rect -539 4403 -529 4437
rect -491 4403 -471 4437
rect -471 4403 -457 4437
rect -419 4403 -403 4437
rect -403 4403 -385 4437
rect -347 4403 -335 4437
rect -335 4403 -313 4437
rect -275 4403 -267 4437
rect -267 4403 -241 4437
rect -203 4403 -199 4437
rect -199 4403 -169 4437
rect -131 4403 -97 4437
rect -59 4403 -29 4437
rect -29 4403 -25 4437
rect 13 4403 39 4437
rect 39 4403 47 4437
rect 85 4403 107 4437
rect 107 4403 119 4437
rect 157 4403 175 4437
rect 175 4403 191 4437
rect 229 4403 243 4437
rect 243 4403 263 4437
rect 301 4403 311 4437
rect 311 4403 335 4437
rect 373 4403 379 4437
rect 379 4403 407 4437
rect 445 4403 447 4437
rect 447 4403 479 4437
rect 517 4403 549 4437
rect 549 4403 551 4437
rect 589 4403 617 4437
rect 617 4403 623 4437
rect 661 4403 685 4437
rect 685 4403 695 4437
rect 733 4403 753 4437
rect 753 4403 767 4437
rect 805 4403 821 4437
rect 821 4403 839 4437
rect 877 4403 889 4437
rect 889 4403 911 4437
rect 949 4403 957 4437
rect 957 4403 983 4437
rect 1021 4403 1025 4437
rect 1025 4403 1055 4437
rect 1093 4403 1127 4437
rect 1165 4403 1195 4437
rect 1195 4403 1199 4437
rect 1237 4403 1263 4437
rect 1263 4403 1271 4437
rect 1309 4403 1331 4437
rect 1331 4403 1343 4437
rect 1381 4403 1399 4437
rect 1399 4403 1415 4437
rect 1453 4403 1467 4437
rect 1467 4403 1487 4437
rect 1525 4403 1535 4437
rect 1535 4403 1559 4437
rect 1597 4403 1603 4437
rect 1603 4403 1631 4437
rect 1669 4403 1671 4437
rect 1671 4403 1703 4437
rect 1741 4403 1773 4437
rect 1773 4403 1775 4437
rect 1813 4403 1841 4437
rect 1841 4403 1847 4437
rect 1885 4403 1909 4437
rect 1909 4403 1919 4437
rect 1957 4403 1977 4437
rect 1977 4403 1991 4437
rect 2029 4403 2045 4437
rect 2045 4403 2063 4437
rect 2101 4403 2113 4437
rect 2113 4403 2135 4437
rect 2173 4403 2181 4437
rect 2181 4403 2207 4437
rect 2245 4403 2249 4437
rect 2249 4403 2279 4437
rect 2317 4403 2351 4437
rect 2389 4403 2419 4437
rect 2419 4403 2423 4437
rect 2461 4403 2487 4437
rect 2487 4403 2495 4437
rect 2533 4403 2555 4437
rect 2555 4403 2567 4437
rect 2605 4403 2623 4437
rect 2623 4403 2639 4437
rect 2677 4403 2691 4437
rect 2691 4403 2711 4437
rect 2749 4403 2759 4437
rect 2759 4403 2783 4437
rect 2821 4403 2827 4437
rect 2827 4403 2855 4437
rect 2893 4403 2895 4437
rect 2895 4403 2927 4437
rect 2965 4403 2997 4437
rect 2997 4403 2999 4437
rect 3037 4403 3065 4437
rect 3065 4403 3071 4437
rect 3109 4403 3133 4437
rect 3133 4403 3143 4437
rect 3181 4403 3201 4437
rect 3201 4403 3215 4437
rect 3253 4403 3269 4437
rect 3269 4403 3287 4437
rect 3325 4403 3337 4437
rect 3337 4403 3359 4437
rect 3397 4403 3405 4437
rect 3405 4403 3431 4437
rect 3469 4403 3473 4437
rect 3473 4403 3503 4437
rect 3541 4403 3575 4437
rect 3613 4403 3643 4437
rect 3643 4403 3647 4437
rect 3685 4403 3711 4437
rect 3711 4403 3719 4437
rect 3757 4403 3779 4437
rect 3779 4403 3791 4437
rect 3829 4403 3847 4437
rect 3847 4403 3863 4437
rect 3901 4403 3915 4437
rect 3915 4403 3935 4437
rect 3973 4403 3983 4437
rect 3983 4403 4007 4437
rect 4045 4403 4051 4437
rect 4051 4403 4079 4437
rect 4117 4403 4119 4437
rect 4119 4403 4151 4437
rect 4189 4403 4221 4437
rect 4221 4403 4223 4437
rect 4261 4403 4289 4437
rect 4289 4403 4295 4437
rect 4333 4403 4357 4437
rect 4357 4403 4367 4437
rect 4405 4403 4425 4437
rect 4425 4403 4439 4437
rect 4477 4403 4493 4437
rect 4493 4403 4511 4437
rect 4549 4403 4561 4437
rect 4561 4403 4583 4437
rect 4621 4403 4629 4437
rect 4629 4403 4655 4437
rect 4693 4403 4697 4437
rect 4697 4403 4727 4437
rect 4765 4403 4799 4437
rect 4837 4403 4867 4437
rect 4867 4403 4871 4437
rect 4909 4403 4935 4437
rect 4935 4403 4943 4437
rect 4981 4403 5003 4437
rect 5003 4403 5015 4437
rect 5053 4403 5071 4437
rect 5071 4403 5087 4437
rect 5125 4403 5139 4437
rect 5139 4403 5159 4437
rect 5197 4403 5207 4437
rect 5207 4403 5231 4437
rect 5269 4403 5275 4437
rect 5275 4403 5303 4437
rect 5341 4403 5343 4437
rect 5343 4403 5375 4437
rect 5413 4403 5445 4437
rect 5445 4403 5447 4437
rect 5485 4403 5513 4437
rect 5513 4403 5519 4437
rect 5557 4403 5581 4437
rect 5581 4403 5591 4437
rect 5629 4403 5649 4437
rect 5649 4403 5663 4437
rect 5701 4403 5717 4437
rect 5717 4403 5735 4437
rect 5773 4403 5785 4437
rect 5785 4403 5807 4437
rect 5845 4403 5853 4437
rect 5853 4403 5879 4437
rect 5917 4403 5921 4437
rect 5921 4403 5951 4437
rect 5989 4403 6023 4437
rect 6061 4403 6091 4437
rect 6091 4403 6095 4437
rect 6133 4403 6159 4437
rect 6159 4403 6167 4437
rect 6205 4403 6227 4437
rect 6227 4403 6239 4437
rect 6277 4403 6295 4437
rect 6295 4403 6311 4437
rect 6349 4403 6363 4437
rect 6363 4403 6383 4437
rect 6421 4403 6431 4437
rect 6431 4403 6455 4437
rect 6493 4403 6499 4437
rect 6499 4403 6527 4437
rect 6565 4403 6567 4437
rect 6567 4403 6599 4437
rect 6637 4403 6669 4437
rect 6669 4403 6671 4437
rect 6709 4403 6737 4437
rect 6737 4403 6743 4437
rect 6781 4403 6805 4437
rect 6805 4403 6815 4437
rect 6853 4403 6873 4437
rect 6873 4403 6887 4437
rect 6925 4403 6941 4437
rect 6941 4403 6959 4437
rect 6997 4403 7009 4437
rect 7009 4403 7031 4437
rect 7069 4403 7077 4437
rect 7077 4403 7103 4437
rect 7141 4403 7145 4437
rect 7145 4403 7175 4437
rect 7213 4403 7247 4437
rect 7285 4403 7315 4437
rect 7315 4403 7319 4437
rect 7357 4403 7383 4437
rect 7383 4403 7391 4437
rect 7429 4403 7451 4437
rect 7451 4403 7463 4437
rect 7501 4403 7519 4437
rect 7519 4403 7535 4437
rect 7573 4403 7587 4437
rect 7587 4403 7607 4437
rect 7645 4403 7655 4437
rect 7655 4403 7679 4437
rect 7717 4403 7723 4437
rect 7723 4403 7751 4437
rect 7789 4403 7791 4437
rect 7791 4403 7823 4437
rect 7861 4403 7893 4437
rect 7893 4403 7895 4437
rect 7933 4403 7961 4437
rect 7961 4403 7967 4437
rect 8005 4403 8029 4437
rect 8029 4403 8039 4437
rect 8077 4403 8097 4437
rect 8097 4403 8111 4437
rect 8149 4403 8165 4437
rect 8165 4403 8183 4437
rect 8221 4403 8233 4437
rect 8233 4403 8255 4437
rect 8293 4403 8301 4437
rect 8301 4403 8327 4437
rect 8365 4403 8369 4437
rect 8369 4403 8399 4437
rect 8437 4403 8471 4437
rect 8509 4403 8539 4437
rect 8539 4403 8543 4437
rect 8581 4403 8607 4437
rect 8607 4403 8615 4437
rect 8653 4403 8675 4437
rect 8675 4403 8687 4437
rect 8725 4403 8743 4437
rect 8743 4403 8759 4437
rect 8797 4403 8811 4437
rect 8811 4403 8831 4437
rect 8869 4403 8879 4437
rect 8879 4403 8903 4437
rect 8941 4403 8947 4437
rect 8947 4403 8975 4437
rect 9013 4403 9015 4437
rect 9015 4403 9047 4437
rect 9085 4403 9117 4437
rect 9117 4403 9119 4437
rect 9157 4403 9185 4437
rect 9185 4403 9191 4437
rect 9229 4403 9253 4437
rect 9253 4403 9263 4437
rect 9301 4403 9321 4437
rect 9321 4403 9335 4437
rect 9373 4403 9389 4437
rect 9389 4403 9407 4437
rect 9445 4403 9457 4437
rect 9457 4403 9479 4437
rect 9517 4403 9525 4437
rect 9525 4403 9551 4437
rect 9589 4403 9593 4437
rect 9593 4403 9623 4437
rect 9661 4403 9695 4437
rect 9733 4403 9763 4437
rect 9763 4403 9767 4437
rect 9805 4403 9831 4437
rect 9831 4403 9839 4437
rect 9877 4403 9899 4437
rect 9899 4403 9911 4437
rect 9949 4403 9967 4437
rect 9967 4403 9983 4437
rect 10021 4403 10035 4437
rect 10035 4403 10055 4437
rect 10093 4403 10103 4437
rect 10103 4403 10127 4437
rect 10165 4403 10171 4437
rect 10171 4403 10199 4437
rect 10237 4403 10239 4437
rect 10239 4403 10271 4437
rect 10309 4403 10341 4437
rect 10341 4403 10343 4437
rect 10381 4403 10409 4437
rect 10409 4403 10415 4437
rect 10453 4403 10477 4437
rect 10477 4403 10487 4437
rect 10525 4403 10545 4437
rect 10545 4403 10559 4437
rect 10597 4403 10613 4437
rect 10613 4403 10631 4437
rect 10669 4403 10681 4437
rect 10681 4403 10703 4437
rect 10741 4403 10749 4437
rect 10749 4403 10775 4437
rect 10813 4403 10817 4437
rect 10817 4403 10847 4437
rect 10885 4403 10919 4437
rect -2347 4103 -2313 4137
rect -1867 4103 -1833 4137
rect -1427 4103 -1393 4137
rect -967 4103 -933 4137
rect -507 4103 -473 4137
rect -47 4103 -13 4137
rect 413 4103 447 4137
rect 2933 4103 2967 4137
rect 3393 4103 3427 4137
rect 3853 4103 3887 4137
rect 4313 4103 4347 4137
rect 4753 4103 4787 4137
rect 5233 4103 5267 4137
rect 5713 4103 5747 4137
rect 7953 4103 7987 4137
rect 8393 4103 8427 4137
rect 8853 4103 8887 4137
rect 9313 4103 9347 4137
rect 9773 4103 9807 4137
rect 10233 4103 10267 4137
rect 10693 4103 10727 4137
rect -2577 3719 -2543 3753
rect -2577 3647 -2543 3681
rect -1657 3719 -1623 3753
rect -1657 3647 -1623 3681
rect -737 3699 -703 3733
rect -737 3627 -703 3661
rect 163 3719 197 3753
rect 163 3647 197 3681
rect 743 3709 777 3743
rect 743 3637 777 3671
rect 2703 3699 2737 3733
rect 2703 3627 2737 3661
rect 3623 3725 3657 3759
rect 3623 3653 3657 3687
rect 3623 3581 3657 3615
rect 4543 3725 4577 3759
rect 4543 3653 4577 3687
rect 4543 3581 4577 3615
rect 5463 3725 5497 3759
rect 5463 3653 5497 3687
rect 6023 3709 6057 3743
rect 6023 3637 6057 3671
rect 7603 3689 7637 3723
rect 5463 3581 5497 3615
rect 7603 3617 7637 3651
rect 7723 3679 7757 3713
rect 7723 3607 7757 3641
rect 8643 3679 8677 3713
rect 8643 3607 8677 3641
rect 9563 3679 9597 3713
rect 9563 3607 9597 3641
rect 10483 3679 10517 3713
rect 10483 3607 10517 3641
rect -2097 2993 -2063 3027
rect -1197 2993 -1163 3027
rect -277 2993 -243 3027
rect 643 2993 677 3027
rect 3163 2979 3197 3013
rect 3163 2907 3197 2941
rect 4083 2979 4117 3013
rect 4083 2907 4117 2941
rect 5003 2979 5037 3013
rect 5003 2907 5037 2941
rect 5903 2979 5937 3013
rect 5903 2907 5937 2941
rect 8163 2833 8197 2867
rect 9083 2833 9117 2867
rect 10003 2833 10037 2867
rect 10903 2833 10937 2867
rect -511 2573 -477 2607
rect -439 2573 -405 2607
rect -1277 2303 -1243 2337
rect 4027 2303 4061 2337
rect 4099 2303 4133 2337
rect 6913 2263 6947 2297
rect 1294 2101 1328 2135
rect 1366 2101 1400 2135
rect 4047 2103 4081 2137
rect 4119 2103 4153 2137
rect 6887 2103 6921 2137
rect 6959 2103 6993 2137
rect 1294 1980 1328 2014
rect 1366 1980 1400 2014
rect 4073 2003 4107 2037
rect 6897 2003 6931 2037
rect 6969 2003 7003 2037
rect 2306 1852 2340 1886
rect 3363 1853 3397 1887
rect 4686 1878 4720 1912
rect 4686 1806 4720 1840
rect 6163 1853 6197 1887
rect 2053 1714 2087 1748
rect 2125 1714 2159 1748
rect 3567 1723 3601 1757
rect 3639 1723 3673 1757
rect 6897 1723 6931 1757
rect 6969 1723 7003 1757
rect 2083 1131 2117 1165
rect 6897 1163 6931 1197
rect 6969 1163 7003 1197
rect 2083 1059 2117 1093
rect 2083 987 2117 1021
rect 6143 1023 6177 1057
rect 2083 915 2117 949
rect 6607 903 6641 937
rect 6679 903 6713 937
rect 7527 903 7561 937
rect 7599 903 7633 937
rect 1063 799 1097 833
rect 4967 823 5001 857
rect 5039 823 5073 857
rect 6643 783 6677 817
rect 1063 727 1097 761
rect 2875 686 2909 720
rect 5383 683 5417 717
rect 3703 543 3737 577
rect 2083 437 2117 471
rect 3693 443 3727 477
rect -1897 349 -1863 383
rect -1897 277 -1863 311
rect -1797 349 -1763 383
rect -1797 277 -1763 311
rect -1337 352 -1303 386
rect -1337 280 -1303 314
rect -17 329 17 363
rect -17 257 17 291
rect 83 339 117 373
rect 83 267 117 301
rect 547 338 581 372
rect 547 266 581 300
rect 2083 365 2117 399
rect 2083 293 2117 327
rect 2083 221 2117 255
rect 311 131 345 165
rect 2083 149 2117 183
rect 5763 183 5797 217
rect -1593 53 -1559 87
rect -1521 53 -1487 87
rect 2783 -631 2817 -597
rect 2783 -703 2817 -669
rect 3703 -631 3737 -597
rect 3703 -703 3737 -669
rect 4623 -611 4657 -577
rect 4623 -683 4657 -649
rect 5543 -611 5577 -577
rect 5543 -683 5577 -649
rect 6643 -621 6677 -587
rect 6643 -693 6677 -659
rect 7563 -621 7597 -587
rect 7563 -693 7597 -659
rect 8483 -601 8517 -567
rect 8483 -673 8517 -639
rect 9403 -601 9437 -567
rect 9403 -673 9437 -639
rect 3243 -1127 3277 -1093
rect 4163 -1127 4197 -1093
rect 5083 -1127 5117 -1093
rect 6003 -1127 6037 -1093
rect 6103 -1137 6137 -1103
rect 7103 -1127 7137 -1093
rect 8023 -1127 8057 -1093
rect 8943 -1127 8977 -1093
rect 9863 -1127 9897 -1093
rect 9963 -1117 9997 -1083
rect 2987 -1337 3021 -1303
rect 3059 -1337 3093 -1303
rect 3467 -1337 3501 -1303
rect 3539 -1337 3573 -1303
rect 3907 -1337 3941 -1303
rect 3979 -1337 4013 -1303
rect 4367 -1337 4401 -1303
rect 4439 -1337 4473 -1303
rect 4847 -1337 4881 -1303
rect 4919 -1337 4953 -1303
rect 5287 -1337 5321 -1303
rect 5359 -1337 5393 -1303
rect 5747 -1337 5781 -1303
rect 5819 -1337 5853 -1303
rect 6847 -1337 6881 -1303
rect 6919 -1337 6953 -1303
rect 7327 -1337 7361 -1303
rect 7399 -1337 7433 -1303
rect 7767 -1337 7801 -1303
rect 7839 -1337 7873 -1303
rect 8227 -1337 8261 -1303
rect 8299 -1337 8333 -1303
rect 8687 -1337 8721 -1303
rect 8759 -1337 8793 -1303
rect 9167 -1337 9201 -1303
rect 9239 -1337 9273 -1303
rect 9627 -1337 9661 -1303
rect 9699 -1337 9733 -1303
rect -1777 -2297 -1743 -2263
rect -857 -2297 -823 -2263
rect 63 -2297 97 -2263
rect 983 -2297 1017 -2263
rect 1903 -2297 1937 -2263
rect 2803 -2297 2837 -2263
rect 4963 -2327 4997 -2293
rect 5883 -2327 5917 -2293
rect 6803 -2327 6837 -2293
rect 7723 -2327 7757 -2293
rect 8643 -2327 8677 -2293
rect 9543 -2347 9577 -2313
rect 10463 -2347 10497 -2313
rect -2177 -3177 -2143 -3143
rect -2057 -3141 -2023 -3107
rect -2057 -3213 -2023 -3179
rect -1877 -3187 -1843 -3153
rect -1317 -3177 -1283 -3143
rect -397 -3177 -363 -3143
rect 523 -3177 557 -3143
rect 1443 -3177 1477 -3143
rect 2343 -3177 2377 -3143
rect 3893 -3177 3927 -3143
rect 4863 -3177 4897 -3143
rect 5423 -3177 5457 -3143
rect 6343 -3177 6377 -3143
rect 7263 -3177 7297 -3143
rect 8163 -3177 8197 -3143
rect 9083 -3177 9117 -3143
rect 10003 -3177 10037 -3143
rect -2637 -3367 -2603 -3333
rect -2463 -3477 -2429 -3443
rect -2391 -3477 -2357 -3443
rect -1583 -3477 -1549 -3443
rect -1511 -3477 -1477 -3443
rect -1123 -3477 -1089 -3443
rect -1051 -3477 -1017 -3443
rect -663 -3477 -629 -3443
rect -591 -3477 -557 -3443
rect -243 -3477 -209 -3443
rect -171 -3477 -137 -3443
rect 237 -3477 271 -3443
rect 309 -3477 343 -3443
rect 697 -3477 731 -3443
rect 769 -3477 803 -3443
rect 1157 -3477 1191 -3443
rect 1229 -3477 1263 -3443
rect 1617 -3477 1651 -3443
rect 1689 -3477 1723 -3443
rect 2077 -3477 2111 -3443
rect 2149 -3477 2183 -3443
rect 2557 -3477 2591 -3443
rect 2629 -3477 2663 -3443
rect 5167 -3477 5201 -3443
rect 5239 -3477 5273 -3443
rect 5627 -3477 5661 -3443
rect 5699 -3477 5733 -3443
rect 6087 -3477 6121 -3443
rect 6159 -3477 6193 -3443
rect 6547 -3477 6581 -3443
rect 6619 -3477 6653 -3443
rect 7007 -3477 7041 -3443
rect 7079 -3477 7113 -3443
rect 7447 -3477 7481 -3443
rect 7519 -3477 7553 -3443
rect 7907 -3477 7941 -3443
rect 7979 -3477 8013 -3443
rect 8367 -3477 8401 -3443
rect 8439 -3477 8473 -3443
rect 8847 -3477 8881 -3443
rect 8919 -3477 8953 -3443
rect 9287 -3477 9321 -3443
rect 9359 -3477 9393 -3443
rect 9747 -3477 9781 -3443
rect 9819 -3477 9853 -3443
rect 10207 -3477 10241 -3443
rect 10279 -3477 10313 -3443
rect -2639 -3777 -2616 -3743
rect -2616 -3777 -2605 -3743
rect -2567 -3777 -2548 -3743
rect -2548 -3777 -2533 -3743
rect -2495 -3777 -2480 -3743
rect -2480 -3777 -2461 -3743
rect -2423 -3777 -2412 -3743
rect -2412 -3777 -2389 -3743
rect -2351 -3777 -2344 -3743
rect -2344 -3777 -2317 -3743
rect -2279 -3777 -2276 -3743
rect -2276 -3777 -2245 -3743
rect -2207 -3777 -2174 -3743
rect -2174 -3777 -2173 -3743
rect -2135 -3777 -2106 -3743
rect -2106 -3777 -2101 -3743
rect -2063 -3777 -2038 -3743
rect -2038 -3777 -2029 -3743
rect -1991 -3777 -1970 -3743
rect -1970 -3777 -1957 -3743
rect -1919 -3777 -1902 -3743
rect -1902 -3777 -1885 -3743
rect -1847 -3777 -1834 -3743
rect -1834 -3777 -1813 -3743
rect -1775 -3777 -1766 -3743
rect -1766 -3777 -1741 -3743
rect -1703 -3777 -1698 -3743
rect -1698 -3777 -1669 -3743
rect -1631 -3777 -1603 -3743
rect -1603 -3777 -1597 -3743
rect -1559 -3777 -1525 -3743
rect -1487 -3777 -1453 -3743
rect -1415 -3777 -1381 -3743
rect -1343 -3777 -1309 -3743
rect -1271 -3777 -1237 -3743
rect -1199 -3777 -1165 -3743
rect -1127 -3777 -1093 -3743
rect -1055 -3777 -1021 -3743
rect -983 -3777 -949 -3743
rect -911 -3777 -877 -3743
rect -839 -3777 -805 -3743
rect -767 -3777 -733 -3743
rect -695 -3777 -661 -3743
rect -623 -3777 -589 -3743
rect -551 -3777 -517 -3743
rect -479 -3777 -445 -3743
rect -407 -3777 -373 -3743
rect -335 -3777 -301 -3743
rect -263 -3777 -229 -3743
rect -191 -3777 -157 -3743
rect -119 -3777 -85 -3743
rect -47 -3777 -13 -3743
rect 25 -3777 59 -3743
rect 97 -3777 131 -3743
rect 169 -3777 203 -3743
rect 241 -3777 275 -3743
rect 313 -3777 347 -3743
rect 385 -3777 419 -3743
rect 457 -3777 491 -3743
rect 529 -3777 563 -3743
rect 601 -3777 635 -3743
rect 673 -3777 707 -3743
rect 745 -3777 779 -3743
rect 817 -3777 851 -3743
rect 889 -3777 923 -3743
rect 961 -3777 995 -3743
rect 1033 -3777 1067 -3743
rect 1105 -3777 1139 -3743
rect 1177 -3777 1211 -3743
rect 1249 -3777 1283 -3743
rect 1321 -3777 1355 -3743
rect 1393 -3777 1427 -3743
rect 1465 -3777 1499 -3743
rect 1537 -3777 1571 -3743
rect 1609 -3777 1643 -3743
rect 1681 -3777 1715 -3743
rect 1753 -3777 1787 -3743
rect 1825 -3777 1859 -3743
rect 1897 -3777 1931 -3743
rect 1969 -3777 2003 -3743
rect 2041 -3777 2075 -3743
rect 2113 -3777 2147 -3743
rect 2185 -3777 2219 -3743
rect 2257 -3777 2291 -3743
rect 2329 -3777 2363 -3743
rect 2401 -3777 2435 -3743
rect 2473 -3777 2507 -3743
rect 2545 -3777 2579 -3743
rect 2617 -3777 2651 -3743
rect 2689 -3777 2723 -3743
rect 2761 -3777 2783 -3743
rect 2783 -3777 2795 -3743
rect 2833 -3777 2852 -3743
rect 2852 -3777 2867 -3743
rect 2905 -3777 2920 -3743
rect 2920 -3777 2939 -3743
rect 2977 -3777 2988 -3743
rect 2988 -3777 3011 -3743
rect 3049 -3777 3056 -3743
rect 3056 -3777 3083 -3743
rect 3121 -3777 3124 -3743
rect 3124 -3777 3155 -3743
rect 3193 -3777 3226 -3743
rect 3226 -3777 3227 -3743
rect 3265 -3777 3294 -3743
rect 3294 -3777 3299 -3743
rect 3337 -3777 3362 -3743
rect 3362 -3777 3371 -3743
rect 3409 -3777 3430 -3743
rect 3430 -3777 3443 -3743
rect 3481 -3777 3498 -3743
rect 3498 -3777 3515 -3743
rect 3553 -3777 3566 -3743
rect 3566 -3777 3587 -3743
rect 3625 -3777 3634 -3743
rect 3634 -3777 3659 -3743
rect 3697 -3777 3702 -3743
rect 3702 -3777 3731 -3743
rect 3769 -3777 3770 -3743
rect 3770 -3777 3803 -3743
rect 3841 -3777 3872 -3743
rect 3872 -3777 3875 -3743
rect 3913 -3777 3940 -3743
rect 3940 -3777 3947 -3743
rect 3985 -3777 4008 -3743
rect 4008 -3777 4019 -3743
rect 4057 -3777 4076 -3743
rect 4076 -3777 4091 -3743
rect 4129 -3777 4144 -3743
rect 4144 -3777 4163 -3743
rect 4201 -3777 4212 -3743
rect 4212 -3777 4235 -3743
rect 4273 -3777 4280 -3743
rect 4280 -3777 4307 -3743
rect 4345 -3777 4348 -3743
rect 4348 -3777 4379 -3743
rect 4417 -3777 4450 -3743
rect 4450 -3777 4451 -3743
rect 4489 -3777 4518 -3743
rect 4518 -3777 4523 -3743
rect 4561 -3777 4586 -3743
rect 4586 -3777 4595 -3743
rect 4633 -3777 4654 -3743
rect 4654 -3777 4667 -3743
rect 4705 -3777 4722 -3743
rect 4722 -3777 4739 -3743
rect 4777 -3777 4790 -3743
rect 4790 -3777 4811 -3743
rect 4849 -3777 4858 -3743
rect 4858 -3777 4883 -3743
rect 4921 -3777 4926 -3743
rect 4926 -3777 4955 -3743
rect 4993 -3777 4994 -3743
rect 4994 -3777 5027 -3743
rect 5065 -3777 5096 -3743
rect 5096 -3777 5099 -3743
rect 5137 -3777 5164 -3743
rect 5164 -3777 5171 -3743
rect 5209 -3777 5232 -3743
rect 5232 -3777 5243 -3743
rect 5281 -3777 5300 -3743
rect 5300 -3777 5315 -3743
rect 5353 -3777 5368 -3743
rect 5368 -3777 5387 -3743
rect 5425 -3777 5436 -3743
rect 5436 -3777 5459 -3743
rect 5497 -3777 5504 -3743
rect 5504 -3777 5531 -3743
rect 5569 -3777 5572 -3743
rect 5572 -3777 5603 -3743
rect 5641 -3777 5674 -3743
rect 5674 -3777 5675 -3743
rect 5713 -3777 5742 -3743
rect 5742 -3777 5747 -3743
rect 5785 -3777 5810 -3743
rect 5810 -3777 5819 -3743
rect 5857 -3777 5878 -3743
rect 5878 -3777 5891 -3743
rect 5929 -3777 5946 -3743
rect 5946 -3777 5963 -3743
rect 6001 -3777 6014 -3743
rect 6014 -3777 6035 -3743
rect 6073 -3777 6082 -3743
rect 6082 -3777 6107 -3743
rect 6145 -3777 6150 -3743
rect 6150 -3777 6179 -3743
rect 6217 -3777 6218 -3743
rect 6218 -3777 6251 -3743
rect 6289 -3777 6320 -3743
rect 6320 -3777 6323 -3743
rect 6361 -3777 6388 -3743
rect 6388 -3777 6395 -3743
rect 6433 -3777 6456 -3743
rect 6456 -3777 6467 -3743
rect 6505 -3777 6524 -3743
rect 6524 -3777 6539 -3743
rect 6577 -3777 6592 -3743
rect 6592 -3777 6611 -3743
rect 6649 -3777 6660 -3743
rect 6660 -3777 6683 -3743
rect 6721 -3777 6728 -3743
rect 6728 -3777 6755 -3743
rect 6793 -3777 6796 -3743
rect 6796 -3777 6827 -3743
rect 6865 -3777 6898 -3743
rect 6898 -3777 6899 -3743
rect 6937 -3777 6966 -3743
rect 6966 -3777 6971 -3743
rect 7009 -3777 7034 -3743
rect 7034 -3777 7043 -3743
rect 7081 -3777 7102 -3743
rect 7102 -3777 7115 -3743
rect 7153 -3777 7170 -3743
rect 7170 -3777 7187 -3743
rect 7225 -3777 7238 -3743
rect 7238 -3777 7259 -3743
rect 7297 -3777 7306 -3743
rect 7306 -3777 7331 -3743
rect 7369 -3777 7374 -3743
rect 7374 -3777 7403 -3743
rect 7441 -3777 7442 -3743
rect 7442 -3777 7475 -3743
rect 7513 -3777 7544 -3743
rect 7544 -3777 7547 -3743
rect 7585 -3777 7612 -3743
rect 7612 -3777 7619 -3743
rect 7657 -3777 7680 -3743
rect 7680 -3777 7691 -3743
rect 7729 -3777 7748 -3743
rect 7748 -3777 7763 -3743
rect 7801 -3777 7816 -3743
rect 7816 -3777 7835 -3743
rect 7873 -3777 7884 -3743
rect 7884 -3777 7907 -3743
rect 7945 -3777 7952 -3743
rect 7952 -3777 7979 -3743
rect 8017 -3777 8020 -3743
rect 8020 -3777 8051 -3743
rect 8089 -3777 8122 -3743
rect 8122 -3777 8123 -3743
rect 8161 -3777 8190 -3743
rect 8190 -3777 8195 -3743
rect 8233 -3777 8258 -3743
rect 8258 -3777 8267 -3743
rect 8305 -3777 8326 -3743
rect 8326 -3777 8339 -3743
rect 8377 -3777 8394 -3743
rect 8394 -3777 8411 -3743
rect 8449 -3777 8462 -3743
rect 8462 -3777 8483 -3743
rect 8521 -3777 8530 -3743
rect 8530 -3777 8555 -3743
rect 8593 -3777 8598 -3743
rect 8598 -3777 8627 -3743
rect 8665 -3777 8666 -3743
rect 8666 -3777 8699 -3743
rect 8737 -3777 8768 -3743
rect 8768 -3777 8771 -3743
rect 8809 -3777 8836 -3743
rect 8836 -3777 8843 -3743
rect 8881 -3777 8904 -3743
rect 8904 -3777 8915 -3743
rect 8953 -3777 8972 -3743
rect 8972 -3777 8987 -3743
rect 9025 -3777 9040 -3743
rect 9040 -3777 9059 -3743
rect 9097 -3777 9108 -3743
rect 9108 -3777 9131 -3743
rect 9169 -3777 9176 -3743
rect 9176 -3777 9203 -3743
rect 9241 -3777 9244 -3743
rect 9244 -3777 9275 -3743
rect 9313 -3777 9346 -3743
rect 9346 -3777 9347 -3743
rect 9385 -3777 9414 -3743
rect 9414 -3777 9419 -3743
rect 9457 -3777 9482 -3743
rect 9482 -3777 9491 -3743
rect 9529 -3777 9550 -3743
rect 9550 -3777 9563 -3743
rect 9601 -3777 9618 -3743
rect 9618 -3777 9635 -3743
rect 9673 -3777 9686 -3743
rect 9686 -3777 9707 -3743
rect 9745 -3777 9754 -3743
rect 9754 -3777 9779 -3743
rect 9817 -3777 9822 -3743
rect 9822 -3777 9851 -3743
rect 9889 -3777 9890 -3743
rect 9890 -3777 9923 -3743
rect 9961 -3777 9992 -3743
rect 9992 -3777 9995 -3743
rect 10033 -3777 10060 -3743
rect 10060 -3777 10067 -3743
rect 10105 -3777 10128 -3743
rect 10128 -3777 10139 -3743
rect 10177 -3777 10196 -3743
rect 10196 -3777 10211 -3743
rect 10249 -3777 10264 -3743
rect 10264 -3777 10283 -3743
rect 10321 -3777 10332 -3743
rect 10332 -3777 10355 -3743
rect 10393 -3777 10400 -3743
rect 10400 -3777 10427 -3743
rect 10465 -3777 10468 -3743
rect 10468 -3777 10499 -3743
<< metal1 >>
rect -2700 4437 11060 4520
rect -3480 4340 -3040 4420
rect -2700 4403 -2579 4437
rect -2545 4403 -2507 4437
rect -2473 4403 -2435 4437
rect -2401 4403 -2363 4437
rect -2329 4403 -2291 4437
rect -2257 4403 -2219 4437
rect -2185 4403 -2147 4437
rect -2113 4403 -2075 4437
rect -2041 4403 -2003 4437
rect -1969 4403 -1931 4437
rect -1897 4403 -1859 4437
rect -1825 4403 -1787 4437
rect -1753 4403 -1715 4437
rect -1681 4403 -1643 4437
rect -1609 4403 -1571 4437
rect -1537 4403 -1499 4437
rect -1465 4403 -1427 4437
rect -1393 4403 -1355 4437
rect -1321 4403 -1283 4437
rect -1249 4403 -1211 4437
rect -1177 4403 -1139 4437
rect -1105 4403 -1067 4437
rect -1033 4403 -995 4437
rect -961 4403 -923 4437
rect -889 4403 -851 4437
rect -817 4403 -779 4437
rect -745 4403 -707 4437
rect -673 4403 -635 4437
rect -601 4403 -563 4437
rect -529 4403 -491 4437
rect -457 4403 -419 4437
rect -385 4403 -347 4437
rect -313 4403 -275 4437
rect -241 4403 -203 4437
rect -169 4403 -131 4437
rect -97 4403 -59 4437
rect -25 4403 13 4437
rect 47 4403 85 4437
rect 119 4403 157 4437
rect 191 4403 229 4437
rect 263 4403 301 4437
rect 335 4403 373 4437
rect 407 4403 445 4437
rect 479 4403 517 4437
rect 551 4403 589 4437
rect 623 4403 661 4437
rect 695 4403 733 4437
rect 767 4403 805 4437
rect 839 4403 877 4437
rect 911 4403 949 4437
rect 983 4403 1021 4437
rect 1055 4403 1093 4437
rect 1127 4403 1165 4437
rect 1199 4403 1237 4437
rect 1271 4403 1309 4437
rect 1343 4403 1381 4437
rect 1415 4403 1453 4437
rect 1487 4403 1525 4437
rect 1559 4403 1597 4437
rect 1631 4403 1669 4437
rect 1703 4403 1741 4437
rect 1775 4403 1813 4437
rect 1847 4403 1885 4437
rect 1919 4403 1957 4437
rect 1991 4403 2029 4437
rect 2063 4403 2101 4437
rect 2135 4403 2173 4437
rect 2207 4403 2245 4437
rect 2279 4403 2317 4437
rect 2351 4403 2389 4437
rect 2423 4403 2461 4437
rect 2495 4403 2533 4437
rect 2567 4403 2605 4437
rect 2639 4403 2677 4437
rect 2711 4403 2749 4437
rect 2783 4403 2821 4437
rect 2855 4403 2893 4437
rect 2927 4403 2965 4437
rect 2999 4403 3037 4437
rect 3071 4403 3109 4437
rect 3143 4403 3181 4437
rect 3215 4403 3253 4437
rect 3287 4403 3325 4437
rect 3359 4403 3397 4437
rect 3431 4403 3469 4437
rect 3503 4403 3541 4437
rect 3575 4403 3613 4437
rect 3647 4403 3685 4437
rect 3719 4403 3757 4437
rect 3791 4403 3829 4437
rect 3863 4403 3901 4437
rect 3935 4403 3973 4437
rect 4007 4403 4045 4437
rect 4079 4403 4117 4437
rect 4151 4403 4189 4437
rect 4223 4403 4261 4437
rect 4295 4403 4333 4437
rect 4367 4403 4405 4437
rect 4439 4403 4477 4437
rect 4511 4403 4549 4437
rect 4583 4403 4621 4437
rect 4655 4403 4693 4437
rect 4727 4403 4765 4437
rect 4799 4403 4837 4437
rect 4871 4403 4909 4437
rect 4943 4403 4981 4437
rect 5015 4403 5053 4437
rect 5087 4403 5125 4437
rect 5159 4403 5197 4437
rect 5231 4403 5269 4437
rect 5303 4403 5341 4437
rect 5375 4403 5413 4437
rect 5447 4403 5485 4437
rect 5519 4403 5557 4437
rect 5591 4403 5629 4437
rect 5663 4403 5701 4437
rect 5735 4403 5773 4437
rect 5807 4403 5845 4437
rect 5879 4403 5917 4437
rect 5951 4403 5989 4437
rect 6023 4403 6061 4437
rect 6095 4403 6133 4437
rect 6167 4403 6205 4437
rect 6239 4403 6277 4437
rect 6311 4403 6349 4437
rect 6383 4403 6421 4437
rect 6455 4403 6493 4437
rect 6527 4403 6565 4437
rect 6599 4403 6637 4437
rect 6671 4403 6709 4437
rect 6743 4403 6781 4437
rect 6815 4403 6853 4437
rect 6887 4403 6925 4437
rect 6959 4403 6997 4437
rect 7031 4403 7069 4437
rect 7103 4403 7141 4437
rect 7175 4403 7213 4437
rect 7247 4403 7285 4437
rect 7319 4403 7357 4437
rect 7391 4403 7429 4437
rect 7463 4403 7501 4437
rect 7535 4403 7573 4437
rect 7607 4403 7645 4437
rect 7679 4403 7717 4437
rect 7751 4403 7789 4437
rect 7823 4403 7861 4437
rect 7895 4403 7933 4437
rect 7967 4403 8005 4437
rect 8039 4403 8077 4437
rect 8111 4403 8149 4437
rect 8183 4403 8221 4437
rect 8255 4403 8293 4437
rect 8327 4403 8365 4437
rect 8399 4403 8437 4437
rect 8471 4403 8509 4437
rect 8543 4403 8581 4437
rect 8615 4403 8653 4437
rect 8687 4403 8725 4437
rect 8759 4403 8797 4437
rect 8831 4403 8869 4437
rect 8903 4403 8941 4437
rect 8975 4403 9013 4437
rect 9047 4403 9085 4437
rect 9119 4403 9157 4437
rect 9191 4403 9229 4437
rect 9263 4403 9301 4437
rect 9335 4403 9373 4437
rect 9407 4403 9445 4437
rect 9479 4403 9517 4437
rect 9551 4403 9589 4437
rect 9623 4403 9661 4437
rect 9695 4403 9733 4437
rect 9767 4403 9805 4437
rect 9839 4403 9877 4437
rect 9911 4403 9949 4437
rect 9983 4403 10021 4437
rect 10055 4403 10093 4437
rect 10127 4403 10165 4437
rect 10199 4403 10237 4437
rect 10271 4403 10309 4437
rect 10343 4403 10381 4437
rect 10415 4403 10453 4437
rect 10487 4403 10525 4437
rect 10559 4403 10597 4437
rect 10631 4403 10669 4437
rect 10703 4403 10741 4437
rect 10775 4403 10813 4437
rect 10847 4403 10885 4437
rect 10919 4403 11060 4437
rect -2700 4340 11060 4403
rect -3480 4338 -2520 4340
rect -3480 4222 -3340 4338
rect -3160 4240 -2520 4338
rect -3160 4222 -3040 4240
rect -3480 4120 -3040 4222
rect -2620 3800 -2520 4240
rect -2420 4137 10920 4160
rect -2420 4103 -2347 4137
rect -2313 4103 -1867 4137
rect -1833 4103 -1427 4137
rect -1393 4103 -967 4137
rect -933 4103 -507 4137
rect -473 4103 -47 4137
rect -13 4103 413 4137
rect 447 4103 2933 4137
rect 2967 4103 3393 4137
rect 3427 4103 3853 4137
rect 3887 4103 4313 4137
rect 4347 4103 4753 4137
rect 4787 4103 5233 4137
rect 5267 4103 5713 4137
rect 5747 4103 7953 4137
rect 7987 4103 8393 4137
rect 8427 4103 8853 4137
rect 8887 4103 9313 4137
rect 9347 4103 9773 4137
rect 9807 4103 10233 4137
rect 10267 4103 10693 4137
rect 10727 4103 10920 4137
rect -2420 4080 10920 4103
rect 2680 3800 5960 3820
rect -2620 3759 10560 3800
rect -2620 3753 3623 3759
rect -2620 3719 -2577 3753
rect -2543 3719 -1657 3753
rect -1623 3733 163 3753
rect -1623 3719 -737 3733
rect -2620 3699 -737 3719
rect -703 3719 163 3733
rect 197 3743 3623 3753
rect 197 3719 743 3743
rect -703 3709 743 3719
rect 777 3733 3623 3743
rect 777 3709 2703 3733
rect -703 3699 2703 3709
rect 2737 3725 3623 3733
rect 3657 3725 4543 3759
rect 4577 3725 5463 3759
rect 5497 3743 10560 3759
rect 5497 3725 6023 3743
rect 2737 3709 6023 3725
rect 6057 3723 10560 3743
rect 6057 3709 7603 3723
rect 2737 3699 7603 3709
rect -2620 3689 7603 3699
rect 7637 3713 10560 3723
rect 7637 3689 7723 3713
rect -2620 3687 7723 3689
rect -2620 3681 3623 3687
rect -2620 3647 -2577 3681
rect -2543 3647 -1657 3681
rect -1623 3661 163 3681
rect -1623 3647 -737 3661
rect -2620 3627 -737 3647
rect -703 3647 163 3661
rect 197 3671 3623 3681
rect 197 3647 743 3671
rect -703 3637 743 3647
rect 777 3661 3623 3671
rect 777 3637 2703 3661
rect -703 3627 2703 3637
rect 2737 3653 3623 3661
rect 3657 3653 4543 3687
rect 4577 3653 5463 3687
rect 5497 3679 7723 3687
rect 7757 3679 8643 3713
rect 8677 3679 9563 3713
rect 9597 3679 10483 3713
rect 10517 3679 10560 3713
rect 5497 3671 10560 3679
rect 5497 3653 6023 3671
rect 2737 3637 6023 3653
rect 6057 3651 10560 3671
rect 6057 3637 7603 3651
rect 2737 3627 7603 3637
rect -2620 3617 7603 3627
rect 7637 3641 10560 3651
rect 7637 3617 7723 3641
rect -2620 3615 7723 3617
rect -2620 3581 3623 3615
rect 3657 3581 4543 3615
rect 4577 3581 5463 3615
rect 5497 3607 7723 3615
rect 7757 3607 8643 3641
rect 8677 3607 9563 3641
rect 9597 3607 10483 3641
rect 10517 3607 10560 3641
rect 5497 3581 10560 3607
rect -2620 3540 10560 3581
rect -2120 3120 700 3140
rect -2120 3027 1480 3120
rect -2120 2993 -2097 3027
rect -2063 2993 -1197 3027
rect -1163 2993 -277 3027
rect -243 2993 643 3027
rect 677 2993 1480 3027
rect -2120 2880 1480 2993
rect 1200 2660 1480 2880
rect 3140 3013 5960 3200
rect 3140 2979 3163 3013
rect 3197 2979 4083 3013
rect 4117 2979 5003 3013
rect 5037 2979 5903 3013
rect 5937 2979 5960 3013
rect 3140 2941 5960 2979
rect 3140 2907 3163 2941
rect 3197 2907 4083 2941
rect 4117 2907 5003 2941
rect 5037 2907 5903 2941
rect 5937 2907 5960 2941
rect 3140 2840 5960 2907
rect 6800 2867 10960 3000
rect -561 2607 -371 2627
rect -561 2573 -511 2607
rect -477 2573 -439 2607
rect -405 2573 -371 2607
rect -1340 2346 -1160 2380
rect -1340 2294 -1296 2346
rect -1244 2337 -1160 2346
rect -1243 2303 -1160 2337
rect -1244 2294 -1160 2303
rect -1340 2220 -1160 2294
rect -1340 1038 -1260 2220
rect -561 1750 -371 2573
rect 1200 2135 1487 2660
rect 1200 2101 1294 2135
rect 1328 2101 1366 2135
rect 1400 2101 1487 2135
rect 1200 2014 1487 2101
rect 1200 1980 1294 2014
rect 1328 1980 1366 2014
rect 1400 1980 1487 2014
rect 3980 2337 4200 2840
rect 3980 2336 4027 2337
rect 4061 2336 4099 2337
rect 4133 2336 4200 2337
rect 3980 2284 3990 2336
rect 4042 2284 4054 2303
rect 4106 2284 4118 2303
rect 4170 2284 4200 2336
rect 3980 2137 4200 2284
rect 3980 2103 4047 2137
rect 4081 2103 4119 2137
rect 4153 2103 4200 2137
rect 3980 2037 4200 2103
rect 3980 2003 4073 2037
rect 4107 2003 4200 2037
rect 3980 1980 4200 2003
rect 6800 2833 8163 2867
rect 8197 2833 9083 2867
rect 9117 2833 10003 2867
rect 10037 2833 10903 2867
rect 10937 2833 10960 2867
rect 6800 2720 10960 2833
rect 6800 2338 7100 2720
rect 6800 2222 6840 2338
rect 7020 2222 7100 2338
rect 6800 2137 7100 2222
rect 6800 2103 6887 2137
rect 6921 2103 6959 2137
rect 6993 2103 7100 2137
rect 6800 2037 7100 2103
rect 6800 2003 6897 2037
rect 6931 2003 6969 2037
rect 7003 2003 7100 2037
rect 4665 1980 5040 1983
rect 6800 1980 7100 2003
rect 1200 1968 1487 1980
rect 2780 1979 3420 1980
rect 2301 1974 3420 1979
rect 2275 1887 3420 1974
rect 2275 1886 3363 1887
rect 2275 1852 2306 1886
rect 2340 1853 3363 1886
rect 3397 1853 3420 1887
rect 2340 1852 3420 1853
rect 2275 1780 3420 1852
rect 4665 1912 6220 1980
rect 4665 1878 4686 1912
rect 4720 1887 6220 1912
rect 4720 1878 6163 1887
rect 4665 1853 6163 1878
rect 6197 1853 6220 1887
rect 4665 1840 6220 1853
rect 4665 1806 4686 1840
rect 4720 1806 6220 1840
rect 2275 1767 2878 1780
rect 2014 1750 2184 1760
rect -561 1748 2188 1750
rect -561 1714 2053 1748
rect 2087 1714 2125 1748
rect 2159 1714 2188 1748
rect -561 1676 2188 1714
rect -561 1668 -371 1676
rect 2014 1556 2179 1676
rect 2301 1556 2440 1767
rect 2014 1434 2180 1556
rect -1348 989 -1260 1038
rect 2020 1165 2180 1434
rect 2020 1131 2083 1165
rect 2117 1131 2180 1165
rect 2020 1093 2180 1131
rect 2020 1059 2083 1093
rect 2117 1059 2180 1093
rect 2020 1021 2180 1059
rect -1800 440 -1740 500
rect -1920 383 -1740 440
rect -1920 349 -1897 383
rect -1863 349 -1797 383
rect -1763 349 -1740 383
rect -1920 311 -1740 349
rect -1920 277 -1897 311
rect -1863 277 -1797 311
rect -1763 277 -1740 311
rect -1920 240 -1740 277
rect -1348 386 -1261 989
rect 2020 987 2083 1021
rect 2117 987 2180 1021
rect 2020 949 2180 987
rect 2020 915 2083 949
rect 2117 915 2180 949
rect 526 886 603 888
rect 526 880 947 886
rect 526 838 1180 880
rect 2020 860 2180 915
rect 526 722 990 838
rect 1170 722 1180 838
rect 526 664 1180 722
rect 60 420 120 500
rect -1348 352 -1337 386
rect -1303 352 -1261 386
rect -1348 314 -1261 352
rect -1348 280 -1337 314
rect -1303 280 -1261 314
rect -1348 255 -1261 280
rect -40 373 140 420
rect -40 363 83 373
rect -40 329 -17 363
rect 17 339 83 363
rect 117 339 140 373
rect 17 329 140 339
rect -40 301 140 329
rect -40 291 83 301
rect -40 257 -17 291
rect 17 267 83 291
rect 117 267 140 301
rect 17 257 140 267
rect -1800 -2200 -1740 240
rect -40 220 140 257
rect 526 372 603 664
rect 725 660 1180 664
rect 526 338 547 372
rect 581 338 603 372
rect 526 300 603 338
rect 526 266 547 300
rect 581 266 603 300
rect 526 246 603 266
rect 2020 471 2200 540
rect 2020 437 2083 471
rect 2117 437 2200 471
rect 2020 399 2200 437
rect 2020 365 2083 399
rect 2117 365 2200 399
rect 2020 327 2200 365
rect 2020 293 2083 327
rect 2117 293 2200 327
rect 2020 255 2200 293
rect 2020 221 2083 255
rect 2117 221 2200 255
rect -1640 87 -1440 120
rect -1640 53 -1593 87
rect -1559 53 -1521 87
rect -1487 53 -1440 87
rect -1640 -120 -1440 53
rect -920 -82 -480 0
rect -920 -120 -780 -82
rect -1640 -198 -780 -120
rect -600 -198 -480 -82
rect -1640 -240 -480 -198
rect -1640 -320 -1440 -240
rect -920 -300 -480 -240
rect 60 -2200 120 220
rect 240 165 442 190
rect 240 131 311 165
rect 345 131 442 165
rect 240 96 442 131
rect 2020 183 2200 221
rect 2020 149 2083 183
rect 2117 149 2200 183
rect 2020 120 2200 149
rect 2020 100 2180 120
rect 240 -120 440 96
rect 840 -120 1280 -40
rect 240 -122 1280 -120
rect 240 -238 980 -122
rect 1160 -238 1280 -122
rect 240 -240 1280 -238
rect 240 -320 440 -240
rect 840 -340 1280 -240
rect 2060 -1580 2140 100
rect 2300 -1580 2440 1556
rect 3460 1757 3780 1780
rect 4665 1763 6220 1806
rect 4976 1760 6220 1763
rect 3460 1723 3567 1757
rect 3601 1723 3639 1757
rect 3673 1723 3780 1757
rect 3460 1260 3780 1723
rect 6800 1757 7080 1780
rect 6800 1723 6897 1757
rect 6931 1723 6969 1757
rect 7003 1723 7080 1757
rect 6800 1500 7080 1723
rect 9301 1504 9741 1579
rect 8749 1500 9741 1504
rect 6800 1497 9741 1500
rect 6800 1381 9441 1497
rect 9621 1381 9741 1497
rect 6800 1361 9741 1381
rect 6800 1360 8263 1361
rect 4860 1320 5840 1340
rect 4860 1280 4920 1320
rect 5080 1280 5840 1320
rect 4860 1260 5840 1280
rect 3500 1098 3700 1260
rect 2853 1020 3700 1098
rect 2853 1019 3697 1020
rect 2859 720 2930 1019
rect 4860 857 5180 1260
rect 4860 823 4967 857
rect 5001 823 5039 857
rect 5073 823 5180 857
rect 4860 800 5180 823
rect 2859 686 2875 720
rect 2909 686 2930 720
rect 2859 654 2930 686
rect 5360 726 5440 760
rect 5360 674 5374 726
rect 5426 674 5440 726
rect 5360 620 5440 674
rect 3680 577 3760 600
rect 3680 543 3703 577
rect 3737 543 3760 577
rect 3680 500 3760 543
rect 3620 477 3800 500
rect 3620 443 3693 477
rect 3727 443 3800 477
rect 3620 420 3800 443
rect 3700 -500 3740 420
rect 5720 217 5840 1260
rect 6800 1197 7080 1360
rect 9170 1359 9741 1361
rect 9301 1279 9741 1359
rect 6800 1163 6897 1197
rect 6931 1163 6969 1197
rect 7003 1163 7080 1197
rect 6800 1140 7080 1163
rect 6100 1066 6220 1080
rect 6100 1014 6134 1066
rect 6186 1014 6220 1066
rect 6100 1000 6220 1014
rect 6560 937 6760 960
rect 6560 903 6607 937
rect 6641 903 6679 937
rect 6713 903 6760 937
rect 6560 880 6760 903
rect 7460 937 7680 960
rect 7460 903 7527 937
rect 7561 903 7599 937
rect 7633 903 7680 937
rect 7460 880 7680 903
rect 6640 840 6680 880
rect 6600 817 6720 840
rect 6600 783 6643 817
rect 6677 783 6720 817
rect 6600 760 6720 783
rect 5720 183 5763 217
rect 5797 183 5840 217
rect 5720 160 5840 183
rect 6640 -500 6680 760
rect 7560 -500 7600 880
rect 2760 -577 5600 -500
rect 2760 -597 4623 -577
rect 2760 -631 2783 -597
rect 2817 -631 3703 -597
rect 3737 -611 4623 -597
rect 4657 -611 5543 -577
rect 5577 -611 5600 -577
rect 3737 -631 5600 -611
rect 2760 -649 5600 -631
rect 2760 -669 4623 -649
rect 2760 -703 2783 -669
rect 2817 -703 3703 -669
rect 3737 -683 4623 -669
rect 4657 -683 5543 -649
rect 5577 -683 5600 -649
rect 3737 -703 5600 -683
rect 2760 -760 5600 -703
rect 6620 -567 9460 -500
rect 6620 -587 8483 -567
rect 6620 -621 6643 -587
rect 6677 -621 7563 -587
rect 7597 -601 8483 -587
rect 8517 -601 9403 -567
rect 9437 -601 9460 -567
rect 7597 -621 9460 -601
rect 6620 -639 9460 -621
rect 6620 -659 8483 -639
rect 6620 -693 6643 -659
rect 6677 -693 7563 -659
rect 7597 -673 8483 -659
rect 8517 -673 9403 -639
rect 9437 -673 9460 -639
rect 7597 -693 9460 -673
rect 6620 -760 9460 -693
rect 6620 -780 6700 -760
rect 3220 -1083 10920 -1020
rect 3220 -1093 9963 -1083
rect 3220 -1127 3243 -1093
rect 3277 -1127 4163 -1093
rect 4197 -1127 5083 -1093
rect 5117 -1127 6003 -1093
rect 6037 -1103 7103 -1093
rect 6037 -1127 6103 -1103
rect 3220 -1137 6103 -1127
rect 6137 -1127 7103 -1103
rect 7137 -1127 8023 -1093
rect 8057 -1127 8943 -1093
rect 8977 -1127 9863 -1093
rect 9897 -1117 9963 -1093
rect 9997 -1117 10920 -1083
rect 9897 -1127 10920 -1117
rect 6137 -1137 10920 -1127
rect 3220 -1180 10920 -1137
rect 2840 -1303 9840 -1260
rect 2840 -1337 2987 -1303
rect 3021 -1337 3059 -1303
rect 3093 -1337 3467 -1303
rect 3501 -1337 3539 -1303
rect 3573 -1337 3907 -1303
rect 3941 -1337 3979 -1303
rect 4013 -1337 4367 -1303
rect 4401 -1337 4439 -1303
rect 4473 -1337 4847 -1303
rect 4881 -1337 4919 -1303
rect 4953 -1337 5287 -1303
rect 5321 -1337 5359 -1303
rect 5393 -1337 5747 -1303
rect 5781 -1337 5819 -1303
rect 5853 -1337 6847 -1303
rect 6881 -1337 6919 -1303
rect 6953 -1337 7327 -1303
rect 7361 -1337 7399 -1303
rect 7433 -1337 7767 -1303
rect 7801 -1337 7839 -1303
rect 7873 -1337 8227 -1303
rect 8261 -1337 8299 -1303
rect 8333 -1337 8687 -1303
rect 8721 -1337 8759 -1303
rect 8793 -1337 9167 -1303
rect 9201 -1337 9239 -1303
rect 9273 -1337 9627 -1303
rect 9661 -1337 9699 -1303
rect 9733 -1337 9840 -1303
rect 2840 -1360 9840 -1337
rect 2060 -1740 4000 -1580
rect 3820 -2180 4000 -1740
rect -1800 -2263 2860 -2200
rect -1800 -2297 -1777 -2263
rect -1743 -2297 -857 -2263
rect -823 -2297 63 -2263
rect 97 -2297 983 -2263
rect 1017 -2297 1903 -2263
rect 1937 -2297 2803 -2263
rect 2837 -2297 2860 -2263
rect -1800 -2380 2860 -2297
rect 3820 -2293 10520 -2180
rect 3820 -2327 4963 -2293
rect 4997 -2327 5883 -2293
rect 5917 -2327 6803 -2293
rect 6837 -2327 7723 -2293
rect 7757 -2327 8643 -2293
rect 8677 -2313 10520 -2293
rect 8677 -2327 9543 -2313
rect 3820 -2347 9543 -2327
rect 9577 -2347 10463 -2313
rect 10497 -2347 10520 -2313
rect 3820 -2440 10520 -2347
rect -2080 -3100 -2000 -3080
rect -1920 -3100 -1840 -3080
rect 10720 -3100 10920 -1180
rect -2200 -3107 10920 -3100
rect -2200 -3141 -2057 -3107
rect -2023 -3134 10920 -3107
rect -2023 -3141 3884 -3134
rect -2200 -3143 3884 -3141
rect 3936 -3143 10920 -3134
rect -2200 -3177 -2177 -3143
rect -2143 -3153 -1317 -3143
rect -2143 -3177 -1877 -3153
rect -2200 -3179 -1877 -3177
rect -3520 -3262 -3080 -3180
rect -2200 -3213 -2057 -3179
rect -2023 -3187 -1877 -3179
rect -1843 -3177 -1317 -3153
rect -1283 -3177 -397 -3143
rect -363 -3177 523 -3143
rect 557 -3177 1443 -3143
rect 1477 -3177 2343 -3143
rect 2377 -3177 3884 -3143
rect 3936 -3177 4863 -3143
rect 4897 -3177 5423 -3143
rect 5457 -3177 6343 -3143
rect 6377 -3177 7263 -3143
rect 7297 -3177 8163 -3143
rect 8197 -3177 9083 -3143
rect 9117 -3177 10003 -3143
rect 10037 -3177 10920 -3143
rect -1843 -3186 3884 -3177
rect 3936 -3186 10920 -3177
rect -1843 -3187 10920 -3186
rect -2023 -3213 10920 -3187
rect -2200 -3220 10920 -3213
rect -2080 -3240 -2000 -3220
rect -1920 -3240 -1820 -3220
rect -3520 -3378 -3380 -3262
rect -3200 -3280 -3080 -3262
rect -3200 -3333 -2580 -3280
rect -3200 -3367 -2637 -3333
rect -2603 -3367 -2580 -3333
rect -3200 -3378 -2580 -3367
rect -3520 -3420 -2580 -3378
rect -3520 -3480 -3080 -3420
rect -2660 -3443 10460 -3420
rect -2660 -3477 -2463 -3443
rect -2429 -3477 -2391 -3443
rect -2357 -3477 -1583 -3443
rect -1549 -3477 -1511 -3443
rect -1477 -3477 -1123 -3443
rect -1089 -3477 -1051 -3443
rect -1017 -3477 -663 -3443
rect -629 -3477 -591 -3443
rect -557 -3477 -243 -3443
rect -209 -3477 -171 -3443
rect -137 -3477 237 -3443
rect 271 -3477 309 -3443
rect 343 -3477 697 -3443
rect 731 -3477 769 -3443
rect 803 -3477 1157 -3443
rect 1191 -3477 1229 -3443
rect 1263 -3477 1617 -3443
rect 1651 -3477 1689 -3443
rect 1723 -3477 2077 -3443
rect 2111 -3477 2149 -3443
rect 2183 -3477 2557 -3443
rect 2591 -3477 2629 -3443
rect 2663 -3477 5167 -3443
rect 5201 -3477 5239 -3443
rect 5273 -3477 5627 -3443
rect 5661 -3477 5699 -3443
rect 5733 -3477 6087 -3443
rect 6121 -3477 6159 -3443
rect 6193 -3477 6547 -3443
rect 6581 -3477 6619 -3443
rect 6653 -3477 7007 -3443
rect 7041 -3477 7079 -3443
rect 7113 -3477 7447 -3443
rect 7481 -3477 7519 -3443
rect 7553 -3477 7907 -3443
rect 7941 -3477 7979 -3443
rect 8013 -3477 8367 -3443
rect 8401 -3477 8439 -3443
rect 8473 -3477 8847 -3443
rect 8881 -3477 8919 -3443
rect 8953 -3477 9287 -3443
rect 9321 -3477 9359 -3443
rect 9393 -3477 9747 -3443
rect 9781 -3477 9819 -3443
rect 9853 -3477 10207 -3443
rect 10241 -3477 10279 -3443
rect 10313 -3477 10460 -3443
rect -2660 -3500 10460 -3477
rect -2780 -3734 10640 -3620
rect -2780 -3743 3874 -3734
rect 3926 -3743 10640 -3734
rect -2780 -3777 -2639 -3743
rect -2605 -3777 -2567 -3743
rect -2533 -3777 -2495 -3743
rect -2461 -3777 -2423 -3743
rect -2389 -3777 -2351 -3743
rect -2317 -3777 -2279 -3743
rect -2245 -3777 -2207 -3743
rect -2173 -3777 -2135 -3743
rect -2101 -3777 -2063 -3743
rect -2029 -3777 -1991 -3743
rect -1957 -3777 -1919 -3743
rect -1885 -3777 -1847 -3743
rect -1813 -3777 -1775 -3743
rect -1741 -3777 -1703 -3743
rect -1669 -3777 -1631 -3743
rect -1597 -3777 -1559 -3743
rect -1525 -3777 -1487 -3743
rect -1453 -3777 -1415 -3743
rect -1381 -3777 -1343 -3743
rect -1309 -3777 -1271 -3743
rect -1237 -3777 -1199 -3743
rect -1165 -3777 -1127 -3743
rect -1093 -3777 -1055 -3743
rect -1021 -3777 -983 -3743
rect -949 -3777 -911 -3743
rect -877 -3777 -839 -3743
rect -805 -3777 -767 -3743
rect -733 -3777 -695 -3743
rect -661 -3777 -623 -3743
rect -589 -3777 -551 -3743
rect -517 -3777 -479 -3743
rect -445 -3777 -407 -3743
rect -373 -3777 -335 -3743
rect -301 -3777 -263 -3743
rect -229 -3777 -191 -3743
rect -157 -3777 -119 -3743
rect -85 -3777 -47 -3743
rect -13 -3777 25 -3743
rect 59 -3777 97 -3743
rect 131 -3777 169 -3743
rect 203 -3777 241 -3743
rect 275 -3777 313 -3743
rect 347 -3777 385 -3743
rect 419 -3777 457 -3743
rect 491 -3777 529 -3743
rect 563 -3777 601 -3743
rect 635 -3777 673 -3743
rect 707 -3777 745 -3743
rect 779 -3777 817 -3743
rect 851 -3777 889 -3743
rect 923 -3777 961 -3743
rect 995 -3777 1033 -3743
rect 1067 -3777 1105 -3743
rect 1139 -3777 1177 -3743
rect 1211 -3777 1249 -3743
rect 1283 -3777 1321 -3743
rect 1355 -3777 1393 -3743
rect 1427 -3777 1465 -3743
rect 1499 -3777 1537 -3743
rect 1571 -3777 1609 -3743
rect 1643 -3777 1681 -3743
rect 1715 -3777 1753 -3743
rect 1787 -3777 1825 -3743
rect 1859 -3777 1897 -3743
rect 1931 -3777 1969 -3743
rect 2003 -3777 2041 -3743
rect 2075 -3777 2113 -3743
rect 2147 -3777 2185 -3743
rect 2219 -3777 2257 -3743
rect 2291 -3777 2329 -3743
rect 2363 -3777 2401 -3743
rect 2435 -3777 2473 -3743
rect 2507 -3777 2545 -3743
rect 2579 -3777 2617 -3743
rect 2651 -3777 2689 -3743
rect 2723 -3777 2761 -3743
rect 2795 -3777 2833 -3743
rect 2867 -3777 2905 -3743
rect 2939 -3777 2977 -3743
rect 3011 -3777 3049 -3743
rect 3083 -3777 3121 -3743
rect 3155 -3777 3193 -3743
rect 3227 -3777 3265 -3743
rect 3299 -3777 3337 -3743
rect 3371 -3777 3409 -3743
rect 3443 -3777 3481 -3743
rect 3515 -3777 3553 -3743
rect 3587 -3777 3625 -3743
rect 3659 -3777 3697 -3743
rect 3731 -3777 3769 -3743
rect 3803 -3777 3841 -3743
rect 3947 -3777 3985 -3743
rect 4019 -3777 4057 -3743
rect 4091 -3777 4129 -3743
rect 4163 -3777 4201 -3743
rect 4235 -3777 4273 -3743
rect 4307 -3777 4345 -3743
rect 4379 -3777 4417 -3743
rect 4451 -3777 4489 -3743
rect 4523 -3777 4561 -3743
rect 4595 -3777 4633 -3743
rect 4667 -3777 4705 -3743
rect 4739 -3777 4777 -3743
rect 4811 -3777 4849 -3743
rect 4883 -3777 4921 -3743
rect 4955 -3777 4993 -3743
rect 5027 -3777 5065 -3743
rect 5099 -3777 5137 -3743
rect 5171 -3777 5209 -3743
rect 5243 -3777 5281 -3743
rect 5315 -3777 5353 -3743
rect 5387 -3777 5425 -3743
rect 5459 -3777 5497 -3743
rect 5531 -3777 5569 -3743
rect 5603 -3777 5641 -3743
rect 5675 -3777 5713 -3743
rect 5747 -3777 5785 -3743
rect 5819 -3777 5857 -3743
rect 5891 -3777 5929 -3743
rect 5963 -3777 6001 -3743
rect 6035 -3777 6073 -3743
rect 6107 -3777 6145 -3743
rect 6179 -3777 6217 -3743
rect 6251 -3777 6289 -3743
rect 6323 -3777 6361 -3743
rect 6395 -3777 6433 -3743
rect 6467 -3777 6505 -3743
rect 6539 -3777 6577 -3743
rect 6611 -3777 6649 -3743
rect 6683 -3777 6721 -3743
rect 6755 -3777 6793 -3743
rect 6827 -3777 6865 -3743
rect 6899 -3777 6937 -3743
rect 6971 -3777 7009 -3743
rect 7043 -3777 7081 -3743
rect 7115 -3777 7153 -3743
rect 7187 -3777 7225 -3743
rect 7259 -3777 7297 -3743
rect 7331 -3777 7369 -3743
rect 7403 -3777 7441 -3743
rect 7475 -3777 7513 -3743
rect 7547 -3777 7585 -3743
rect 7619 -3777 7657 -3743
rect 7691 -3777 7729 -3743
rect 7763 -3777 7801 -3743
rect 7835 -3777 7873 -3743
rect 7907 -3777 7945 -3743
rect 7979 -3777 8017 -3743
rect 8051 -3777 8089 -3743
rect 8123 -3777 8161 -3743
rect 8195 -3777 8233 -3743
rect 8267 -3777 8305 -3743
rect 8339 -3777 8377 -3743
rect 8411 -3777 8449 -3743
rect 8483 -3777 8521 -3743
rect 8555 -3777 8593 -3743
rect 8627 -3777 8665 -3743
rect 8699 -3777 8737 -3743
rect 8771 -3777 8809 -3743
rect 8843 -3777 8881 -3743
rect 8915 -3777 8953 -3743
rect 8987 -3777 9025 -3743
rect 9059 -3777 9097 -3743
rect 9131 -3777 9169 -3743
rect 9203 -3777 9241 -3743
rect 9275 -3777 9313 -3743
rect 9347 -3777 9385 -3743
rect 9419 -3777 9457 -3743
rect 9491 -3777 9529 -3743
rect 9563 -3777 9601 -3743
rect 9635 -3777 9673 -3743
rect 9707 -3777 9745 -3743
rect 9779 -3777 9817 -3743
rect 9851 -3777 9889 -3743
rect 9923 -3777 9961 -3743
rect 9995 -3777 10033 -3743
rect 10067 -3777 10105 -3743
rect 10139 -3777 10177 -3743
rect 10211 -3777 10249 -3743
rect 10283 -3777 10321 -3743
rect 10355 -3777 10393 -3743
rect 10427 -3777 10465 -3743
rect 10499 -3777 10640 -3743
rect -2780 -3786 3874 -3777
rect 3926 -3786 10640 -3777
rect -2780 -3880 10640 -3786
rect -1820 -4060 -1700 -3880
rect -2000 -4142 -1560 -4060
rect -2000 -4258 -1860 -4142
rect -1680 -4258 -1560 -4142
rect -2000 -4360 -1560 -4258
<< via1 >>
rect -3340 4222 -3160 4338
rect -1296 2337 -1244 2346
rect -1296 2303 -1277 2337
rect -1277 2303 -1244 2337
rect -1296 2294 -1244 2303
rect 3990 2303 4027 2336
rect 4027 2303 4042 2336
rect 4054 2303 4061 2336
rect 4061 2303 4099 2336
rect 4099 2303 4106 2336
rect 4118 2303 4133 2336
rect 4133 2303 4170 2336
rect 3990 2284 4042 2303
rect 4054 2284 4106 2303
rect 4118 2284 4170 2303
rect 6840 2297 7020 2338
rect 6840 2263 6913 2297
rect 6913 2263 6947 2297
rect 6947 2263 7020 2297
rect 6840 2222 7020 2263
rect 990 833 1170 838
rect 990 799 1063 833
rect 1063 799 1097 833
rect 1097 799 1170 833
rect 990 761 1170 799
rect 990 727 1063 761
rect 1063 727 1097 761
rect 1097 727 1170 761
rect 990 722 1170 727
rect -780 -198 -600 -82
rect 980 -238 1160 -122
rect 9441 1381 9621 1497
rect 5374 717 5426 726
rect 5374 683 5383 717
rect 5383 683 5417 717
rect 5417 683 5426 717
rect 5374 674 5426 683
rect 6134 1057 6186 1066
rect 6134 1023 6143 1057
rect 6143 1023 6177 1057
rect 6177 1023 6186 1057
rect 6134 1014 6186 1023
rect 3884 -3143 3936 -3134
rect 3884 -3177 3893 -3143
rect 3893 -3177 3927 -3143
rect 3927 -3177 3936 -3143
rect 3884 -3186 3936 -3177
rect -3380 -3378 -3200 -3262
rect 3874 -3743 3926 -3734
rect 3874 -3777 3875 -3743
rect 3875 -3777 3913 -3743
rect 3913 -3777 3926 -3743
rect 3874 -3786 3926 -3777
rect -1860 -4258 -1680 -4142
<< metal2 >>
rect -3500 4348 -3000 4460
rect -3500 4212 -3358 4348
rect -3142 4212 -3000 4348
rect -3500 4080 -3000 4212
rect 246 2380 644 2385
rect 960 2380 1728 2383
rect -1340 2346 4200 2380
rect -1340 2294 -1296 2346
rect -1244 2336 4200 2346
rect -1244 2294 3990 2336
rect -1340 2284 3990 2294
rect 4042 2284 4054 2336
rect 4106 2284 4118 2336
rect 4170 2284 4200 2336
rect -1340 2223 4200 2284
rect -1340 2220 319 2223
rect 553 2220 4200 2223
rect 5680 2338 7100 2380
rect 5680 2222 6840 2338
rect 7020 2222 7100 2338
rect 5680 2200 7100 2222
rect 5680 1540 5900 2200
rect 980 1340 5900 1540
rect 9281 1507 9781 1619
rect 9281 1371 9423 1507
rect 9639 1371 9781 1507
rect 980 838 1180 1340
rect 9281 1239 9781 1371
rect 6100 1066 6220 1120
rect 6100 1014 6134 1066
rect 6186 1014 6220 1066
rect 6100 920 6220 1014
rect 980 722 990 838
rect 1170 722 1180 838
rect 6120 780 6200 920
rect 980 680 1180 722
rect 5340 726 6200 780
rect 5340 674 5374 726
rect 5426 674 6200 726
rect 5340 620 6200 674
rect -940 -72 -440 40
rect -940 -208 -798 -72
rect -582 -208 -440 -72
rect -940 -340 -440 -208
rect 820 -112 1320 0
rect 820 -248 962 -112
rect 1178 -248 1320 -112
rect 820 -380 1320 -248
rect 3840 -3134 3980 -3100
rect -3540 -3252 -3040 -3140
rect -3540 -3388 -3398 -3252
rect -3182 -3388 -3040 -3252
rect -3540 -3520 -3040 -3388
rect 3840 -3186 3884 -3134
rect 3936 -3186 3980 -3134
rect 3840 -3734 3980 -3186
rect 3840 -3786 3874 -3734
rect 3926 -3786 3980 -3734
rect 3840 -3840 3980 -3786
rect -2020 -4132 -1520 -4020
rect -2020 -4268 -1878 -4132
rect -1662 -4268 -1520 -4132
rect -2020 -4400 -1520 -4268
<< via2 >>
rect -3358 4338 -3142 4348
rect -3358 4222 -3340 4338
rect -3340 4222 -3160 4338
rect -3160 4222 -3142 4338
rect -3358 4212 -3142 4222
rect 9423 1497 9639 1507
rect 9423 1381 9441 1497
rect 9441 1381 9621 1497
rect 9621 1381 9639 1497
rect 9423 1371 9639 1381
rect -798 -82 -582 -72
rect -798 -198 -780 -82
rect -780 -198 -600 -82
rect -600 -198 -582 -82
rect -798 -208 -582 -198
rect 962 -122 1178 -112
rect 962 -238 980 -122
rect 980 -238 1160 -122
rect 1160 -238 1178 -122
rect 962 -248 1178 -238
rect -3398 -3262 -3182 -3252
rect -3398 -3378 -3380 -3262
rect -3380 -3378 -3200 -3262
rect -3200 -3378 -3182 -3262
rect -3398 -3388 -3182 -3378
rect -1878 -4142 -1662 -4132
rect -1878 -4258 -1860 -4142
rect -1860 -4258 -1680 -4142
rect -1680 -4258 -1662 -4142
rect -1878 -4268 -1662 -4258
<< metal3 >>
rect -3520 4348 -2980 4460
rect -3520 4342 -3358 4348
rect -3142 4342 -2980 4348
rect -3520 4198 -3362 4342
rect -3138 4198 -2980 4342
rect -3520 4060 -2980 4198
rect 9261 1507 9801 1619
rect 9261 1501 9423 1507
rect 9639 1501 9801 1507
rect 9261 1357 9419 1501
rect 9643 1357 9801 1501
rect 9261 1219 9801 1357
rect -960 -72 -420 40
rect -960 -78 -798 -72
rect -582 -78 -420 -72
rect -960 -222 -802 -78
rect -578 -222 -420 -78
rect -960 -360 -420 -222
rect 800 -112 1340 0
rect 800 -118 962 -112
rect 1178 -118 1340 -112
rect 800 -262 958 -118
rect 1182 -262 1340 -118
rect 800 -400 1340 -262
rect -3560 -3252 -3020 -3140
rect -3560 -3258 -3398 -3252
rect -3182 -3258 -3020 -3252
rect -3560 -3402 -3402 -3258
rect -3178 -3402 -3020 -3258
rect -3560 -3540 -3020 -3402
rect -2040 -4132 -1500 -4020
rect -2040 -4138 -1878 -4132
rect -1662 -4138 -1500 -4132
rect -2040 -4282 -1882 -4138
rect -1658 -4282 -1500 -4138
rect -2040 -4420 -1500 -4282
<< via3 >>
rect -3362 4212 -3358 4342
rect -3358 4212 -3142 4342
rect -3142 4212 -3138 4342
rect -3362 4198 -3138 4212
rect 9419 1371 9423 1501
rect 9423 1371 9639 1501
rect 9639 1371 9643 1501
rect 9419 1357 9643 1371
rect -802 -208 -798 -78
rect -798 -208 -582 -78
rect -582 -208 -578 -78
rect -802 -222 -578 -208
rect 958 -248 962 -118
rect 962 -248 1178 -118
rect 1178 -248 1182 -118
rect 958 -262 1182 -248
rect -3402 -3388 -3398 -3258
rect -3398 -3388 -3182 -3258
rect -3182 -3388 -3178 -3258
rect -3402 -3402 -3178 -3388
rect -1882 -4268 -1878 -4138
rect -1878 -4268 -1662 -4138
rect -1662 -4268 -1658 -4138
rect -1882 -4282 -1658 -4268
<< metal4 >>
rect -3540 4388 -2940 4480
rect -3540 4152 -3368 4388
rect -3132 4152 -2940 4388
rect -3540 4040 -2940 4152
rect 9241 1547 9841 1639
rect 9241 1311 9413 1547
rect 9649 1311 9841 1547
rect 9241 1199 9841 1311
rect -980 -32 -380 60
rect -980 -268 -808 -32
rect -572 -268 -380 -32
rect -980 -380 -380 -268
rect 780 -72 1380 20
rect 780 -308 952 -72
rect 1188 -308 1380 -72
rect 780 -420 1380 -308
rect -3580 -3212 -2980 -3120
rect -3580 -3448 -3408 -3212
rect -3172 -3448 -2980 -3212
rect -3580 -3560 -2980 -3448
rect -2060 -4092 -1460 -4000
rect -2060 -4328 -1888 -4092
rect -1652 -4328 -1460 -4092
rect -2060 -4440 -1460 -4328
<< via4 >>
rect -3368 4342 -3132 4388
rect -3368 4198 -3362 4342
rect -3362 4198 -3138 4342
rect -3138 4198 -3132 4342
rect -3368 4152 -3132 4198
rect 9413 1501 9649 1547
rect 9413 1357 9419 1501
rect 9419 1357 9643 1501
rect 9643 1357 9649 1501
rect 9413 1311 9649 1357
rect -808 -78 -572 -32
rect -808 -222 -802 -78
rect -802 -222 -578 -78
rect -578 -222 -572 -78
rect -808 -268 -572 -222
rect 952 -118 1188 -72
rect 952 -262 958 -118
rect 958 -262 1182 -118
rect 1182 -262 1188 -118
rect 952 -308 1188 -262
rect -3408 -3258 -3172 -3212
rect -3408 -3402 -3402 -3258
rect -3402 -3402 -3178 -3258
rect -3178 -3402 -3172 -3258
rect -3408 -3448 -3172 -3402
rect -1888 -4138 -1652 -4092
rect -1888 -4282 -1882 -4138
rect -1882 -4282 -1658 -4138
rect -1658 -4282 -1652 -4138
rect -1888 -4328 -1652 -4282
<< metal5 >>
rect -3560 4388 -2920 4500
rect -3560 4152 -3368 4388
rect -3132 4152 -2920 4388
rect -3560 4020 -2920 4152
rect 9221 1547 9861 1659
rect 9221 1311 9413 1547
rect 9649 1311 9861 1547
rect 9221 1179 9861 1311
rect -1000 -32 -360 80
rect -1000 -268 -808 -32
rect -572 -268 -360 -32
rect -1000 -400 -360 -268
rect 760 -72 1400 40
rect 760 -308 952 -72
rect 1188 -308 1400 -72
rect 760 -440 1400 -308
rect -3600 -3212 -2960 -3100
rect -3600 -3448 -3408 -3212
rect -3172 -3448 -2960 -3212
rect -3600 -3580 -2960 -3448
rect -2080 -4092 -1440 -3980
rect -2080 -4328 -1888 -4092
rect -1652 -4328 -1440 -4092
rect -2080 -4460 -1440 -4328
use sky130_fd_pr__nfet_01v8_lvt_4oweb9  sky130_fd_pr__nfet_01v8_lvt_4oweb9_0
timestamp 1611881054
transform 1 0 -2384 0 1 -2710
box -360 -874 360 874
use sky130_fd_pr__nfet_01v8_lvt_9YHVJG  sky130_fd_pr__nfet_01v8_lvt_9YHVJG_0
timestamp 1611881054
transform 1 0 535 0 1 -2709
box -2421 -874 2421 874
use sky130_fd_pr__nfet_01v8_lvt_6vyjkp  sky130_fd_pr__nfet_01v8_lvt_6vyjkp_0
timestamp 1611881054
transform 1 0 7735 0 1 -2710
box -2879 -874 2879 874
use sky130_fd_pr__res_high_po_0p35_rfxuin  sky130_fd_pr__res_high_po_0p35_rfxuin_0
timestamp 1611881054
transform 1 0 2101 0 1 689
box -165 -693 165 693
use sky130_fd_pr__nfet_01v8_im9uye  sky130_fd_pr__nfet_01v8_im9uye_0
timestamp 1611881054
transform 1 0 4410 0 1 -570
box -1734 -874 1734 874
use sky130_fd_pr__nfet_01v8_lvt_2ZZGCN  sky130_fd_pr__nfet_01v8_lvt_2ZZGCN_1
timestamp 1611881054
transform 1 0 -1549 0 1 337
box -360 -374 360 374
use sky130_fd_pr__nfet_01v8_lvt_2ZZGCN  sky130_fd_pr__nfet_01v8_lvt_2ZZGCN_0
timestamp 1611881054
transform 1 0 328 0 1 403
box -360 -374 360 374
use sky130_fd_pr__nfet_01v8_cvwdxd  sky130_fd_pr__nfet_01v8_cvwdxd_0
timestamp 1611881054
transform 1 0 8270 0 1 -570
box -1734 -874 1734 874
use sky130_fd_pr__pfet_01v8_lvt_M62V36  sky130_fd_pr__pfet_01v8_lvt_M62V36_0
timestamp 1611881054
transform 0 1 1249 -1 0 1865
box -296 -1219 296 1219
use sky130_fd_pr__nfet_01v8_lvt_VCXKU2  sky130_fd_pr__nfet_01v8_lvt_VCXKU2_1
timestamp 1611881054
transform 0 1 4154 -1 0 706
box -260 -1374 260 1374
use sky130_fd_pr__nfet_01v8_lvt_VCXKU2  sky130_fd_pr__nfet_01v8_lvt_VCXKU2_0
timestamp 1611881054
transform 0 1 7427 -1 0 1038
box -260 -1374 260 1374
use sky130_fd_pr__pfet_01v8_lvt_RAZ4RL  sky130_fd_pr__pfet_01v8_lvt_RAZ4RL_1
timestamp 1611881054
transform 0 1 6843 -1 0 1878
box -296 -819 296 819
use sky130_fd_pr__pfet_01v8_lvt_RAZ4RL  sky130_fd_pr__pfet_01v8_lvt_RAZ4RL_0
timestamp 1611881054
transform 0 1 4042 -1 0 1878
box -296 -819 296 819
use sky130_fd_pr__res_xhigh_po_0p35_6FRE74  sky130_fd_pr__res_xhigh_po_0p35_6FRE74_0
timestamp 1611881054
transform 0 1 4284 -1 0 1301
box -165 -1020 165 1020
use sky130_fd_pr__pfet_01v8_NLQV3P  sky130_fd_pr__pfet_01v8_NLQV3P_1
timestamp 1611881054
transform 1 0 -953 0 1 3347
box -1770 -919 1770 919
use sky130_fd_pr__pfet_01v8_NLQV3P  sky130_fd_pr__pfet_01v8_NLQV3P_0
timestamp 1611881054
transform 1 0 4313 0 1 3349
box -1770 -919 1770 919
use sky130_fd_pr__pfet_01v8_U5BVXJ  sky130_fd_pr__pfet_01v8_U5BVXJ_0
timestamp 1611881054
transform 1 0 9337 0 1 3351
box -1770 -919 1770 919
<< labels >>
rlabel metal1 s -2600 4260 -2540 4320 4 VDD
port 1 nsew
rlabel metal1 s 6860 1360 7060 1480 4 VOUT
port 2 nsew
rlabel metal1 s -1580 -220 -1480 -120 4 VINP
port 3 nsew
rlabel metal1 s 300 -240 380 -120 4 VINN
port 4 nsew
rlabel metal1 s -2880 -3380 -2800 -3320 4 IBP
port 5 nsew
rlabel metal1 s -1800 -3840 -1700 -3680 4 VSS
port 6 nsew
<< end >>
