magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< poly >>
rect 1386 -298 1482 -238
rect 1988 -244 2068 -238
rect 1988 -292 2078 -244
rect 1988 -298 2068 -292
rect 2084 -298 2114 -290
<< locali >>
rect 186 2022 3244 2060
rect 186 1988 261 2022
rect 295 2020 2477 2022
rect 295 2016 2037 2020
rect 295 1988 571 2016
rect 186 1982 571 1988
rect 605 2010 1363 2016
rect 605 1982 887 2010
rect 186 1976 887 1982
rect 921 1982 1363 2010
rect 1397 1986 2037 2016
rect 2071 1988 2477 2020
rect 2511 1988 2771 2022
rect 2805 1988 3073 2022
rect 3107 1988 3244 2022
rect 2071 1986 3244 1988
rect 1397 1982 3244 1986
rect 921 1976 3244 1982
rect 186 1936 3244 1976
rect 113 1578 183 1597
rect 113 1544 131 1578
rect 165 1544 183 1578
rect 113 1506 183 1544
rect 113 1472 131 1506
rect 165 1472 183 1506
rect 113 1434 183 1472
rect 113 1400 131 1434
rect 165 1400 183 1434
rect 113 1362 183 1400
rect 113 1328 131 1362
rect 165 1328 183 1362
rect 113 1290 183 1328
rect 113 1256 131 1290
rect 165 1256 183 1290
rect 113 1218 183 1256
rect 113 1184 131 1218
rect 165 1184 183 1218
rect 113 1165 183 1184
rect 431 1578 501 1597
rect 431 1544 449 1578
rect 483 1544 501 1578
rect 431 1506 501 1544
rect 431 1472 449 1506
rect 483 1472 501 1506
rect 431 1434 501 1472
rect 431 1400 449 1434
rect 483 1400 501 1434
rect 431 1362 501 1400
rect 431 1328 449 1362
rect 483 1328 501 1362
rect 431 1290 501 1328
rect 431 1256 449 1290
rect 483 1256 501 1290
rect 431 1218 501 1256
rect 431 1184 449 1218
rect 483 1184 501 1218
rect 431 1165 501 1184
rect 749 1578 819 1597
rect 749 1544 767 1578
rect 801 1544 819 1578
rect 749 1506 819 1544
rect 749 1472 767 1506
rect 801 1472 819 1506
rect 749 1434 819 1472
rect 749 1400 767 1434
rect 801 1400 819 1434
rect 749 1362 819 1400
rect 749 1328 767 1362
rect 801 1328 819 1362
rect 749 1290 819 1328
rect 749 1256 767 1290
rect 801 1256 819 1290
rect 749 1218 819 1256
rect 749 1184 767 1218
rect 801 1184 819 1218
rect 749 1165 819 1184
rect 1067 1578 1137 1597
rect 1067 1544 1085 1578
rect 1119 1544 1137 1578
rect 1067 1506 1137 1544
rect 1067 1472 1085 1506
rect 1119 1472 1137 1506
rect 1067 1434 1137 1472
rect 1067 1400 1085 1434
rect 1119 1400 1137 1434
rect 1067 1362 1137 1400
rect 1067 1328 1085 1362
rect 1119 1328 1137 1362
rect 1067 1290 1137 1328
rect 1067 1256 1085 1290
rect 1119 1256 1137 1290
rect 1067 1218 1137 1256
rect 1067 1184 1085 1218
rect 1119 1184 1137 1218
rect 1067 1165 1137 1184
rect 2316 1573 2386 1592
rect 2316 1539 2334 1573
rect 2368 1539 2386 1573
rect 2316 1501 2386 1539
rect 2316 1467 2334 1501
rect 2368 1467 2386 1501
rect 2316 1429 2386 1467
rect 2316 1395 2334 1429
rect 2368 1395 2386 1429
rect 2316 1357 2386 1395
rect 2316 1323 2334 1357
rect 2368 1323 2386 1357
rect 2316 1285 2386 1323
rect 2316 1251 2334 1285
rect 2368 1251 2386 1285
rect 2316 1213 2386 1251
rect 2316 1179 2334 1213
rect 2368 1179 2386 1213
rect 2316 1160 2386 1179
rect 2634 1573 2704 1592
rect 2634 1539 2652 1573
rect 2686 1539 2704 1573
rect 2634 1501 2704 1539
rect 2634 1467 2652 1501
rect 2686 1467 2704 1501
rect 2634 1429 2704 1467
rect 2634 1395 2652 1429
rect 2686 1395 2704 1429
rect 2634 1357 2704 1395
rect 2634 1323 2652 1357
rect 2686 1323 2704 1357
rect 2634 1285 2704 1323
rect 2634 1251 2652 1285
rect 2686 1251 2704 1285
rect 2634 1213 2704 1251
rect 2634 1179 2652 1213
rect 2686 1179 2704 1213
rect 2634 1160 2704 1179
rect 2952 1573 3022 1592
rect 2952 1539 2970 1573
rect 3004 1539 3022 1573
rect 2952 1501 3022 1539
rect 2952 1467 2970 1501
rect 3004 1467 3022 1501
rect 2952 1429 3022 1467
rect 2952 1395 2970 1429
rect 3004 1395 3022 1429
rect 2952 1357 3022 1395
rect 2952 1323 2970 1357
rect 3004 1323 3022 1357
rect 2952 1285 3022 1323
rect 2952 1251 2970 1285
rect 3004 1251 3022 1285
rect 2952 1213 3022 1251
rect 2952 1179 2970 1213
rect 3004 1179 3022 1213
rect 2952 1160 3022 1179
rect 3270 1573 3340 1592
rect 3270 1539 3288 1573
rect 3322 1539 3340 1573
rect 3270 1501 3340 1539
rect 3270 1467 3288 1501
rect 3322 1467 3340 1501
rect 3270 1429 3340 1467
rect 3270 1395 3288 1429
rect 3322 1395 3340 1429
rect 3270 1357 3340 1395
rect 3270 1323 3288 1357
rect 3322 1323 3340 1357
rect 3270 1285 3340 1323
rect 3270 1251 3288 1285
rect 3322 1251 3340 1285
rect 3270 1213 3340 1251
rect 3270 1179 3288 1213
rect 3322 1179 3340 1213
rect 3270 1160 3340 1179
rect 113 526 183 545
rect 113 492 131 526
rect 165 492 183 526
rect 113 454 183 492
rect 113 420 131 454
rect 165 420 183 454
rect 113 382 183 420
rect 113 348 131 382
rect 165 348 183 382
rect 113 310 183 348
rect 113 276 131 310
rect 165 276 183 310
rect 113 238 183 276
rect 113 204 131 238
rect 165 204 183 238
rect 113 166 183 204
rect 113 132 131 166
rect 165 132 183 166
rect 113 113 183 132
rect 431 526 501 545
rect 431 492 449 526
rect 483 492 501 526
rect 431 454 501 492
rect 431 420 449 454
rect 483 420 501 454
rect 431 382 501 420
rect 431 348 449 382
rect 483 348 501 382
rect 431 310 501 348
rect 431 276 449 310
rect 483 276 501 310
rect 431 238 501 276
rect 431 204 449 238
rect 483 204 501 238
rect 431 166 501 204
rect 431 132 449 166
rect 483 132 501 166
rect 431 113 501 132
rect 749 526 819 545
rect 749 492 767 526
rect 801 492 819 526
rect 749 454 819 492
rect 749 420 767 454
rect 801 420 819 454
rect 749 382 819 420
rect 749 348 767 382
rect 801 348 819 382
rect 749 310 819 348
rect 749 276 767 310
rect 801 276 819 310
rect 749 238 819 276
rect 749 204 767 238
rect 801 204 819 238
rect 749 166 819 204
rect 749 132 767 166
rect 801 132 819 166
rect 749 113 819 132
rect 1067 526 1137 545
rect 1067 492 1085 526
rect 1119 492 1137 526
rect 1067 454 1137 492
rect 1067 420 1085 454
rect 1119 420 1137 454
rect 1067 382 1137 420
rect 1067 348 1085 382
rect 1119 348 1137 382
rect 1067 310 1137 348
rect 1067 276 1085 310
rect 1119 276 1137 310
rect 1067 238 1137 276
rect 1067 204 1085 238
rect 1119 204 1137 238
rect 1067 166 1137 204
rect 1067 132 1085 166
rect 1119 132 1137 166
rect 1067 113 1137 132
rect 2316 521 2386 540
rect 2316 487 2334 521
rect 2368 487 2386 521
rect 2316 449 2386 487
rect 2316 415 2334 449
rect 2368 415 2386 449
rect 2316 377 2386 415
rect 2316 343 2334 377
rect 2368 343 2386 377
rect 2316 305 2386 343
rect 2316 271 2334 305
rect 2368 271 2386 305
rect 2316 233 2386 271
rect 2316 199 2334 233
rect 2368 199 2386 233
rect 2316 161 2386 199
rect 2316 127 2334 161
rect 2368 127 2386 161
rect 2316 108 2386 127
rect 2634 521 2704 540
rect 2634 487 2652 521
rect 2686 487 2704 521
rect 2634 449 2704 487
rect 2634 415 2652 449
rect 2686 415 2704 449
rect 2634 377 2704 415
rect 2634 343 2652 377
rect 2686 343 2704 377
rect 2634 305 2704 343
rect 2634 271 2652 305
rect 2686 271 2704 305
rect 2634 233 2704 271
rect 2634 199 2652 233
rect 2686 199 2704 233
rect 2634 161 2704 199
rect 2634 127 2652 161
rect 2686 127 2704 161
rect 2634 108 2704 127
rect 2952 521 3022 540
rect 2952 487 2970 521
rect 3004 487 3022 521
rect 2952 449 3022 487
rect 2952 415 2970 449
rect 3004 415 3022 449
rect 2952 377 3022 415
rect 2952 343 2970 377
rect 3004 343 3022 377
rect 2952 305 3022 343
rect 2952 271 2970 305
rect 3004 271 3022 305
rect 2952 233 3022 271
rect 2952 199 2970 233
rect 3004 199 3022 233
rect 2952 161 3022 199
rect 2952 127 2970 161
rect 3004 127 3022 161
rect 2952 108 3022 127
rect 3270 521 3340 540
rect 3270 487 3288 521
rect 3322 487 3340 521
rect 3270 449 3340 487
rect 3270 415 3288 449
rect 3322 415 3340 449
rect 3270 377 3340 415
rect 3270 343 3288 377
rect 3322 343 3340 377
rect 3270 305 3340 343
rect 3270 271 3288 305
rect 3322 271 3340 305
rect 3270 233 3340 271
rect 3270 199 3288 233
rect 3322 199 3340 233
rect 3270 161 3340 199
rect 3270 127 3288 161
rect 3322 127 3340 161
rect 3270 108 3340 127
rect 240 19 312 20
rect 240 -15 259 19
rect 293 -15 312 19
rect 240 -16 312 -15
rect 608 19 680 20
rect 608 -15 627 19
rect 661 -15 680 19
rect 608 -16 680 -15
rect 920 19 992 20
rect 920 -15 939 19
rect 973 -15 992 19
rect 920 -16 992 -15
rect 2282 -22 2307 12
rect 2341 -22 2379 12
rect 2413 -22 2451 12
rect 2485 -22 2523 12
rect 2557 -22 2595 12
rect 2629 -22 2667 12
rect 2701 -22 2739 12
rect 2773 -22 2811 12
rect 2845 -22 2883 12
rect 2917 -22 2955 12
rect 2989 -22 3027 12
rect 3061 -22 3099 12
rect 3133 -22 3171 12
rect 3205 -22 3243 12
rect 3277 -22 3315 12
rect 3349 -22 3374 12
rect 1644 -360 1680 -346
rect 1644 -394 1645 -360
rect 1679 -394 1680 -360
rect 1644 -408 1680 -394
rect 1826 -366 1862 -352
rect 1826 -400 1827 -366
rect 1861 -400 1862 -366
rect 1826 -414 1862 -400
rect 2246 -356 2282 -342
rect 2246 -390 2247 -356
rect 2281 -390 2282 -356
rect 2246 -404 2282 -390
rect 490 -908 493 -874
rect 527 -908 565 -874
rect 599 -908 637 -874
rect 671 -908 709 -874
rect 743 -908 781 -874
rect 815 -908 853 -874
rect 887 -908 925 -874
rect 959 -908 997 -874
rect 1031 -908 1069 -874
rect 1103 -908 1141 -874
rect 1175 -908 1213 -874
rect 1247 -908 1285 -874
rect 1319 -908 1357 -874
rect 1391 -908 1429 -874
rect 1463 -908 1466 -874
rect 2236 -894 2243 -860
rect 2277 -894 2284 -860
rect 406 -959 440 -936
rect 406 -1031 440 -993
rect 406 -1103 440 -1065
rect 406 -1175 440 -1137
rect 406 -1247 440 -1209
rect 406 -1304 440 -1281
rect 1516 -959 1550 -936
rect 1516 -1031 1550 -993
rect 1516 -1103 1550 -1065
rect 1516 -1175 1550 -1137
rect 1516 -1247 1550 -1209
rect 1516 -1304 1550 -1281
rect 1968 -947 2002 -924
rect 1968 -1019 2002 -981
rect 1968 -1091 2002 -1053
rect 1968 -1163 2002 -1125
rect 1968 -1235 2002 -1197
rect 1968 -1292 2002 -1269
rect 934 -1366 949 -1332
rect 983 -1366 1021 -1332
rect 1055 -1366 1070 -1332
rect 2494 -1354 2507 -1320
rect 2541 -1354 2579 -1320
rect 2613 -1354 2626 -1320
rect 400 -1480 421 -1446
rect 455 -1480 493 -1446
rect 527 -1480 565 -1446
rect 599 -1480 637 -1446
rect 671 -1480 709 -1446
rect 743 -1480 781 -1446
rect 815 -1480 853 -1446
rect 887 -1480 925 -1446
rect 959 -1480 997 -1446
rect 1031 -1480 1069 -1446
rect 1103 -1480 1141 -1446
rect 1175 -1480 1213 -1446
rect 1247 -1480 1285 -1446
rect 1319 -1480 1357 -1446
rect 1391 -1480 1429 -1446
rect 1463 -1480 1501 -1446
rect 1535 -1480 1556 -1446
rect 1962 -1468 1983 -1434
rect 2017 -1468 2055 -1434
rect 2089 -1468 2127 -1434
rect 2161 -1468 2199 -1434
rect 2233 -1468 2271 -1434
rect 2305 -1468 2343 -1434
rect 2377 -1468 2415 -1434
rect 2449 -1468 2487 -1434
rect 2521 -1468 2559 -1434
rect 2593 -1468 2631 -1434
rect 2665 -1468 2703 -1434
rect 2737 -1468 2775 -1434
rect 2809 -1468 2847 -1434
rect 2881 -1468 2919 -1434
rect 2953 -1468 2991 -1434
rect 3025 -1468 3063 -1434
rect 3097 -1468 3118 -1434
<< viali >>
rect 261 1988 295 2022
rect 571 1982 605 2016
rect 887 1976 921 2010
rect 1363 1982 1397 2016
rect 2037 1986 2071 2020
rect 2477 1988 2511 2022
rect 2771 1988 2805 2022
rect 3073 1988 3107 2022
rect 131 1544 165 1578
rect 131 1472 165 1506
rect 131 1400 165 1434
rect 131 1328 165 1362
rect 131 1256 165 1290
rect 131 1184 165 1218
rect 449 1544 483 1578
rect 449 1472 483 1506
rect 449 1400 483 1434
rect 449 1328 483 1362
rect 449 1256 483 1290
rect 449 1184 483 1218
rect 767 1544 801 1578
rect 767 1472 801 1506
rect 767 1400 801 1434
rect 767 1328 801 1362
rect 767 1256 801 1290
rect 767 1184 801 1218
rect 1085 1544 1119 1578
rect 1085 1472 1119 1506
rect 1085 1400 1119 1434
rect 1085 1328 1119 1362
rect 1085 1256 1119 1290
rect 1085 1184 1119 1218
rect 2334 1539 2368 1573
rect 2334 1467 2368 1501
rect 2334 1395 2368 1429
rect 2334 1323 2368 1357
rect 2334 1251 2368 1285
rect 2334 1179 2368 1213
rect 2652 1539 2686 1573
rect 2652 1467 2686 1501
rect 2652 1395 2686 1429
rect 2652 1323 2686 1357
rect 2652 1251 2686 1285
rect 2652 1179 2686 1213
rect 2970 1539 3004 1573
rect 2970 1467 3004 1501
rect 2970 1395 3004 1429
rect 2970 1323 3004 1357
rect 2970 1251 3004 1285
rect 2970 1179 3004 1213
rect 3288 1539 3322 1573
rect 3288 1467 3322 1501
rect 3288 1395 3322 1429
rect 3288 1323 3322 1357
rect 3288 1251 3322 1285
rect 3288 1179 3322 1213
rect 131 492 165 526
rect 131 420 165 454
rect 131 348 165 382
rect 131 276 165 310
rect 131 204 165 238
rect 131 132 165 166
rect 449 492 483 526
rect 449 420 483 454
rect 449 348 483 382
rect 449 276 483 310
rect 449 204 483 238
rect 449 132 483 166
rect 767 492 801 526
rect 767 420 801 454
rect 767 348 801 382
rect 767 276 801 310
rect 767 204 801 238
rect 767 132 801 166
rect 1085 492 1119 526
rect 1085 420 1119 454
rect 1085 348 1119 382
rect 1085 276 1119 310
rect 1085 204 1119 238
rect 1085 132 1119 166
rect 2334 487 2368 521
rect 2334 415 2368 449
rect 2334 343 2368 377
rect 2334 271 2368 305
rect 2334 199 2368 233
rect 2334 127 2368 161
rect 2652 487 2686 521
rect 2652 415 2686 449
rect 2652 343 2686 377
rect 2652 271 2686 305
rect 2652 199 2686 233
rect 2652 127 2686 161
rect 2970 487 3004 521
rect 2970 415 3004 449
rect 2970 343 3004 377
rect 2970 271 3004 305
rect 2970 199 3004 233
rect 2970 127 3004 161
rect 3288 487 3322 521
rect 3288 415 3322 449
rect 3288 343 3322 377
rect 3288 271 3322 305
rect 3288 199 3322 233
rect 3288 127 3322 161
rect 259 -15 293 19
rect 627 -15 661 19
rect 939 -15 973 19
rect 2307 -22 2341 12
rect 2379 -22 2413 12
rect 2451 -22 2485 12
rect 2523 -22 2557 12
rect 2595 -22 2629 12
rect 2667 -22 2701 12
rect 2739 -22 2773 12
rect 2811 -22 2845 12
rect 2883 -22 2917 12
rect 2955 -22 2989 12
rect 3027 -22 3061 12
rect 3099 -22 3133 12
rect 3171 -22 3205 12
rect 3243 -22 3277 12
rect 3315 -22 3349 12
rect 1645 -394 1679 -360
rect 1827 -400 1861 -366
rect 2247 -390 2281 -356
rect 1386 -500 1420 -466
rect 1988 -500 2022 -466
rect 493 -908 527 -874
rect 565 -908 599 -874
rect 637 -908 671 -874
rect 709 -908 743 -874
rect 781 -908 815 -874
rect 853 -908 887 -874
rect 925 -908 959 -874
rect 997 -908 1031 -874
rect 1069 -908 1103 -874
rect 1141 -908 1175 -874
rect 1213 -908 1247 -874
rect 1285 -908 1319 -874
rect 1357 -908 1391 -874
rect 1429 -908 1463 -874
rect 2243 -894 2277 -860
rect 406 -993 440 -959
rect 406 -1065 440 -1031
rect 406 -1137 440 -1103
rect 406 -1209 440 -1175
rect 406 -1281 440 -1247
rect 1516 -993 1550 -959
rect 1516 -1065 1550 -1031
rect 1516 -1137 1550 -1103
rect 1516 -1209 1550 -1175
rect 1516 -1281 1550 -1247
rect 1968 -981 2002 -947
rect 1968 -1053 2002 -1019
rect 1968 -1125 2002 -1091
rect 1968 -1197 2002 -1163
rect 1968 -1269 2002 -1235
rect 949 -1366 983 -1332
rect 1021 -1366 1055 -1332
rect 2507 -1354 2541 -1320
rect 2579 -1354 2613 -1320
rect 421 -1480 455 -1446
rect 493 -1480 527 -1446
rect 565 -1480 599 -1446
rect 637 -1480 671 -1446
rect 709 -1480 743 -1446
rect 781 -1480 815 -1446
rect 853 -1480 887 -1446
rect 925 -1480 959 -1446
rect 997 -1480 1031 -1446
rect 1069 -1480 1103 -1446
rect 1141 -1480 1175 -1446
rect 1213 -1480 1247 -1446
rect 1285 -1480 1319 -1446
rect 1357 -1480 1391 -1446
rect 1429 -1480 1463 -1446
rect 1501 -1480 1535 -1446
rect 1983 -1468 2017 -1434
rect 2055 -1468 2089 -1434
rect 2127 -1468 2161 -1434
rect 2199 -1468 2233 -1434
rect 2271 -1468 2305 -1434
rect 2343 -1468 2377 -1434
rect 2415 -1468 2449 -1434
rect 2487 -1468 2521 -1434
rect 2559 -1468 2593 -1434
rect 2631 -1468 2665 -1434
rect 2703 -1468 2737 -1434
rect 2775 -1468 2809 -1434
rect 2847 -1468 2881 -1434
rect 2919 -1468 2953 -1434
rect 2991 -1468 3025 -1434
rect 3063 -1468 3097 -1434
<< metal1 >>
rect 94 2106 3230 2114
rect 94 2022 3360 2106
rect 94 1988 261 2022
rect 295 2020 2477 2022
rect 295 2016 2037 2020
rect 295 1988 571 2016
rect 94 1982 571 1988
rect 605 2010 1363 2016
rect 605 1982 887 2010
rect 94 1976 887 1982
rect 921 1982 1363 2010
rect 1397 1986 2037 2016
rect 2071 1988 2477 2020
rect 2511 1988 2771 2022
rect 2805 1988 3073 2022
rect 3107 1988 3360 2022
rect 2071 1986 3360 1988
rect 1397 1982 3360 1986
rect 921 1976 3360 1982
rect 94 1888 3360 1976
rect 94 1578 206 1888
rect 94 1544 131 1578
rect 165 1544 206 1578
rect 94 1506 206 1544
rect 94 1472 131 1506
rect 165 1472 206 1506
rect 94 1434 206 1472
rect 94 1400 131 1434
rect 165 1400 206 1434
rect 94 1362 206 1400
rect 94 1328 131 1362
rect 165 1328 206 1362
rect 94 1290 206 1328
rect 94 1256 131 1290
rect 165 1256 206 1290
rect 94 1218 206 1256
rect 94 1184 131 1218
rect 165 1184 206 1218
rect 94 1142 206 1184
rect 404 1578 842 1626
rect 404 1544 449 1578
rect 483 1544 767 1578
rect 801 1544 842 1578
rect 404 1506 842 1544
rect 404 1472 449 1506
rect 483 1472 767 1506
rect 801 1472 842 1506
rect 404 1434 842 1472
rect 404 1400 449 1434
rect 483 1400 767 1434
rect 801 1400 842 1434
rect 404 1362 842 1400
rect 404 1328 449 1362
rect 483 1328 767 1362
rect 801 1328 842 1362
rect 404 1290 842 1328
rect 404 1256 449 1290
rect 483 1256 767 1290
rect 801 1256 842 1290
rect 404 1218 842 1256
rect 404 1184 449 1218
rect 483 1184 767 1218
rect 801 1184 842 1218
rect 404 1136 842 1184
rect 1044 1578 1476 1622
rect 1044 1544 1085 1578
rect 1119 1544 1476 1578
rect 1044 1506 1476 1544
rect 1044 1472 1085 1506
rect 1119 1472 1476 1506
rect 1044 1434 1476 1472
rect 1044 1400 1085 1434
rect 1119 1400 1476 1434
rect 1044 1362 1476 1400
rect 1044 1328 1085 1362
rect 1119 1328 1476 1362
rect 1044 1290 1476 1328
rect 1044 1256 1085 1290
rect 1119 1256 1476 1290
rect 1044 1218 1476 1256
rect 1044 1184 1085 1218
rect 1119 1184 1476 1218
rect 1044 1148 1476 1184
rect 88 526 524 564
rect 88 492 131 526
rect 165 492 449 526
rect 483 492 524 526
rect 88 454 524 492
rect 88 420 131 454
rect 165 420 449 454
rect 483 420 524 454
rect 88 382 524 420
rect 88 348 131 382
rect 165 348 449 382
rect 483 348 524 382
rect 88 310 524 348
rect 88 276 131 310
rect 165 276 449 310
rect 483 276 524 310
rect 88 238 524 276
rect 88 204 131 238
rect 165 204 449 238
rect 483 204 524 238
rect 88 166 524 204
rect 88 132 131 166
rect 165 132 449 166
rect 483 132 524 166
rect 88 90 524 132
rect 732 526 1154 560
rect 732 492 767 526
rect 801 492 1085 526
rect 1119 492 1154 526
rect 732 454 1154 492
rect 732 420 767 454
rect 801 420 1085 454
rect 1119 420 1154 454
rect 732 382 1154 420
rect 732 348 767 382
rect 801 348 1085 382
rect 1119 348 1154 382
rect 732 310 1154 348
rect 732 276 767 310
rect 801 276 1085 310
rect 1119 276 1154 310
rect 732 238 1154 276
rect 732 204 767 238
rect 801 204 1085 238
rect 1119 204 1154 238
rect 732 166 1154 204
rect 732 132 767 166
rect 801 132 1085 166
rect 1119 132 1154 166
rect 732 102 1154 132
rect 964 28 1206 30
rect 68 19 1206 28
rect 68 -15 259 19
rect 293 -15 627 19
rect 661 -15 939 19
rect 973 -15 1206 19
rect 68 -28 1206 -15
rect 224 -1402 350 -28
rect 1428 -198 1476 1148
rect 2004 1573 2414 1610
rect 2004 1539 2334 1573
rect 2368 1539 2414 1573
rect 2004 1501 2414 1539
rect 2004 1467 2334 1501
rect 2368 1467 2414 1501
rect 2004 1429 2414 1467
rect 2004 1395 2334 1429
rect 2368 1395 2414 1429
rect 2004 1357 2414 1395
rect 2004 1323 2334 1357
rect 2368 1323 2414 1357
rect 2004 1285 2414 1323
rect 2004 1251 2334 1285
rect 2368 1251 2414 1285
rect 2004 1213 2414 1251
rect 2004 1179 2334 1213
rect 2368 1179 2414 1213
rect 2004 1142 2414 1179
rect 2616 1573 3040 1616
rect 2616 1539 2652 1573
rect 2686 1539 2970 1573
rect 3004 1539 3040 1573
rect 2616 1501 3040 1539
rect 2616 1467 2652 1501
rect 2686 1467 2970 1501
rect 3004 1467 3040 1501
rect 2616 1429 3040 1467
rect 2616 1395 2652 1429
rect 2686 1395 2970 1429
rect 3004 1395 3040 1429
rect 2616 1357 3040 1395
rect 2616 1323 2652 1357
rect 2686 1323 2970 1357
rect 3004 1323 3040 1357
rect 2616 1285 3040 1323
rect 2616 1251 2652 1285
rect 2686 1251 2970 1285
rect 3004 1251 3040 1285
rect 2616 1213 3040 1251
rect 2616 1179 2652 1213
rect 2686 1179 2970 1213
rect 3004 1179 3040 1213
rect 2616 1142 3040 1179
rect 3254 1573 3360 1888
rect 3254 1539 3288 1573
rect 3322 1539 3360 1573
rect 3254 1501 3360 1539
rect 3254 1467 3288 1501
rect 3322 1467 3360 1501
rect 3254 1429 3360 1467
rect 3254 1395 3288 1429
rect 3322 1395 3360 1429
rect 3254 1357 3360 1395
rect 3254 1323 3288 1357
rect 3322 1323 3360 1357
rect 3254 1285 3360 1323
rect 3254 1251 3288 1285
rect 3322 1251 3360 1285
rect 3254 1213 3360 1251
rect 3254 1179 3288 1213
rect 3322 1179 3360 1213
rect 3254 1144 3360 1179
rect 1212 -430 1378 -316
rect 1428 -324 1474 -198
rect 1822 -316 1982 -314
rect 1816 -320 1982 -316
rect 1428 -335 1460 -324
rect 1524 -334 1982 -320
rect 2030 -329 2076 1142
rect 2286 521 2724 554
rect 2286 487 2334 521
rect 2368 487 2652 521
rect 2686 487 2724 521
rect 2286 449 2724 487
rect 2286 415 2334 449
rect 2368 415 2652 449
rect 2686 415 2724 449
rect 2286 377 2724 415
rect 2286 343 2334 377
rect 2368 343 2652 377
rect 2686 343 2724 377
rect 2286 305 2724 343
rect 2286 271 2334 305
rect 2368 271 2652 305
rect 2686 271 2724 305
rect 2286 233 2724 271
rect 2286 199 2334 233
rect 2368 199 2652 233
rect 2686 199 2724 233
rect 2286 161 2724 199
rect 2286 127 2334 161
rect 2368 127 2652 161
rect 2686 127 2724 161
rect 2286 86 2724 127
rect 2942 521 3362 560
rect 2942 487 2970 521
rect 3004 487 3288 521
rect 3322 487 3362 521
rect 2942 449 3362 487
rect 2942 415 2970 449
rect 3004 415 3288 449
rect 3322 415 3362 449
rect 2942 377 3362 415
rect 2942 343 2970 377
rect 3004 343 3288 377
rect 3322 343 3362 377
rect 2942 305 3362 343
rect 2942 271 2970 305
rect 3004 271 3288 305
rect 3322 271 3362 305
rect 2942 233 3362 271
rect 2942 199 2970 233
rect 3004 199 3288 233
rect 3322 199 3362 233
rect 2942 161 3362 199
rect 2942 127 2970 161
rect 3004 127 3288 161
rect 3322 127 3362 161
rect 2942 96 3362 127
rect 2270 12 3380 24
rect 2270 -22 2307 12
rect 2341 -22 2379 12
rect 2413 -22 2451 12
rect 2485 -22 2523 12
rect 2557 -22 2595 12
rect 2629 -22 2667 12
rect 2701 -22 2739 12
rect 2773 -22 2811 12
rect 2845 -22 2883 12
rect 2917 -22 2955 12
rect 2989 -22 3027 12
rect 3061 -22 3099 12
rect 3133 -22 3171 12
rect 3205 -22 3243 12
rect 3277 -22 3315 12
rect 3349 -22 3380 12
rect 2270 -42 3380 -22
rect 2158 -314 2294 -310
rect 1524 -360 1940 -334
rect 1524 -394 1645 -360
rect 1679 -366 1940 -360
rect 1679 -394 1827 -366
rect 1524 -400 1827 -394
rect 1861 -400 1940 -366
rect 1524 -420 1940 -400
rect 1974 -420 1982 -334
rect 1524 -428 1982 -420
rect 2126 -334 2294 -314
rect 2126 -420 2132 -334
rect 2166 -356 2294 -334
rect 2166 -390 2247 -356
rect 2281 -390 2294 -356
rect 2166 -420 2294 -390
rect 1212 -444 1306 -430
rect 1524 -440 1926 -428
rect 2126 -440 2294 -420
rect 1524 -442 1886 -440
rect 1524 -448 1880 -442
rect 1524 -450 1694 -448
rect 1372 -466 1440 -460
rect 1372 -500 1386 -466
rect 1420 -500 1440 -466
rect 1372 -510 1440 -500
rect 1972 -466 2034 -456
rect 1972 -500 1988 -466
rect 2022 -500 2034 -466
rect 1972 -512 2034 -500
rect 384 -874 1566 -858
rect 384 -908 493 -874
rect 527 -908 565 -874
rect 599 -908 637 -874
rect 671 -908 709 -874
rect 743 -908 781 -874
rect 815 -908 853 -874
rect 887 -908 925 -874
rect 959 -908 997 -874
rect 1031 -908 1069 -874
rect 1103 -908 1141 -874
rect 1175 -908 1213 -874
rect 1247 -908 1285 -874
rect 1319 -908 1357 -874
rect 1391 -908 1429 -874
rect 1463 -902 1566 -874
rect 2228 -860 2294 -440
rect 2228 -894 2243 -860
rect 2277 -894 2294 -860
rect 1463 -908 2012 -902
rect 2228 -906 2294 -894
rect 384 -922 2012 -908
rect 384 -959 470 -922
rect 384 -993 406 -959
rect 440 -993 470 -959
rect 384 -1031 470 -993
rect 384 -1065 406 -1031
rect 440 -1065 470 -1031
rect 384 -1103 470 -1065
rect 384 -1137 406 -1103
rect 440 -1137 470 -1103
rect 384 -1175 470 -1137
rect 384 -1209 406 -1175
rect 440 -1209 470 -1175
rect 384 -1247 470 -1209
rect 384 -1281 406 -1247
rect 440 -1281 470 -1247
rect 384 -1320 470 -1281
rect 1510 -947 2012 -922
rect 1510 -959 1968 -947
rect 1510 -993 1516 -959
rect 1550 -981 1968 -959
rect 2002 -981 2012 -947
rect 1550 -993 2012 -981
rect 1510 -1019 2012 -993
rect 1510 -1031 1968 -1019
rect 1510 -1065 1516 -1031
rect 1550 -1053 1968 -1031
rect 2002 -1053 2012 -1019
rect 1550 -1065 2012 -1053
rect 1510 -1091 2012 -1065
rect 1510 -1103 1968 -1091
rect 1510 -1137 1516 -1103
rect 1550 -1125 1968 -1103
rect 2002 -1125 2012 -1091
rect 1550 -1137 2012 -1125
rect 1510 -1163 2012 -1137
rect 1510 -1175 1968 -1163
rect 1510 -1209 1516 -1175
rect 1550 -1197 1968 -1175
rect 2002 -1197 2012 -1163
rect 1550 -1209 2012 -1197
rect 1510 -1235 2012 -1209
rect 1510 -1247 1968 -1235
rect 1510 -1281 1516 -1247
rect 1550 -1269 1968 -1247
rect 2002 -1269 2012 -1235
rect 1550 -1281 2012 -1269
rect 1510 -1326 2012 -1281
rect 2436 -1320 2714 -1312
rect 884 -1332 1132 -1326
rect 884 -1366 949 -1332
rect 983 -1366 1021 -1332
rect 1055 -1366 1132 -1332
rect 884 -1402 1132 -1366
rect 2436 -1354 2507 -1320
rect 2541 -1354 2579 -1320
rect 2613 -1354 2714 -1320
rect 222 -1404 1668 -1402
rect 2436 -1404 2714 -1354
rect 3146 -1402 3228 -42
rect 3030 -1404 3238 -1402
rect 222 -1434 3238 -1404
rect 222 -1446 1983 -1434
rect 222 -1480 421 -1446
rect 455 -1480 493 -1446
rect 527 -1480 565 -1446
rect 599 -1480 637 -1446
rect 671 -1480 709 -1446
rect 743 -1480 781 -1446
rect 815 -1480 853 -1446
rect 887 -1480 925 -1446
rect 959 -1480 997 -1446
rect 1031 -1480 1069 -1446
rect 1103 -1480 1141 -1446
rect 1175 -1480 1213 -1446
rect 1247 -1480 1285 -1446
rect 1319 -1480 1357 -1446
rect 1391 -1480 1429 -1446
rect 1463 -1480 1501 -1446
rect 1535 -1468 1983 -1446
rect 2017 -1468 2055 -1434
rect 2089 -1468 2127 -1434
rect 2161 -1468 2199 -1434
rect 2233 -1468 2271 -1434
rect 2305 -1468 2343 -1434
rect 2377 -1468 2415 -1434
rect 2449 -1468 2487 -1434
rect 2521 -1468 2559 -1434
rect 2593 -1468 2631 -1434
rect 2665 -1468 2703 -1434
rect 2737 -1468 2775 -1434
rect 2809 -1468 2847 -1434
rect 2881 -1468 2919 -1434
rect 2953 -1468 2991 -1434
rect 3025 -1468 3063 -1434
rect 3097 -1468 3238 -1434
rect 1535 -1480 3238 -1468
rect 222 -1582 3238 -1480
rect 1660 -1584 3106 -1582
use sky130_fd_pr__nfet_01v8_lvt_F9NR5A  sky130_fd_pr__nfet_01v8_lvt_F9NR5A_0
timestamp 1611881054
transform 0 1 976 -1 0 -1120
box -360 -674 360 674
use sky130_fd_pr__res_xhigh_po_0p35_RRCNTY  sky130_fd_pr__res_xhigh_po_0p35_RRCNTY_0
timestamp 1611881054
transform 1 0 625 0 1 855
box -642 -872 642 872
use sky130_fd_pr__nfet_01v8_N9UHYA  sky130_fd_pr__nfet_01v8_N9UHYA_0
timestamp 1611881054
transform 1 0 1451 0 1 -374
box -227 -228 227 228
use sky130_fd_pr__nfet_01v8_N9UHYA  sky130_fd_pr__nfet_01v8_N9UHYA_1
timestamp 1611881054
transform 1 0 2053 0 1 -374
box -227 -228 227 228
use sky130_fd_pr__nfet_01v8_lvt_F9NR5A  sky130_fd_pr__nfet_01v8_lvt_F9NR5A_1
timestamp 1611881054
transform 0 1 2542 -1 0 -1106
box -360 -674 360 674
use sky130_fd_pr__res_xhigh_po_0p35_RRCNTY  sky130_fd_pr__res_xhigh_po_0p35_RRCNTY_1
timestamp 1611881054
transform 1 0 2828 0 1 850
box -642 -872 642 872
<< labels >>
rlabel metal1 s 2244 -690 2270 -666 4 Itail_a
rlabel metal1 s 1676 1966 1770 2038 4 Vdd
port 1 nsew
rlabel metal1 s 2018 1326 2108 1452 4 ON2a
port 2 nsew
rlabel metal1 s 1370 1334 1460 1460 4 ON1a
port 3 nsew
rlabel poly s 1390 -276 1408 -252 4 VP
port 4 nsew
rlabel poly s 1996 -272 2014 -248 4 VN
port 5 nsew
rlabel metal1 s 1720 -1526 1794 -1482 4 Gnd
port 6 nsew
rlabel metal1 s 1720 -1144 1792 -1080 4 vbiasn
port 7 nsew
<< end >>
