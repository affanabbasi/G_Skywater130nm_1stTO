magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< locali >>
rect 3174 662 3226 664
rect -102 618 3226 662
rect -102 614 3132 618
rect -100 366 -52 614
rect 458 527 466 561
rect -100 332 28 366
rect 202 253 242 254
rect 202 219 205 253
rect 239 219 242 253
rect 202 218 242 219
rect 440 216 612 260
rect 740 254 754 260
rect 1092 252 1308 260
rect 614 216 616 220
rect 442 215 616 216
rect 650 216 654 220
rect 740 218 754 220
rect 650 215 666 216
rect 1102 218 1308 252
rect 1446 252 1662 260
rect 1448 218 1662 252
rect 1092 216 1308 218
rect 1446 216 1662 218
rect 1796 216 2012 260
rect 2148 254 2364 260
rect 2500 254 2716 260
rect 3174 258 3226 618
rect 2150 220 2364 254
rect 2148 216 2364 220
rect 2504 220 2716 254
rect 2500 216 2716 220
rect 2728 249 2762 250
rect 2852 220 3226 258
rect 2852 216 3180 220
rect 442 200 566 215
rect 458 -17 466 17
<< viali >>
rect 32 340 66 374
rect 205 219 239 253
rect 720 220 754 254
rect 968 215 1002 249
rect 1068 218 1102 252
rect 1314 222 1348 256
rect 1414 218 1448 252
rect 1664 220 1698 254
rect 1762 220 1796 254
rect 2016 220 2050 254
rect 2116 220 2150 254
rect 2376 218 2410 252
rect 2470 220 2504 254
rect 2728 215 2762 249
rect 2818 216 2852 250
<< metal1 >>
rect 3172 708 4272 714
rect -118 625 4272 708
rect -118 622 4043 625
rect -118 390 -36 622
rect 4 582 1630 594
rect 1634 582 3118 592
rect 4 578 3118 582
rect 4 526 26 578
rect 78 526 90 578
rect 142 526 154 578
rect 206 526 218 578
rect 270 526 282 578
rect 334 526 346 578
rect 398 526 410 578
rect 462 526 474 578
rect 526 526 538 578
rect 590 526 602 578
rect 654 526 666 578
rect 718 526 730 578
rect 782 526 794 578
rect 846 526 858 578
rect 910 526 922 578
rect 974 526 986 578
rect 1038 526 1050 578
rect 1102 526 1114 578
rect 1166 526 1178 578
rect 1230 526 1242 578
rect 1294 526 1306 578
rect 1358 526 1370 578
rect 1422 526 1434 578
rect 1486 526 1498 578
rect 1550 526 1562 578
rect 1614 526 1626 578
rect 1678 526 1690 578
rect 1742 526 1754 578
rect 1806 526 1818 578
rect 1870 526 1882 578
rect 1934 526 1946 578
rect 1998 526 2010 578
rect 2062 526 2074 578
rect 2126 526 2138 578
rect 2190 526 2202 578
rect 2254 526 2266 578
rect 2318 526 2330 578
rect 2382 526 2394 578
rect 2446 526 2458 578
rect 2510 526 2522 578
rect 2574 526 2586 578
rect 2638 526 2650 578
rect 2702 526 2714 578
rect 2766 526 2778 578
rect 2830 526 2842 578
rect 2894 526 2906 578
rect 2958 526 2970 578
rect 3022 526 3034 578
rect 3086 526 3118 578
rect 4 522 3118 526
rect 4 498 1630 522
rect 460 496 464 498
rect 1634 496 3118 522
rect -118 374 86 390
rect -118 340 32 374
rect 66 340 86 374
rect -118 324 86 340
rect -658 273 -250 304
rect -658 221 -595 273
rect -543 221 -531 273
rect -479 221 -467 273
rect -415 221 -403 273
rect -351 221 -339 273
rect -287 260 -250 273
rect -287 253 256 260
rect -287 221 205 253
rect -658 219 205 221
rect 239 219 256 253
rect -658 212 256 219
rect 698 254 1020 266
rect 698 220 720 254
rect 754 249 1020 254
rect 754 220 968 249
rect 698 215 968 220
rect 1002 215 1020 249
rect -658 184 -250 212
rect 698 198 1020 215
rect 1052 256 1372 264
rect 1052 252 1314 256
rect 1052 218 1068 252
rect 1102 222 1314 252
rect 1348 222 1372 256
rect 1102 218 1372 222
rect 1052 196 1372 218
rect 1400 254 1720 266
rect 1400 252 1664 254
rect 1400 218 1414 252
rect 1448 220 1664 252
rect 1698 220 1720 254
rect 1448 218 1720 220
rect 1400 198 1720 218
rect 1756 254 2076 266
rect 1756 220 1762 254
rect 1796 220 2016 254
rect 2050 220 2076 254
rect 1756 198 2076 220
rect 2106 254 2426 268
rect 2106 220 2116 254
rect 2150 252 2426 254
rect 2150 220 2376 252
rect 2106 218 2376 220
rect 2410 218 2426 252
rect 2106 200 2426 218
rect 2462 254 2782 268
rect 3172 264 4043 622
rect 2462 220 2470 254
rect 2504 249 2782 254
rect 2504 220 2728 249
rect 2462 215 2728 220
rect 2762 215 2782 249
rect 2462 200 2782 215
rect 2812 253 4043 264
rect 4159 253 4272 625
rect 2812 250 4272 253
rect 2812 216 2818 250
rect 2852 216 4272 250
rect 2812 188 4272 216
rect 0 -594 3118 48
rect 0 -646 59 -594
rect 111 -646 123 -594
rect 175 -646 187 -594
rect 239 -646 251 -594
rect 303 -646 315 -594
rect 367 -646 379 -594
rect 431 -646 443 -594
rect 495 -646 507 -594
rect 559 -646 571 -594
rect 623 -646 635 -594
rect 687 -646 699 -594
rect 751 -646 763 -594
rect 815 -646 827 -594
rect 879 -646 891 -594
rect 943 -646 955 -594
rect 1007 -646 1019 -594
rect 1071 -646 1083 -594
rect 1135 -646 1147 -594
rect 1199 -646 1211 -594
rect 1263 -646 1275 -594
rect 1327 -646 1339 -594
rect 1391 -646 1403 -594
rect 1455 -646 1467 -594
rect 1519 -646 1531 -594
rect 1583 -646 1595 -594
rect 1647 -646 1659 -594
rect 1711 -646 1723 -594
rect 1775 -646 1787 -594
rect 1839 -646 1851 -594
rect 1903 -646 1915 -594
rect 1967 -646 1979 -594
rect 2031 -646 2043 -594
rect 2095 -646 2107 -594
rect 2159 -646 2171 -594
rect 2223 -646 2235 -594
rect 2287 -646 2299 -594
rect 2351 -646 2363 -594
rect 2415 -646 2427 -594
rect 2479 -646 2491 -594
rect 2543 -646 2555 -594
rect 2607 -646 2619 -594
rect 2671 -646 2683 -594
rect 2735 -646 2747 -594
rect 2799 -646 2811 -594
rect 2863 -646 2875 -594
rect 2927 -646 2939 -594
rect 2991 -646 3003 -594
rect 3055 -646 3118 -594
rect 0 -686 3118 -646
<< via1 >>
rect 26 526 78 578
rect 90 526 142 578
rect 154 526 206 578
rect 218 526 270 578
rect 282 526 334 578
rect 346 526 398 578
rect 410 526 462 578
rect 474 526 526 578
rect 538 526 590 578
rect 602 526 654 578
rect 666 526 718 578
rect 730 526 782 578
rect 794 526 846 578
rect 858 526 910 578
rect 922 526 974 578
rect 986 526 1038 578
rect 1050 526 1102 578
rect 1114 526 1166 578
rect 1178 526 1230 578
rect 1242 526 1294 578
rect 1306 526 1358 578
rect 1370 526 1422 578
rect 1434 526 1486 578
rect 1498 526 1550 578
rect 1562 526 1614 578
rect 1626 526 1678 578
rect 1690 526 1742 578
rect 1754 526 1806 578
rect 1818 526 1870 578
rect 1882 526 1934 578
rect 1946 526 1998 578
rect 2010 526 2062 578
rect 2074 526 2126 578
rect 2138 526 2190 578
rect 2202 526 2254 578
rect 2266 526 2318 578
rect 2330 526 2382 578
rect 2394 526 2446 578
rect 2458 526 2510 578
rect 2522 526 2574 578
rect 2586 526 2638 578
rect 2650 526 2702 578
rect 2714 526 2766 578
rect 2778 526 2830 578
rect 2842 526 2894 578
rect 2906 526 2958 578
rect 2970 526 3022 578
rect 3034 526 3086 578
rect -595 221 -543 273
rect -531 221 -479 273
rect -467 221 -415 273
rect -403 221 -351 273
rect -339 221 -287 273
rect 4043 253 4159 625
rect 59 -646 111 -594
rect 123 -646 175 -594
rect 187 -646 239 -594
rect 251 -646 303 -594
rect 315 -646 367 -594
rect 379 -646 431 -594
rect 443 -646 495 -594
rect 507 -646 559 -594
rect 571 -646 623 -594
rect 635 -646 687 -594
rect 699 -646 751 -594
rect 763 -646 815 -594
rect 827 -646 879 -594
rect 891 -646 943 -594
rect 955 -646 1007 -594
rect 1019 -646 1071 -594
rect 1083 -646 1135 -594
rect 1147 -646 1199 -594
rect 1211 -646 1263 -594
rect 1275 -646 1327 -594
rect 1339 -646 1391 -594
rect 1403 -646 1455 -594
rect 1467 -646 1519 -594
rect 1531 -646 1583 -594
rect 1595 -646 1647 -594
rect 1659 -646 1711 -594
rect 1723 -646 1775 -594
rect 1787 -646 1839 -594
rect 1851 -646 1903 -594
rect 1915 -646 1967 -594
rect 1979 -646 2031 -594
rect 2043 -646 2095 -594
rect 2107 -646 2159 -594
rect 2171 -646 2223 -594
rect 2235 -646 2287 -594
rect 2299 -646 2351 -594
rect 2363 -646 2415 -594
rect 2427 -646 2479 -594
rect 2491 -646 2543 -594
rect 2555 -646 2607 -594
rect 2619 -646 2671 -594
rect 2683 -646 2735 -594
rect 2747 -646 2799 -594
rect 2811 -646 2863 -594
rect 2875 -646 2927 -594
rect 2939 -646 2991 -594
rect 3003 -646 3055 -594
<< metal2 >>
rect -10 1422 3140 1462
rect -10 1339 3184 1422
rect -10 1283 163 1339
rect 219 1283 243 1339
rect 299 1283 323 1339
rect 379 1283 403 1339
rect 459 1283 483 1339
rect 539 1283 563 1339
rect 619 1283 643 1339
rect 699 1283 723 1339
rect 779 1283 803 1339
rect 859 1283 883 1339
rect 939 1283 963 1339
rect 1019 1283 1043 1339
rect 1099 1283 1123 1339
rect 1179 1283 1203 1339
rect 1259 1283 1283 1339
rect 1339 1283 1363 1339
rect 1419 1283 1443 1339
rect 1499 1283 1523 1339
rect 1579 1283 1603 1339
rect 1659 1283 1683 1339
rect 1739 1283 1763 1339
rect 1819 1283 1843 1339
rect 1899 1283 1923 1339
rect 1979 1283 2003 1339
rect 2059 1283 2083 1339
rect 2139 1283 2163 1339
rect 2219 1283 2243 1339
rect 2299 1283 2323 1339
rect 2379 1283 2403 1339
rect 2459 1283 2483 1339
rect 2539 1283 2563 1339
rect 2619 1283 2643 1339
rect 2699 1283 2723 1339
rect 2779 1283 2803 1339
rect 2859 1283 2883 1339
rect 2939 1283 2963 1339
rect 3019 1283 3043 1339
rect 3099 1283 3123 1339
rect 3179 1283 3184 1339
rect -10 1244 3184 1283
rect -10 578 3140 1244
rect -10 526 26 578
rect 78 526 90 578
rect 142 526 154 578
rect 206 526 218 578
rect 270 526 282 578
rect 334 526 346 578
rect 398 526 410 578
rect 462 526 474 578
rect 526 526 538 578
rect 590 526 602 578
rect 654 526 666 578
rect 718 526 730 578
rect 782 526 794 578
rect 846 526 858 578
rect 910 526 922 578
rect 974 526 986 578
rect 1038 526 1050 578
rect 1102 526 1114 578
rect 1166 526 1178 578
rect 1230 526 1242 578
rect 1294 526 1306 578
rect 1358 526 1370 578
rect 1422 526 1434 578
rect 1486 526 1498 578
rect 1550 526 1562 578
rect 1614 526 1626 578
rect 1678 526 1690 578
rect 1742 526 1754 578
rect 1806 526 1818 578
rect 1870 526 1882 578
rect 1934 526 1946 578
rect 1998 526 2010 578
rect 2062 526 2074 578
rect 2126 526 2138 578
rect 2190 526 2202 578
rect 2254 526 2266 578
rect 2318 526 2330 578
rect 2382 526 2394 578
rect 2446 526 2458 578
rect 2510 526 2522 578
rect 2574 526 2586 578
rect 2638 526 2650 578
rect 2702 526 2714 578
rect 2766 526 2778 578
rect 2830 526 2842 578
rect 2894 526 2906 578
rect 2958 526 2970 578
rect 3022 526 3034 578
rect 3086 526 3140 578
rect -10 486 3140 526
rect 3938 687 4314 798
rect -696 405 -246 482
rect -696 349 -626 405
rect -570 349 -546 405
rect -490 349 -466 405
rect -410 349 -386 405
rect -330 349 -246 405
rect -696 273 -246 349
rect -696 221 -595 273
rect -543 221 -531 273
rect -479 221 -467 273
rect -415 221 -403 273
rect -351 221 -339 273
rect -287 221 -246 273
rect -696 178 -246 221
rect 3938 231 4009 687
rect 4225 231 4314 687
rect 3938 128 4314 231
rect 0 -592 3118 -508
rect 0 -648 49 -592
rect 105 -594 129 -592
rect 185 -594 209 -592
rect 265 -594 289 -592
rect 345 -594 369 -592
rect 425 -594 449 -592
rect 505 -594 529 -592
rect 585 -594 609 -592
rect 665 -594 689 -592
rect 745 -594 769 -592
rect 825 -594 849 -592
rect 905 -594 929 -592
rect 985 -594 1009 -592
rect 1065 -594 1089 -592
rect 1145 -594 1169 -592
rect 1225 -594 1249 -592
rect 1305 -594 1329 -592
rect 1385 -594 1409 -592
rect 1465 -594 1489 -592
rect 1545 -594 1569 -592
rect 1625 -594 1649 -592
rect 1705 -594 1729 -592
rect 1785 -594 1809 -592
rect 1865 -594 1889 -592
rect 1945 -594 1969 -592
rect 2025 -594 2049 -592
rect 2105 -594 2129 -592
rect 2185 -594 2209 -592
rect 2265 -594 2289 -592
rect 2345 -594 2369 -592
rect 2425 -594 2449 -592
rect 2505 -594 2529 -592
rect 2585 -594 2609 -592
rect 2665 -594 2689 -592
rect 2745 -594 2769 -592
rect 2825 -594 2849 -592
rect 2905 -594 2929 -592
rect 2985 -594 3009 -592
rect 111 -646 123 -594
rect 185 -646 187 -594
rect 367 -646 369 -594
rect 431 -646 443 -594
rect 505 -646 507 -594
rect 687 -646 689 -594
rect 751 -646 763 -594
rect 825 -646 827 -594
rect 1007 -646 1009 -594
rect 1071 -646 1083 -594
rect 1145 -646 1147 -594
rect 1327 -646 1329 -594
rect 1391 -646 1403 -594
rect 1465 -646 1467 -594
rect 1647 -646 1649 -594
rect 1711 -646 1723 -594
rect 1785 -646 1787 -594
rect 1967 -646 1969 -594
rect 2031 -646 2043 -594
rect 2105 -646 2107 -594
rect 2287 -646 2289 -594
rect 2351 -646 2363 -594
rect 2425 -646 2427 -594
rect 2607 -646 2609 -594
rect 2671 -646 2683 -594
rect 2745 -646 2747 -594
rect 2927 -646 2929 -594
rect 2991 -646 3003 -594
rect 105 -648 129 -646
rect 185 -648 209 -646
rect 265 -648 289 -646
rect 345 -648 369 -646
rect 425 -648 449 -646
rect 505 -648 529 -646
rect 585 -648 609 -646
rect 665 -648 689 -646
rect 745 -648 769 -646
rect 825 -648 849 -646
rect 905 -648 929 -646
rect 985 -648 1009 -646
rect 1065 -648 1089 -646
rect 1145 -648 1169 -646
rect 1225 -648 1249 -646
rect 1305 -648 1329 -646
rect 1385 -648 1409 -646
rect 1465 -648 1489 -646
rect 1545 -648 1569 -646
rect 1625 -648 1649 -646
rect 1705 -648 1729 -646
rect 1785 -648 1809 -646
rect 1865 -648 1889 -646
rect 1945 -648 1969 -646
rect 2025 -648 2049 -646
rect 2105 -648 2129 -646
rect 2185 -648 2209 -646
rect 2265 -648 2289 -646
rect 2345 -648 2369 -646
rect 2425 -648 2449 -646
rect 2505 -648 2529 -646
rect 2585 -648 2609 -646
rect 2665 -648 2689 -646
rect 2745 -648 2769 -646
rect 2825 -648 2849 -646
rect 2905 -648 2929 -646
rect 2985 -648 3009 -646
rect 3065 -648 3118 -592
rect 0 -686 3118 -648
<< via2 >>
rect 163 1283 219 1339
rect 243 1283 299 1339
rect 323 1283 379 1339
rect 403 1283 459 1339
rect 483 1283 539 1339
rect 563 1283 619 1339
rect 643 1283 699 1339
rect 723 1283 779 1339
rect 803 1283 859 1339
rect 883 1283 939 1339
rect 963 1283 1019 1339
rect 1043 1283 1099 1339
rect 1123 1283 1179 1339
rect 1203 1283 1259 1339
rect 1283 1283 1339 1339
rect 1363 1283 1419 1339
rect 1443 1283 1499 1339
rect 1523 1283 1579 1339
rect 1603 1283 1659 1339
rect 1683 1283 1739 1339
rect 1763 1283 1819 1339
rect 1843 1283 1899 1339
rect 1923 1283 1979 1339
rect 2003 1283 2059 1339
rect 2083 1283 2139 1339
rect 2163 1283 2219 1339
rect 2243 1283 2299 1339
rect 2323 1283 2379 1339
rect 2403 1283 2459 1339
rect 2483 1283 2539 1339
rect 2563 1283 2619 1339
rect 2643 1283 2699 1339
rect 2723 1283 2779 1339
rect 2803 1283 2859 1339
rect 2883 1283 2939 1339
rect 2963 1283 3019 1339
rect 3043 1283 3099 1339
rect 3123 1283 3179 1339
rect -626 349 -570 405
rect -546 349 -490 405
rect -466 349 -410 405
rect -386 349 -330 405
rect 4009 625 4225 687
rect 4009 253 4043 625
rect 4043 253 4159 625
rect 4159 253 4225 625
rect 4009 231 4225 253
rect 49 -594 105 -592
rect 129 -594 185 -592
rect 209 -594 265 -592
rect 289 -594 345 -592
rect 369 -594 425 -592
rect 449 -594 505 -592
rect 529 -594 585 -592
rect 609 -594 665 -592
rect 689 -594 745 -592
rect 769 -594 825 -592
rect 849 -594 905 -592
rect 929 -594 985 -592
rect 1009 -594 1065 -592
rect 1089 -594 1145 -592
rect 1169 -594 1225 -592
rect 1249 -594 1305 -592
rect 1329 -594 1385 -592
rect 1409 -594 1465 -592
rect 1489 -594 1545 -592
rect 1569 -594 1625 -592
rect 1649 -594 1705 -592
rect 1729 -594 1785 -592
rect 1809 -594 1865 -592
rect 1889 -594 1945 -592
rect 1969 -594 2025 -592
rect 2049 -594 2105 -592
rect 2129 -594 2185 -592
rect 2209 -594 2265 -592
rect 2289 -594 2345 -592
rect 2369 -594 2425 -592
rect 2449 -594 2505 -592
rect 2529 -594 2585 -592
rect 2609 -594 2665 -592
rect 2689 -594 2745 -592
rect 2769 -594 2825 -592
rect 2849 -594 2905 -592
rect 2929 -594 2985 -592
rect 3009 -594 3065 -592
rect 49 -646 59 -594
rect 59 -646 105 -594
rect 129 -646 175 -594
rect 175 -646 185 -594
rect 209 -646 239 -594
rect 239 -646 251 -594
rect 251 -646 265 -594
rect 289 -646 303 -594
rect 303 -646 315 -594
rect 315 -646 345 -594
rect 369 -646 379 -594
rect 379 -646 425 -594
rect 449 -646 495 -594
rect 495 -646 505 -594
rect 529 -646 559 -594
rect 559 -646 571 -594
rect 571 -646 585 -594
rect 609 -646 623 -594
rect 623 -646 635 -594
rect 635 -646 665 -594
rect 689 -646 699 -594
rect 699 -646 745 -594
rect 769 -646 815 -594
rect 815 -646 825 -594
rect 849 -646 879 -594
rect 879 -646 891 -594
rect 891 -646 905 -594
rect 929 -646 943 -594
rect 943 -646 955 -594
rect 955 -646 985 -594
rect 1009 -646 1019 -594
rect 1019 -646 1065 -594
rect 1089 -646 1135 -594
rect 1135 -646 1145 -594
rect 1169 -646 1199 -594
rect 1199 -646 1211 -594
rect 1211 -646 1225 -594
rect 1249 -646 1263 -594
rect 1263 -646 1275 -594
rect 1275 -646 1305 -594
rect 1329 -646 1339 -594
rect 1339 -646 1385 -594
rect 1409 -646 1455 -594
rect 1455 -646 1465 -594
rect 1489 -646 1519 -594
rect 1519 -646 1531 -594
rect 1531 -646 1545 -594
rect 1569 -646 1583 -594
rect 1583 -646 1595 -594
rect 1595 -646 1625 -594
rect 1649 -646 1659 -594
rect 1659 -646 1705 -594
rect 1729 -646 1775 -594
rect 1775 -646 1785 -594
rect 1809 -646 1839 -594
rect 1839 -646 1851 -594
rect 1851 -646 1865 -594
rect 1889 -646 1903 -594
rect 1903 -646 1915 -594
rect 1915 -646 1945 -594
rect 1969 -646 1979 -594
rect 1979 -646 2025 -594
rect 2049 -646 2095 -594
rect 2095 -646 2105 -594
rect 2129 -646 2159 -594
rect 2159 -646 2171 -594
rect 2171 -646 2185 -594
rect 2209 -646 2223 -594
rect 2223 -646 2235 -594
rect 2235 -646 2265 -594
rect 2289 -646 2299 -594
rect 2299 -646 2345 -594
rect 2369 -646 2415 -594
rect 2415 -646 2425 -594
rect 2449 -646 2479 -594
rect 2479 -646 2491 -594
rect 2491 -646 2505 -594
rect 2529 -646 2543 -594
rect 2543 -646 2555 -594
rect 2555 -646 2585 -594
rect 2609 -646 2619 -594
rect 2619 -646 2665 -594
rect 2689 -646 2735 -594
rect 2735 -646 2745 -594
rect 2769 -646 2799 -594
rect 2799 -646 2811 -594
rect 2811 -646 2825 -594
rect 2849 -646 2863 -594
rect 2863 -646 2875 -594
rect 2875 -646 2905 -594
rect 2929 -646 2939 -594
rect 2939 -646 2985 -594
rect 3009 -646 3055 -594
rect 3055 -646 3065 -594
rect 49 -648 105 -646
rect 129 -648 185 -646
rect 209 -648 265 -646
rect 289 -648 345 -646
rect 369 -648 425 -646
rect 449 -648 505 -646
rect 529 -648 585 -646
rect 609 -648 665 -646
rect 689 -648 745 -646
rect 769 -648 825 -646
rect 849 -648 905 -646
rect 929 -648 985 -646
rect 1009 -648 1065 -646
rect 1089 -648 1145 -646
rect 1169 -648 1225 -646
rect 1249 -648 1305 -646
rect 1329 -648 1385 -646
rect 1409 -648 1465 -646
rect 1489 -648 1545 -646
rect 1569 -648 1625 -646
rect 1649 -648 1705 -646
rect 1729 -648 1785 -646
rect 1809 -648 1865 -646
rect 1889 -648 1945 -646
rect 1969 -648 2025 -646
rect 2049 -648 2105 -646
rect 2129 -648 2185 -646
rect 2209 -648 2265 -646
rect 2289 -648 2345 -646
rect 2369 -648 2425 -646
rect 2449 -648 2505 -646
rect 2529 -648 2585 -646
rect 2609 -648 2665 -646
rect 2689 -648 2745 -646
rect 2769 -648 2825 -646
rect 2849 -648 2905 -646
rect 2929 -648 2985 -646
rect 3009 -648 3065 -646
<< metal3 >>
rect 114 1343 3232 1422
rect 114 1279 159 1343
rect 223 1279 239 1343
rect 303 1279 319 1343
rect 383 1279 399 1343
rect 463 1279 479 1343
rect 543 1279 559 1343
rect 623 1279 639 1343
rect 703 1279 719 1343
rect 783 1279 799 1343
rect 863 1279 879 1343
rect 943 1279 959 1343
rect 1023 1279 1039 1343
rect 1103 1279 1119 1343
rect 1183 1279 1199 1343
rect 1263 1279 1279 1343
rect 1343 1279 1359 1343
rect 1423 1279 1439 1343
rect 1503 1279 1519 1343
rect 1583 1279 1599 1343
rect 1663 1279 1679 1343
rect 1743 1279 1759 1343
rect 1823 1279 1839 1343
rect 1903 1279 1919 1343
rect 1983 1279 1999 1343
rect 2063 1279 2079 1343
rect 2143 1279 2159 1343
rect 2223 1279 2239 1343
rect 2303 1279 2319 1343
rect 2383 1279 2399 1343
rect 2463 1279 2479 1343
rect 2543 1279 2559 1343
rect 2623 1279 2639 1343
rect 2703 1279 2719 1343
rect 2783 1279 2799 1343
rect 2863 1279 2879 1343
rect 2943 1279 2959 1343
rect 3023 1279 3039 1343
rect 3103 1279 3119 1343
rect 3183 1279 3232 1343
rect 114 1244 3232 1279
rect 3898 728 4344 854
rect -772 485 -238 564
rect -772 341 -661 485
rect -357 405 -238 485
rect -330 349 -238 405
rect -357 341 -238 349
rect -772 168 -238 341
rect 3898 184 4006 728
rect 4230 184 4344 728
rect 3898 84 4344 184
rect 0 -588 3118 -508
rect 0 -652 45 -588
rect 109 -652 125 -588
rect 189 -652 205 -588
rect 269 -652 285 -588
rect 349 -652 365 -588
rect 429 -652 445 -588
rect 509 -652 525 -588
rect 589 -652 605 -588
rect 669 -652 685 -588
rect 749 -652 765 -588
rect 829 -652 845 -588
rect 909 -652 925 -588
rect 989 -652 1005 -588
rect 1069 -652 1085 -588
rect 1149 -652 1165 -588
rect 1229 -652 1245 -588
rect 1309 -652 1325 -588
rect 1389 -652 1405 -588
rect 1469 -652 1485 -588
rect 1549 -652 1565 -588
rect 1629 -652 1645 -588
rect 1709 -652 1725 -588
rect 1789 -652 1805 -588
rect 1869 -652 1885 -588
rect 1949 -652 1965 -588
rect 2029 -652 2045 -588
rect 2109 -652 2125 -588
rect 2189 -652 2205 -588
rect 2269 -652 2285 -588
rect 2349 -652 2365 -588
rect 2429 -652 2445 -588
rect 2509 -652 2525 -588
rect 2589 -652 2605 -588
rect 2669 -652 2685 -588
rect 2749 -652 2765 -588
rect 2829 -652 2845 -588
rect 2909 -652 2925 -588
rect 2989 -652 3005 -588
rect 3069 -652 3118 -588
rect 0 -686 3118 -652
<< via3 >>
rect 159 1339 223 1343
rect 159 1283 163 1339
rect 163 1283 219 1339
rect 219 1283 223 1339
rect 159 1279 223 1283
rect 239 1339 303 1343
rect 239 1283 243 1339
rect 243 1283 299 1339
rect 299 1283 303 1339
rect 239 1279 303 1283
rect 319 1339 383 1343
rect 319 1283 323 1339
rect 323 1283 379 1339
rect 379 1283 383 1339
rect 319 1279 383 1283
rect 399 1339 463 1343
rect 399 1283 403 1339
rect 403 1283 459 1339
rect 459 1283 463 1339
rect 399 1279 463 1283
rect 479 1339 543 1343
rect 479 1283 483 1339
rect 483 1283 539 1339
rect 539 1283 543 1339
rect 479 1279 543 1283
rect 559 1339 623 1343
rect 559 1283 563 1339
rect 563 1283 619 1339
rect 619 1283 623 1339
rect 559 1279 623 1283
rect 639 1339 703 1343
rect 639 1283 643 1339
rect 643 1283 699 1339
rect 699 1283 703 1339
rect 639 1279 703 1283
rect 719 1339 783 1343
rect 719 1283 723 1339
rect 723 1283 779 1339
rect 779 1283 783 1339
rect 719 1279 783 1283
rect 799 1339 863 1343
rect 799 1283 803 1339
rect 803 1283 859 1339
rect 859 1283 863 1339
rect 799 1279 863 1283
rect 879 1339 943 1343
rect 879 1283 883 1339
rect 883 1283 939 1339
rect 939 1283 943 1339
rect 879 1279 943 1283
rect 959 1339 1023 1343
rect 959 1283 963 1339
rect 963 1283 1019 1339
rect 1019 1283 1023 1339
rect 959 1279 1023 1283
rect 1039 1339 1103 1343
rect 1039 1283 1043 1339
rect 1043 1283 1099 1339
rect 1099 1283 1103 1339
rect 1039 1279 1103 1283
rect 1119 1339 1183 1343
rect 1119 1283 1123 1339
rect 1123 1283 1179 1339
rect 1179 1283 1183 1339
rect 1119 1279 1183 1283
rect 1199 1339 1263 1343
rect 1199 1283 1203 1339
rect 1203 1283 1259 1339
rect 1259 1283 1263 1339
rect 1199 1279 1263 1283
rect 1279 1339 1343 1343
rect 1279 1283 1283 1339
rect 1283 1283 1339 1339
rect 1339 1283 1343 1339
rect 1279 1279 1343 1283
rect 1359 1339 1423 1343
rect 1359 1283 1363 1339
rect 1363 1283 1419 1339
rect 1419 1283 1423 1339
rect 1359 1279 1423 1283
rect 1439 1339 1503 1343
rect 1439 1283 1443 1339
rect 1443 1283 1499 1339
rect 1499 1283 1503 1339
rect 1439 1279 1503 1283
rect 1519 1339 1583 1343
rect 1519 1283 1523 1339
rect 1523 1283 1579 1339
rect 1579 1283 1583 1339
rect 1519 1279 1583 1283
rect 1599 1339 1663 1343
rect 1599 1283 1603 1339
rect 1603 1283 1659 1339
rect 1659 1283 1663 1339
rect 1599 1279 1663 1283
rect 1679 1339 1743 1343
rect 1679 1283 1683 1339
rect 1683 1283 1739 1339
rect 1739 1283 1743 1339
rect 1679 1279 1743 1283
rect 1759 1339 1823 1343
rect 1759 1283 1763 1339
rect 1763 1283 1819 1339
rect 1819 1283 1823 1339
rect 1759 1279 1823 1283
rect 1839 1339 1903 1343
rect 1839 1283 1843 1339
rect 1843 1283 1899 1339
rect 1899 1283 1903 1339
rect 1839 1279 1903 1283
rect 1919 1339 1983 1343
rect 1919 1283 1923 1339
rect 1923 1283 1979 1339
rect 1979 1283 1983 1339
rect 1919 1279 1983 1283
rect 1999 1339 2063 1343
rect 1999 1283 2003 1339
rect 2003 1283 2059 1339
rect 2059 1283 2063 1339
rect 1999 1279 2063 1283
rect 2079 1339 2143 1343
rect 2079 1283 2083 1339
rect 2083 1283 2139 1339
rect 2139 1283 2143 1339
rect 2079 1279 2143 1283
rect 2159 1339 2223 1343
rect 2159 1283 2163 1339
rect 2163 1283 2219 1339
rect 2219 1283 2223 1339
rect 2159 1279 2223 1283
rect 2239 1339 2303 1343
rect 2239 1283 2243 1339
rect 2243 1283 2299 1339
rect 2299 1283 2303 1339
rect 2239 1279 2303 1283
rect 2319 1339 2383 1343
rect 2319 1283 2323 1339
rect 2323 1283 2379 1339
rect 2379 1283 2383 1339
rect 2319 1279 2383 1283
rect 2399 1339 2463 1343
rect 2399 1283 2403 1339
rect 2403 1283 2459 1339
rect 2459 1283 2463 1339
rect 2399 1279 2463 1283
rect 2479 1339 2543 1343
rect 2479 1283 2483 1339
rect 2483 1283 2539 1339
rect 2539 1283 2543 1339
rect 2479 1279 2543 1283
rect 2559 1339 2623 1343
rect 2559 1283 2563 1339
rect 2563 1283 2619 1339
rect 2619 1283 2623 1339
rect 2559 1279 2623 1283
rect 2639 1339 2703 1343
rect 2639 1283 2643 1339
rect 2643 1283 2699 1339
rect 2699 1283 2703 1339
rect 2639 1279 2703 1283
rect 2719 1339 2783 1343
rect 2719 1283 2723 1339
rect 2723 1283 2779 1339
rect 2779 1283 2783 1339
rect 2719 1279 2783 1283
rect 2799 1339 2863 1343
rect 2799 1283 2803 1339
rect 2803 1283 2859 1339
rect 2859 1283 2863 1339
rect 2799 1279 2863 1283
rect 2879 1339 2943 1343
rect 2879 1283 2883 1339
rect 2883 1283 2939 1339
rect 2939 1283 2943 1339
rect 2879 1279 2943 1283
rect 2959 1339 3023 1343
rect 2959 1283 2963 1339
rect 2963 1283 3019 1339
rect 3019 1283 3023 1339
rect 2959 1279 3023 1283
rect 3039 1339 3103 1343
rect 3039 1283 3043 1339
rect 3043 1283 3099 1339
rect 3099 1283 3103 1339
rect 3039 1279 3103 1283
rect 3119 1339 3183 1343
rect 3119 1283 3123 1339
rect 3123 1283 3179 1339
rect 3179 1283 3183 1339
rect 3119 1279 3183 1283
rect -661 405 -357 485
rect -661 349 -626 405
rect -626 349 -570 405
rect -570 349 -546 405
rect -546 349 -490 405
rect -490 349 -466 405
rect -466 349 -410 405
rect -410 349 -386 405
rect -386 349 -357 405
rect -661 341 -357 349
rect 4006 687 4230 728
rect 4006 231 4009 687
rect 4009 231 4225 687
rect 4225 231 4230 687
rect 4006 184 4230 231
rect 45 -592 109 -588
rect 45 -648 49 -592
rect 49 -648 105 -592
rect 105 -648 109 -592
rect 45 -652 109 -648
rect 125 -592 189 -588
rect 125 -648 129 -592
rect 129 -648 185 -592
rect 185 -648 189 -592
rect 125 -652 189 -648
rect 205 -592 269 -588
rect 205 -648 209 -592
rect 209 -648 265 -592
rect 265 -648 269 -592
rect 205 -652 269 -648
rect 285 -592 349 -588
rect 285 -648 289 -592
rect 289 -648 345 -592
rect 345 -648 349 -592
rect 285 -652 349 -648
rect 365 -592 429 -588
rect 365 -648 369 -592
rect 369 -648 425 -592
rect 425 -648 429 -592
rect 365 -652 429 -648
rect 445 -592 509 -588
rect 445 -648 449 -592
rect 449 -648 505 -592
rect 505 -648 509 -592
rect 445 -652 509 -648
rect 525 -592 589 -588
rect 525 -648 529 -592
rect 529 -648 585 -592
rect 585 -648 589 -592
rect 525 -652 589 -648
rect 605 -592 669 -588
rect 605 -648 609 -592
rect 609 -648 665 -592
rect 665 -648 669 -592
rect 605 -652 669 -648
rect 685 -592 749 -588
rect 685 -648 689 -592
rect 689 -648 745 -592
rect 745 -648 749 -592
rect 685 -652 749 -648
rect 765 -592 829 -588
rect 765 -648 769 -592
rect 769 -648 825 -592
rect 825 -648 829 -592
rect 765 -652 829 -648
rect 845 -592 909 -588
rect 845 -648 849 -592
rect 849 -648 905 -592
rect 905 -648 909 -592
rect 845 -652 909 -648
rect 925 -592 989 -588
rect 925 -648 929 -592
rect 929 -648 985 -592
rect 985 -648 989 -592
rect 925 -652 989 -648
rect 1005 -592 1069 -588
rect 1005 -648 1009 -592
rect 1009 -648 1065 -592
rect 1065 -648 1069 -592
rect 1005 -652 1069 -648
rect 1085 -592 1149 -588
rect 1085 -648 1089 -592
rect 1089 -648 1145 -592
rect 1145 -648 1149 -592
rect 1085 -652 1149 -648
rect 1165 -592 1229 -588
rect 1165 -648 1169 -592
rect 1169 -648 1225 -592
rect 1225 -648 1229 -592
rect 1165 -652 1229 -648
rect 1245 -592 1309 -588
rect 1245 -648 1249 -592
rect 1249 -648 1305 -592
rect 1305 -648 1309 -592
rect 1245 -652 1309 -648
rect 1325 -592 1389 -588
rect 1325 -648 1329 -592
rect 1329 -648 1385 -592
rect 1385 -648 1389 -592
rect 1325 -652 1389 -648
rect 1405 -592 1469 -588
rect 1405 -648 1409 -592
rect 1409 -648 1465 -592
rect 1465 -648 1469 -592
rect 1405 -652 1469 -648
rect 1485 -592 1549 -588
rect 1485 -648 1489 -592
rect 1489 -648 1545 -592
rect 1545 -648 1549 -592
rect 1485 -652 1549 -648
rect 1565 -592 1629 -588
rect 1565 -648 1569 -592
rect 1569 -648 1625 -592
rect 1625 -648 1629 -592
rect 1565 -652 1629 -648
rect 1645 -592 1709 -588
rect 1645 -648 1649 -592
rect 1649 -648 1705 -592
rect 1705 -648 1709 -592
rect 1645 -652 1709 -648
rect 1725 -592 1789 -588
rect 1725 -648 1729 -592
rect 1729 -648 1785 -592
rect 1785 -648 1789 -592
rect 1725 -652 1789 -648
rect 1805 -592 1869 -588
rect 1805 -648 1809 -592
rect 1809 -648 1865 -592
rect 1865 -648 1869 -592
rect 1805 -652 1869 -648
rect 1885 -592 1949 -588
rect 1885 -648 1889 -592
rect 1889 -648 1945 -592
rect 1945 -648 1949 -592
rect 1885 -652 1949 -648
rect 1965 -592 2029 -588
rect 1965 -648 1969 -592
rect 1969 -648 2025 -592
rect 2025 -648 2029 -592
rect 1965 -652 2029 -648
rect 2045 -592 2109 -588
rect 2045 -648 2049 -592
rect 2049 -648 2105 -592
rect 2105 -648 2109 -592
rect 2045 -652 2109 -648
rect 2125 -592 2189 -588
rect 2125 -648 2129 -592
rect 2129 -648 2185 -592
rect 2185 -648 2189 -592
rect 2125 -652 2189 -648
rect 2205 -592 2269 -588
rect 2205 -648 2209 -592
rect 2209 -648 2265 -592
rect 2265 -648 2269 -592
rect 2205 -652 2269 -648
rect 2285 -592 2349 -588
rect 2285 -648 2289 -592
rect 2289 -648 2345 -592
rect 2345 -648 2349 -592
rect 2285 -652 2349 -648
rect 2365 -592 2429 -588
rect 2365 -648 2369 -592
rect 2369 -648 2425 -592
rect 2425 -648 2429 -592
rect 2365 -652 2429 -648
rect 2445 -592 2509 -588
rect 2445 -648 2449 -592
rect 2449 -648 2505 -592
rect 2505 -648 2509 -592
rect 2445 -652 2509 -648
rect 2525 -592 2589 -588
rect 2525 -648 2529 -592
rect 2529 -648 2585 -592
rect 2585 -648 2589 -592
rect 2525 -652 2589 -648
rect 2605 -592 2669 -588
rect 2605 -648 2609 -592
rect 2609 -648 2665 -592
rect 2665 -648 2669 -592
rect 2605 -652 2669 -648
rect 2685 -592 2749 -588
rect 2685 -648 2689 -592
rect 2689 -648 2745 -592
rect 2745 -648 2749 -592
rect 2685 -652 2749 -648
rect 2765 -592 2829 -588
rect 2765 -648 2769 -592
rect 2769 -648 2825 -592
rect 2825 -648 2829 -592
rect 2765 -652 2829 -648
rect 2845 -592 2909 -588
rect 2845 -648 2849 -592
rect 2849 -648 2905 -592
rect 2905 -648 2909 -592
rect 2845 -652 2909 -648
rect 2925 -592 2989 -588
rect 2925 -648 2929 -592
rect 2929 -648 2985 -592
rect 2985 -648 2989 -592
rect 2925 -652 2989 -648
rect 3005 -592 3069 -588
rect 3005 -648 3009 -592
rect 3009 -648 3065 -592
rect 3065 -648 3069 -592
rect 3005 -652 3069 -648
<< metal4 >>
rect 158 1526 3184 1538
rect 158 1422 273 1526
rect 114 1343 273 1422
rect 509 1343 593 1526
rect 829 1343 913 1526
rect 1149 1343 1233 1526
rect 1469 1343 1553 1526
rect 1789 1343 1873 1526
rect 2109 1343 2193 1526
rect 2429 1343 2513 1526
rect 2749 1343 2833 1526
rect 3069 1422 3184 1526
rect 3069 1343 3232 1422
rect 114 1279 159 1343
rect 223 1279 239 1343
rect 303 1279 319 1290
rect 383 1279 399 1290
rect 463 1279 479 1290
rect 543 1279 559 1343
rect 623 1279 639 1290
rect 703 1279 719 1290
rect 783 1279 799 1290
rect 863 1279 879 1343
rect 943 1279 959 1290
rect 1023 1279 1039 1290
rect 1103 1279 1119 1290
rect 1183 1279 1199 1343
rect 1263 1279 1279 1290
rect 1343 1279 1359 1290
rect 1423 1279 1439 1290
rect 1503 1279 1519 1343
rect 1583 1279 1599 1290
rect 1663 1279 1679 1290
rect 1743 1279 1759 1290
rect 1823 1279 1839 1343
rect 1903 1279 1919 1290
rect 1983 1279 1999 1290
rect 2063 1279 2079 1290
rect 2143 1279 2159 1343
rect 2223 1279 2239 1290
rect 2303 1279 2319 1290
rect 2383 1279 2399 1290
rect 2463 1279 2479 1343
rect 2543 1279 2559 1290
rect 2623 1279 2639 1290
rect 2703 1279 2719 1290
rect 2783 1279 2799 1343
rect 2863 1279 2879 1290
rect 2943 1279 2959 1290
rect 3023 1279 3039 1290
rect 3103 1279 3119 1343
rect 3183 1279 3232 1343
rect 114 1244 3232 1279
rect 3856 739 4362 898
rect -846 511 -232 626
rect -846 275 -667 511
rect -431 485 -232 511
rect -357 341 -232 485
rect -431 275 -232 341
rect -846 160 -232 275
rect 3856 503 3989 739
rect 4225 728 4362 739
rect 3856 419 4006 503
rect 3856 183 3989 419
rect 4230 184 4362 728
rect 4225 183 4362 184
rect 3856 30 4362 183
rect 44 -405 3070 -392
rect 44 -508 159 -405
rect 0 -588 159 -508
rect 395 -588 479 -405
rect 715 -588 799 -405
rect 1035 -588 1119 -405
rect 1355 -588 1439 -405
rect 1675 -588 1759 -405
rect 1995 -588 2079 -405
rect 2315 -588 2399 -405
rect 2635 -588 2719 -405
rect 2955 -508 3070 -405
rect 2955 -588 3118 -508
rect 0 -652 45 -588
rect 109 -652 125 -588
rect 189 -652 205 -641
rect 269 -652 285 -641
rect 349 -652 365 -641
rect 429 -652 445 -588
rect 509 -652 525 -641
rect 589 -652 605 -641
rect 669 -652 685 -641
rect 749 -652 765 -588
rect 829 -652 845 -641
rect 909 -652 925 -641
rect 989 -652 1005 -641
rect 1069 -652 1085 -588
rect 1149 -652 1165 -641
rect 1229 -652 1245 -641
rect 1309 -652 1325 -641
rect 1389 -652 1405 -588
rect 1469 -652 1485 -641
rect 1549 -652 1565 -641
rect 1629 -652 1645 -641
rect 1709 -652 1725 -588
rect 1789 -652 1805 -641
rect 1869 -652 1885 -641
rect 1949 -652 1965 -641
rect 2029 -652 2045 -588
rect 2109 -652 2125 -641
rect 2189 -652 2205 -641
rect 2269 -652 2285 -641
rect 2349 -652 2365 -588
rect 2429 -652 2445 -641
rect 2509 -652 2525 -641
rect 2589 -652 2605 -641
rect 2669 -652 2685 -588
rect 2749 -652 2765 -641
rect 2829 -652 2845 -641
rect 2909 -652 2925 -641
rect 2989 -652 3005 -588
rect 3069 -652 3118 -588
rect 0 -686 3118 -652
<< via4 >>
rect 273 1343 509 1526
rect 593 1343 829 1526
rect 913 1343 1149 1526
rect 1233 1343 1469 1526
rect 1553 1343 1789 1526
rect 1873 1343 2109 1526
rect 2193 1343 2429 1526
rect 2513 1343 2749 1526
rect 2833 1343 3069 1526
rect 273 1290 303 1343
rect 303 1290 319 1343
rect 319 1290 383 1343
rect 383 1290 399 1343
rect 399 1290 463 1343
rect 463 1290 479 1343
rect 479 1290 509 1343
rect 593 1290 623 1343
rect 623 1290 639 1343
rect 639 1290 703 1343
rect 703 1290 719 1343
rect 719 1290 783 1343
rect 783 1290 799 1343
rect 799 1290 829 1343
rect 913 1290 943 1343
rect 943 1290 959 1343
rect 959 1290 1023 1343
rect 1023 1290 1039 1343
rect 1039 1290 1103 1343
rect 1103 1290 1119 1343
rect 1119 1290 1149 1343
rect 1233 1290 1263 1343
rect 1263 1290 1279 1343
rect 1279 1290 1343 1343
rect 1343 1290 1359 1343
rect 1359 1290 1423 1343
rect 1423 1290 1439 1343
rect 1439 1290 1469 1343
rect 1553 1290 1583 1343
rect 1583 1290 1599 1343
rect 1599 1290 1663 1343
rect 1663 1290 1679 1343
rect 1679 1290 1743 1343
rect 1743 1290 1759 1343
rect 1759 1290 1789 1343
rect 1873 1290 1903 1343
rect 1903 1290 1919 1343
rect 1919 1290 1983 1343
rect 1983 1290 1999 1343
rect 1999 1290 2063 1343
rect 2063 1290 2079 1343
rect 2079 1290 2109 1343
rect 2193 1290 2223 1343
rect 2223 1290 2239 1343
rect 2239 1290 2303 1343
rect 2303 1290 2319 1343
rect 2319 1290 2383 1343
rect 2383 1290 2399 1343
rect 2399 1290 2429 1343
rect 2513 1290 2543 1343
rect 2543 1290 2559 1343
rect 2559 1290 2623 1343
rect 2623 1290 2639 1343
rect 2639 1290 2703 1343
rect 2703 1290 2719 1343
rect 2719 1290 2749 1343
rect 2833 1290 2863 1343
rect 2863 1290 2879 1343
rect 2879 1290 2943 1343
rect 2943 1290 2959 1343
rect 2959 1290 3023 1343
rect 3023 1290 3039 1343
rect 3039 1290 3069 1343
rect -667 485 -431 511
rect -667 341 -661 485
rect -661 341 -431 485
rect -667 275 -431 341
rect 3989 728 4225 739
rect 3989 503 4006 728
rect 4006 503 4225 728
rect 3989 184 4006 419
rect 4006 184 4225 419
rect 3989 183 4225 184
rect 159 -588 395 -405
rect 479 -588 715 -405
rect 799 -588 1035 -405
rect 1119 -588 1355 -405
rect 1439 -588 1675 -405
rect 1759 -588 1995 -405
rect 2079 -588 2315 -405
rect 2399 -588 2635 -405
rect 2719 -588 2955 -405
rect 159 -641 189 -588
rect 189 -641 205 -588
rect 205 -641 269 -588
rect 269 -641 285 -588
rect 285 -641 349 -588
rect 349 -641 365 -588
rect 365 -641 395 -588
rect 479 -641 509 -588
rect 509 -641 525 -588
rect 525 -641 589 -588
rect 589 -641 605 -588
rect 605 -641 669 -588
rect 669 -641 685 -588
rect 685 -641 715 -588
rect 799 -641 829 -588
rect 829 -641 845 -588
rect 845 -641 909 -588
rect 909 -641 925 -588
rect 925 -641 989 -588
rect 989 -641 1005 -588
rect 1005 -641 1035 -588
rect 1119 -641 1149 -588
rect 1149 -641 1165 -588
rect 1165 -641 1229 -588
rect 1229 -641 1245 -588
rect 1245 -641 1309 -588
rect 1309 -641 1325 -588
rect 1325 -641 1355 -588
rect 1439 -641 1469 -588
rect 1469 -641 1485 -588
rect 1485 -641 1549 -588
rect 1549 -641 1565 -588
rect 1565 -641 1629 -588
rect 1629 -641 1645 -588
rect 1645 -641 1675 -588
rect 1759 -641 1789 -588
rect 1789 -641 1805 -588
rect 1805 -641 1869 -588
rect 1869 -641 1885 -588
rect 1885 -641 1949 -588
rect 1949 -641 1965 -588
rect 1965 -641 1995 -588
rect 2079 -641 2109 -588
rect 2109 -641 2125 -588
rect 2125 -641 2189 -588
rect 2189 -641 2205 -588
rect 2205 -641 2269 -588
rect 2269 -641 2285 -588
rect 2285 -641 2315 -588
rect 2399 -641 2429 -588
rect 2429 -641 2445 -588
rect 2445 -641 2509 -588
rect 2509 -641 2525 -588
rect 2525 -641 2589 -588
rect 2589 -641 2605 -588
rect 2605 -641 2635 -588
rect 2719 -641 2749 -588
rect 2749 -641 2765 -588
rect 2765 -641 2829 -588
rect 2829 -641 2845 -588
rect 2845 -641 2909 -588
rect 2909 -641 2925 -588
rect 2925 -641 2955 -588
<< metal5 >>
rect 114 1526 3606 1644
rect 114 1290 273 1526
rect 509 1290 593 1526
rect 829 1290 913 1526
rect 1149 1290 1233 1526
rect 1469 1290 1553 1526
rect 1789 1290 1873 1526
rect 2109 1290 2193 1526
rect 2429 1290 2513 1526
rect 2749 1290 2833 1526
rect 3069 1290 3606 1526
rect 114 1244 3606 1290
rect 3810 739 4384 950
rect -918 511 -214 706
rect -918 275 -667 511
rect -431 275 -214 511
rect -918 134 -214 275
rect 3810 503 3989 739
rect 4225 503 4384 739
rect 3810 419 4384 503
rect 3810 183 3989 419
rect 4225 183 4384 419
rect 3810 -38 4384 183
rect 0 -405 3492 -288
rect 0 -641 159 -405
rect 395 -641 479 -405
rect 715 -641 799 -405
rect 1035 -641 1119 -405
rect 1355 -641 1439 -405
rect 1675 -641 1759 -405
rect 1995 -641 2079 -405
rect 2315 -641 2399 -405
rect 2635 -641 2719 -405
rect 2955 -641 3492 -405
rect 0 -686 3492 -641
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1611881054
transform 1 0 464 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_0
timestamp 1611881054
transform 1 0 0 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1611881054
transform 1 0 536 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1611881054
transform 1 0 888 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1611881054
transform 1 0 1592 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1611881054
transform 1 0 1240 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1611881054
transform 1 0 1944 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1611881054
transform 1 0 2648 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1611881054
transform 1 0 2296 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1611881054
transform 1 0 3000 0 1 0
box -38 -48 130 592
<< labels >>
rlabel metal2 s 480 532 486 536 4 Vdd
port 1 nsew
rlabel metal1 s 480 -4 486 0 4 Gnd
port 2 nsew
rlabel metal1 s -96 226 -90 230 4 en
port 3 nsew
rlabel metal1 s -84 342 -70 362 4 out
port 4 nsew
<< end >>
