magic
tech sky130A
magscale 1 2
timestamp 1607987969
<< error_p >>
rect -365 122 -307 128
rect -173 122 -115 128
rect 19 122 77 128
rect 211 122 269 128
rect 403 122 461 128
rect -365 88 -353 122
rect -173 88 -161 122
rect 19 88 31 122
rect 211 88 223 122
rect 403 88 415 122
rect -365 82 -307 88
rect -173 82 -115 88
rect 19 82 77 88
rect 211 82 269 88
rect 403 82 461 88
rect -461 -88 -403 -82
rect -269 -88 -211 -82
rect -77 -88 -19 -82
rect 115 -88 173 -82
rect 307 -88 365 -82
rect -461 -122 -449 -88
rect -269 -122 -257 -88
rect -77 -122 -65 -88
rect 115 -122 127 -88
rect 307 -122 319 -88
rect -461 -128 -403 -122
rect -269 -128 -211 -122
rect -77 -128 -19 -122
rect 115 -128 173 -122
rect 307 -128 365 -122
<< pwell >>
rect -647 -260 647 260
<< nmoslvt >>
rect -447 -50 -417 50
rect -351 -50 -321 50
rect -255 -50 -225 50
rect -159 -50 -129 50
rect -63 -50 -33 50
rect 33 -50 63 50
rect 129 -50 159 50
rect 225 -50 255 50
rect 321 -50 351 50
rect 417 -50 447 50
<< ndiff >>
rect -509 38 -447 50
rect -509 -38 -497 38
rect -463 -38 -447 38
rect -509 -50 -447 -38
rect -417 38 -351 50
rect -417 -38 -401 38
rect -367 -38 -351 38
rect -417 -50 -351 -38
rect -321 38 -255 50
rect -321 -38 -305 38
rect -271 -38 -255 38
rect -321 -50 -255 -38
rect -225 38 -159 50
rect -225 -38 -209 38
rect -175 -38 -159 38
rect -225 -50 -159 -38
rect -129 38 -63 50
rect -129 -38 -113 38
rect -79 -38 -63 38
rect -129 -50 -63 -38
rect -33 38 33 50
rect -33 -38 -17 38
rect 17 -38 33 38
rect -33 -50 33 -38
rect 63 38 129 50
rect 63 -38 79 38
rect 113 -38 129 38
rect 63 -50 129 -38
rect 159 38 225 50
rect 159 -38 175 38
rect 209 -38 225 38
rect 159 -50 225 -38
rect 255 38 321 50
rect 255 -38 271 38
rect 305 -38 321 38
rect 255 -50 321 -38
rect 351 38 417 50
rect 351 -38 367 38
rect 401 -38 417 38
rect 351 -50 417 -38
rect 447 38 509 50
rect 447 -38 463 38
rect 497 -38 509 38
rect 447 -50 509 -38
<< ndiffc >>
rect -497 -38 -463 38
rect -401 -38 -367 38
rect -305 -38 -271 38
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect 271 -38 305 38
rect 367 -38 401 38
rect 463 -38 497 38
<< psubdiff >>
rect -611 190 -515 224
rect 515 190 611 224
rect -611 128 -577 190
rect 577 128 611 190
rect -611 -190 -577 -128
rect 577 -190 611 -128
rect -611 -224 -515 -190
rect 515 -224 611 -190
<< psubdiffcont >>
rect -515 190 515 224
rect -611 -128 -577 128
rect 577 -128 611 128
rect -515 -224 515 -190
<< poly >>
rect -369 122 -303 138
rect -369 88 -353 122
rect -319 88 -303 122
rect -447 50 -417 76
rect -369 72 -303 88
rect -177 122 -111 138
rect -177 88 -161 122
rect -127 88 -111 122
rect -351 50 -321 72
rect -255 50 -225 76
rect -177 72 -111 88
rect 15 122 81 138
rect 15 88 31 122
rect 65 88 81 122
rect -159 50 -129 72
rect -63 50 -33 76
rect 15 72 81 88
rect 207 122 273 138
rect 207 88 223 122
rect 257 88 273 122
rect 33 50 63 72
rect 129 50 159 76
rect 207 72 273 88
rect 399 122 465 138
rect 399 88 415 122
rect 449 88 465 122
rect 225 50 255 72
rect 321 50 351 76
rect 399 72 465 88
rect 417 50 447 72
rect -447 -72 -417 -50
rect -465 -88 -399 -72
rect -351 -76 -321 -50
rect -255 -72 -225 -50
rect -465 -122 -449 -88
rect -415 -122 -399 -88
rect -465 -138 -399 -122
rect -273 -88 -207 -72
rect -159 -76 -129 -50
rect -63 -72 -33 -50
rect -273 -122 -257 -88
rect -223 -122 -207 -88
rect -273 -138 -207 -122
rect -81 -88 -15 -72
rect 33 -76 63 -50
rect 129 -72 159 -50
rect -81 -122 -65 -88
rect -31 -122 -15 -88
rect -81 -138 -15 -122
rect 111 -88 177 -72
rect 225 -76 255 -50
rect 321 -72 351 -50
rect 111 -122 127 -88
rect 161 -122 177 -88
rect 111 -138 177 -122
rect 303 -88 369 -72
rect 417 -76 447 -50
rect 303 -122 319 -88
rect 353 -122 369 -88
rect 303 -138 369 -122
<< polycont >>
rect -353 88 -319 122
rect -161 88 -127 122
rect 31 88 65 122
rect 223 88 257 122
rect 415 88 449 122
rect -449 -122 -415 -88
rect -257 -122 -223 -88
rect -65 -122 -31 -88
rect 127 -122 161 -88
rect 319 -122 353 -88
<< locali >>
rect -611 190 -515 224
rect 515 190 611 224
rect -611 128 -577 190
rect 577 128 611 190
rect -369 88 -353 122
rect -319 88 -303 122
rect -177 88 -161 122
rect -127 88 -111 122
rect 15 88 31 122
rect 65 88 81 122
rect 207 88 223 122
rect 257 88 273 122
rect 399 88 415 122
rect 449 88 465 122
rect -497 38 -463 54
rect -497 -54 -463 -38
rect -401 38 -367 54
rect -401 -54 -367 -38
rect -305 38 -271 54
rect -305 -54 -271 -38
rect -209 38 -175 54
rect -209 -54 -175 -38
rect -113 38 -79 54
rect -113 -54 -79 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 79 38 113 54
rect 79 -54 113 -38
rect 175 38 209 54
rect 175 -54 209 -38
rect 271 38 305 54
rect 271 -54 305 -38
rect 367 38 401 54
rect 367 -54 401 -38
rect 463 38 497 54
rect 463 -54 497 -38
rect -465 -122 -449 -88
rect -415 -122 -399 -88
rect -273 -122 -257 -88
rect -223 -122 -207 -88
rect -81 -122 -65 -88
rect -31 -122 -15 -88
rect 111 -122 127 -88
rect 161 -122 177 -88
rect 303 -122 319 -88
rect 353 -122 369 -88
rect -611 -224 -577 -128
rect 577 -224 611 -128
<< viali >>
rect -353 88 -319 122
rect -161 88 -127 122
rect 31 88 65 122
rect 223 88 257 122
rect 415 88 449 122
rect -497 -38 -463 38
rect -401 -38 -367 38
rect -305 -38 -271 38
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect 271 -38 305 38
rect 367 -38 401 38
rect 463 -38 497 38
rect -449 -122 -415 -88
rect -257 -122 -223 -88
rect -65 -122 -31 -88
rect 127 -122 161 -88
rect 319 -122 353 -88
rect -577 -224 -515 -190
rect -515 -224 515 -190
rect 515 -224 577 -190
<< metal1 >>
rect -365 122 -307 128
rect -365 88 -353 122
rect -319 88 -307 122
rect -365 82 -307 88
rect -173 122 -115 128
rect -173 88 -161 122
rect -127 88 -115 122
rect -173 82 -115 88
rect 19 122 77 128
rect 19 88 31 122
rect 65 88 77 122
rect 19 82 77 88
rect 211 122 269 128
rect 211 88 223 122
rect 257 88 269 122
rect 211 82 269 88
rect 403 122 461 128
rect 403 88 415 122
rect 449 88 461 122
rect 403 82 461 88
rect -503 38 -457 50
rect -503 -38 -497 38
rect -463 -38 -457 38
rect -503 -50 -457 -38
rect -407 38 -361 50
rect -407 -38 -401 38
rect -367 -38 -361 38
rect -407 -50 -361 -38
rect -311 38 -265 50
rect -311 -38 -305 38
rect -271 -38 -265 38
rect -311 -50 -265 -38
rect -215 38 -169 50
rect -215 -38 -209 38
rect -175 -38 -169 38
rect -215 -50 -169 -38
rect -119 38 -73 50
rect -119 -38 -113 38
rect -79 -38 -73 38
rect -119 -50 -73 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 73 38 119 50
rect 73 -38 79 38
rect 113 -38 119 38
rect 73 -50 119 -38
rect 169 38 215 50
rect 169 -38 175 38
rect 209 -38 215 38
rect 169 -50 215 -38
rect 265 38 311 50
rect 265 -38 271 38
rect 305 -38 311 38
rect 265 -50 311 -38
rect 361 38 407 50
rect 361 -38 367 38
rect 401 -38 407 38
rect 361 -50 407 -38
rect 457 38 503 50
rect 457 -38 463 38
rect 497 -38 503 38
rect 457 -50 503 -38
rect -461 -88 -403 -82
rect -461 -122 -449 -88
rect -415 -122 -403 -88
rect -461 -128 -403 -122
rect -269 -88 -211 -82
rect -269 -122 -257 -88
rect -223 -122 -211 -88
rect -269 -128 -211 -122
rect -77 -88 -19 -82
rect -77 -122 -65 -88
rect -31 -122 -19 -88
rect -77 -128 -19 -122
rect 115 -88 173 -82
rect 115 -122 127 -88
rect 161 -122 173 -88
rect 115 -128 173 -122
rect 307 -88 365 -82
rect 307 -122 319 -88
rect 353 -122 365 -88
rect 307 -128 365 -122
rect -589 -190 589 -184
rect -589 -224 -577 -190
rect 577 -224 589 -190
rect -589 -230 589 -224
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -594 -207 594 207
string parameters w 0.5 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
