magic
tech sky130A
timestamp 1606545195
<< nwell >>
rect -348 -484 348 484
<< pmoslvt >>
rect -250 -375 250 375
<< pdiff >>
rect -279 369 -250 375
rect -279 -369 -273 369
rect -256 -369 -250 369
rect -279 -375 -250 -369
rect 250 369 279 375
rect 250 -369 256 369
rect 273 -369 279 369
rect 250 -375 279 -369
<< pdiffc >>
rect -273 -369 -256 369
rect 256 -369 273 369
<< nsubdiff >>
rect -330 449 -282 466
rect 282 449 330 466
rect -330 418 -313 449
rect 313 418 330 449
rect -330 -449 -313 -418
rect 313 -449 330 -418
rect -330 -466 -282 -449
rect 282 -466 330 -449
<< nsubdiffcont >>
rect -282 449 282 466
rect -330 -418 -313 418
rect 313 -418 330 418
rect -282 -466 282 -449
<< poly >>
rect -250 415 250 423
rect -250 398 -242 415
rect 242 398 250 415
rect -250 375 250 398
rect -250 -398 250 -375
rect -250 -415 -242 -398
rect 242 -415 250 -398
rect -250 -423 250 -415
<< polycont >>
rect -242 398 242 415
rect -242 -415 242 -398
<< locali >>
rect -330 449 -282 466
rect 282 449 330 466
rect -330 418 -313 449
rect 313 418 330 449
rect -250 398 -242 415
rect 242 398 250 415
rect -273 369 -256 377
rect -273 -377 -256 -369
rect 256 369 273 377
rect 256 -377 273 -369
rect -250 -415 -242 -398
rect 242 -415 250 -398
rect -330 -449 -313 -418
rect 313 -449 330 -418
rect -330 -466 -282 -449
rect 282 -466 330 -449
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -321 -458 321 458
string parameters w 7.5 l 5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
