magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -1734 840 1734 874
rect -1734 -840 -1700 840
rect 1700 -840 1734 840
rect -1734 -874 1734 -840
<< nmos >>
rect -1574 -700 -1174 700
rect -1116 -700 -716 700
rect -658 -700 -258 700
rect -200 -700 200 700
rect 258 -700 658 700
rect 716 -700 1116 700
rect 1174 -700 1574 700
<< ndiff >>
rect -1632 663 -1574 700
rect -1632 629 -1620 663
rect -1586 629 -1574 663
rect -1632 595 -1574 629
rect -1632 561 -1620 595
rect -1586 561 -1574 595
rect -1632 527 -1574 561
rect -1632 493 -1620 527
rect -1586 493 -1574 527
rect -1632 459 -1574 493
rect -1632 425 -1620 459
rect -1586 425 -1574 459
rect -1632 391 -1574 425
rect -1632 357 -1620 391
rect -1586 357 -1574 391
rect -1632 323 -1574 357
rect -1632 289 -1620 323
rect -1586 289 -1574 323
rect -1632 255 -1574 289
rect -1632 221 -1620 255
rect -1586 221 -1574 255
rect -1632 187 -1574 221
rect -1632 153 -1620 187
rect -1586 153 -1574 187
rect -1632 119 -1574 153
rect -1632 85 -1620 119
rect -1586 85 -1574 119
rect -1632 51 -1574 85
rect -1632 17 -1620 51
rect -1586 17 -1574 51
rect -1632 -17 -1574 17
rect -1632 -51 -1620 -17
rect -1586 -51 -1574 -17
rect -1632 -85 -1574 -51
rect -1632 -119 -1620 -85
rect -1586 -119 -1574 -85
rect -1632 -153 -1574 -119
rect -1632 -187 -1620 -153
rect -1586 -187 -1574 -153
rect -1632 -221 -1574 -187
rect -1632 -255 -1620 -221
rect -1586 -255 -1574 -221
rect -1632 -289 -1574 -255
rect -1632 -323 -1620 -289
rect -1586 -323 -1574 -289
rect -1632 -357 -1574 -323
rect -1632 -391 -1620 -357
rect -1586 -391 -1574 -357
rect -1632 -425 -1574 -391
rect -1632 -459 -1620 -425
rect -1586 -459 -1574 -425
rect -1632 -493 -1574 -459
rect -1632 -527 -1620 -493
rect -1586 -527 -1574 -493
rect -1632 -561 -1574 -527
rect -1632 -595 -1620 -561
rect -1586 -595 -1574 -561
rect -1632 -629 -1574 -595
rect -1632 -663 -1620 -629
rect -1586 -663 -1574 -629
rect -1632 -700 -1574 -663
rect -1174 663 -1116 700
rect -1174 629 -1162 663
rect -1128 629 -1116 663
rect -1174 595 -1116 629
rect -1174 561 -1162 595
rect -1128 561 -1116 595
rect -1174 527 -1116 561
rect -1174 493 -1162 527
rect -1128 493 -1116 527
rect -1174 459 -1116 493
rect -1174 425 -1162 459
rect -1128 425 -1116 459
rect -1174 391 -1116 425
rect -1174 357 -1162 391
rect -1128 357 -1116 391
rect -1174 323 -1116 357
rect -1174 289 -1162 323
rect -1128 289 -1116 323
rect -1174 255 -1116 289
rect -1174 221 -1162 255
rect -1128 221 -1116 255
rect -1174 187 -1116 221
rect -1174 153 -1162 187
rect -1128 153 -1116 187
rect -1174 119 -1116 153
rect -1174 85 -1162 119
rect -1128 85 -1116 119
rect -1174 51 -1116 85
rect -1174 17 -1162 51
rect -1128 17 -1116 51
rect -1174 -17 -1116 17
rect -1174 -51 -1162 -17
rect -1128 -51 -1116 -17
rect -1174 -85 -1116 -51
rect -1174 -119 -1162 -85
rect -1128 -119 -1116 -85
rect -1174 -153 -1116 -119
rect -1174 -187 -1162 -153
rect -1128 -187 -1116 -153
rect -1174 -221 -1116 -187
rect -1174 -255 -1162 -221
rect -1128 -255 -1116 -221
rect -1174 -289 -1116 -255
rect -1174 -323 -1162 -289
rect -1128 -323 -1116 -289
rect -1174 -357 -1116 -323
rect -1174 -391 -1162 -357
rect -1128 -391 -1116 -357
rect -1174 -425 -1116 -391
rect -1174 -459 -1162 -425
rect -1128 -459 -1116 -425
rect -1174 -493 -1116 -459
rect -1174 -527 -1162 -493
rect -1128 -527 -1116 -493
rect -1174 -561 -1116 -527
rect -1174 -595 -1162 -561
rect -1128 -595 -1116 -561
rect -1174 -629 -1116 -595
rect -1174 -663 -1162 -629
rect -1128 -663 -1116 -629
rect -1174 -700 -1116 -663
rect -716 663 -658 700
rect -716 629 -704 663
rect -670 629 -658 663
rect -716 595 -658 629
rect -716 561 -704 595
rect -670 561 -658 595
rect -716 527 -658 561
rect -716 493 -704 527
rect -670 493 -658 527
rect -716 459 -658 493
rect -716 425 -704 459
rect -670 425 -658 459
rect -716 391 -658 425
rect -716 357 -704 391
rect -670 357 -658 391
rect -716 323 -658 357
rect -716 289 -704 323
rect -670 289 -658 323
rect -716 255 -658 289
rect -716 221 -704 255
rect -670 221 -658 255
rect -716 187 -658 221
rect -716 153 -704 187
rect -670 153 -658 187
rect -716 119 -658 153
rect -716 85 -704 119
rect -670 85 -658 119
rect -716 51 -658 85
rect -716 17 -704 51
rect -670 17 -658 51
rect -716 -17 -658 17
rect -716 -51 -704 -17
rect -670 -51 -658 -17
rect -716 -85 -658 -51
rect -716 -119 -704 -85
rect -670 -119 -658 -85
rect -716 -153 -658 -119
rect -716 -187 -704 -153
rect -670 -187 -658 -153
rect -716 -221 -658 -187
rect -716 -255 -704 -221
rect -670 -255 -658 -221
rect -716 -289 -658 -255
rect -716 -323 -704 -289
rect -670 -323 -658 -289
rect -716 -357 -658 -323
rect -716 -391 -704 -357
rect -670 -391 -658 -357
rect -716 -425 -658 -391
rect -716 -459 -704 -425
rect -670 -459 -658 -425
rect -716 -493 -658 -459
rect -716 -527 -704 -493
rect -670 -527 -658 -493
rect -716 -561 -658 -527
rect -716 -595 -704 -561
rect -670 -595 -658 -561
rect -716 -629 -658 -595
rect -716 -663 -704 -629
rect -670 -663 -658 -629
rect -716 -700 -658 -663
rect -258 663 -200 700
rect -258 629 -246 663
rect -212 629 -200 663
rect -258 595 -200 629
rect -258 561 -246 595
rect -212 561 -200 595
rect -258 527 -200 561
rect -258 493 -246 527
rect -212 493 -200 527
rect -258 459 -200 493
rect -258 425 -246 459
rect -212 425 -200 459
rect -258 391 -200 425
rect -258 357 -246 391
rect -212 357 -200 391
rect -258 323 -200 357
rect -258 289 -246 323
rect -212 289 -200 323
rect -258 255 -200 289
rect -258 221 -246 255
rect -212 221 -200 255
rect -258 187 -200 221
rect -258 153 -246 187
rect -212 153 -200 187
rect -258 119 -200 153
rect -258 85 -246 119
rect -212 85 -200 119
rect -258 51 -200 85
rect -258 17 -246 51
rect -212 17 -200 51
rect -258 -17 -200 17
rect -258 -51 -246 -17
rect -212 -51 -200 -17
rect -258 -85 -200 -51
rect -258 -119 -246 -85
rect -212 -119 -200 -85
rect -258 -153 -200 -119
rect -258 -187 -246 -153
rect -212 -187 -200 -153
rect -258 -221 -200 -187
rect -258 -255 -246 -221
rect -212 -255 -200 -221
rect -258 -289 -200 -255
rect -258 -323 -246 -289
rect -212 -323 -200 -289
rect -258 -357 -200 -323
rect -258 -391 -246 -357
rect -212 -391 -200 -357
rect -258 -425 -200 -391
rect -258 -459 -246 -425
rect -212 -459 -200 -425
rect -258 -493 -200 -459
rect -258 -527 -246 -493
rect -212 -527 -200 -493
rect -258 -561 -200 -527
rect -258 -595 -246 -561
rect -212 -595 -200 -561
rect -258 -629 -200 -595
rect -258 -663 -246 -629
rect -212 -663 -200 -629
rect -258 -700 -200 -663
rect 200 663 258 700
rect 200 629 212 663
rect 246 629 258 663
rect 200 595 258 629
rect 200 561 212 595
rect 246 561 258 595
rect 200 527 258 561
rect 200 493 212 527
rect 246 493 258 527
rect 200 459 258 493
rect 200 425 212 459
rect 246 425 258 459
rect 200 391 258 425
rect 200 357 212 391
rect 246 357 258 391
rect 200 323 258 357
rect 200 289 212 323
rect 246 289 258 323
rect 200 255 258 289
rect 200 221 212 255
rect 246 221 258 255
rect 200 187 258 221
rect 200 153 212 187
rect 246 153 258 187
rect 200 119 258 153
rect 200 85 212 119
rect 246 85 258 119
rect 200 51 258 85
rect 200 17 212 51
rect 246 17 258 51
rect 200 -17 258 17
rect 200 -51 212 -17
rect 246 -51 258 -17
rect 200 -85 258 -51
rect 200 -119 212 -85
rect 246 -119 258 -85
rect 200 -153 258 -119
rect 200 -187 212 -153
rect 246 -187 258 -153
rect 200 -221 258 -187
rect 200 -255 212 -221
rect 246 -255 258 -221
rect 200 -289 258 -255
rect 200 -323 212 -289
rect 246 -323 258 -289
rect 200 -357 258 -323
rect 200 -391 212 -357
rect 246 -391 258 -357
rect 200 -425 258 -391
rect 200 -459 212 -425
rect 246 -459 258 -425
rect 200 -493 258 -459
rect 200 -527 212 -493
rect 246 -527 258 -493
rect 200 -561 258 -527
rect 200 -595 212 -561
rect 246 -595 258 -561
rect 200 -629 258 -595
rect 200 -663 212 -629
rect 246 -663 258 -629
rect 200 -700 258 -663
rect 658 663 716 700
rect 658 629 670 663
rect 704 629 716 663
rect 658 595 716 629
rect 658 561 670 595
rect 704 561 716 595
rect 658 527 716 561
rect 658 493 670 527
rect 704 493 716 527
rect 658 459 716 493
rect 658 425 670 459
rect 704 425 716 459
rect 658 391 716 425
rect 658 357 670 391
rect 704 357 716 391
rect 658 323 716 357
rect 658 289 670 323
rect 704 289 716 323
rect 658 255 716 289
rect 658 221 670 255
rect 704 221 716 255
rect 658 187 716 221
rect 658 153 670 187
rect 704 153 716 187
rect 658 119 716 153
rect 658 85 670 119
rect 704 85 716 119
rect 658 51 716 85
rect 658 17 670 51
rect 704 17 716 51
rect 658 -17 716 17
rect 658 -51 670 -17
rect 704 -51 716 -17
rect 658 -85 716 -51
rect 658 -119 670 -85
rect 704 -119 716 -85
rect 658 -153 716 -119
rect 658 -187 670 -153
rect 704 -187 716 -153
rect 658 -221 716 -187
rect 658 -255 670 -221
rect 704 -255 716 -221
rect 658 -289 716 -255
rect 658 -323 670 -289
rect 704 -323 716 -289
rect 658 -357 716 -323
rect 658 -391 670 -357
rect 704 -391 716 -357
rect 658 -425 716 -391
rect 658 -459 670 -425
rect 704 -459 716 -425
rect 658 -493 716 -459
rect 658 -527 670 -493
rect 704 -527 716 -493
rect 658 -561 716 -527
rect 658 -595 670 -561
rect 704 -595 716 -561
rect 658 -629 716 -595
rect 658 -663 670 -629
rect 704 -663 716 -629
rect 658 -700 716 -663
rect 1116 663 1174 700
rect 1116 629 1128 663
rect 1162 629 1174 663
rect 1116 595 1174 629
rect 1116 561 1128 595
rect 1162 561 1174 595
rect 1116 527 1174 561
rect 1116 493 1128 527
rect 1162 493 1174 527
rect 1116 459 1174 493
rect 1116 425 1128 459
rect 1162 425 1174 459
rect 1116 391 1174 425
rect 1116 357 1128 391
rect 1162 357 1174 391
rect 1116 323 1174 357
rect 1116 289 1128 323
rect 1162 289 1174 323
rect 1116 255 1174 289
rect 1116 221 1128 255
rect 1162 221 1174 255
rect 1116 187 1174 221
rect 1116 153 1128 187
rect 1162 153 1174 187
rect 1116 119 1174 153
rect 1116 85 1128 119
rect 1162 85 1174 119
rect 1116 51 1174 85
rect 1116 17 1128 51
rect 1162 17 1174 51
rect 1116 -17 1174 17
rect 1116 -51 1128 -17
rect 1162 -51 1174 -17
rect 1116 -85 1174 -51
rect 1116 -119 1128 -85
rect 1162 -119 1174 -85
rect 1116 -153 1174 -119
rect 1116 -187 1128 -153
rect 1162 -187 1174 -153
rect 1116 -221 1174 -187
rect 1116 -255 1128 -221
rect 1162 -255 1174 -221
rect 1116 -289 1174 -255
rect 1116 -323 1128 -289
rect 1162 -323 1174 -289
rect 1116 -357 1174 -323
rect 1116 -391 1128 -357
rect 1162 -391 1174 -357
rect 1116 -425 1174 -391
rect 1116 -459 1128 -425
rect 1162 -459 1174 -425
rect 1116 -493 1174 -459
rect 1116 -527 1128 -493
rect 1162 -527 1174 -493
rect 1116 -561 1174 -527
rect 1116 -595 1128 -561
rect 1162 -595 1174 -561
rect 1116 -629 1174 -595
rect 1116 -663 1128 -629
rect 1162 -663 1174 -629
rect 1116 -700 1174 -663
rect 1574 663 1632 700
rect 1574 629 1586 663
rect 1620 629 1632 663
rect 1574 595 1632 629
rect 1574 561 1586 595
rect 1620 561 1632 595
rect 1574 527 1632 561
rect 1574 493 1586 527
rect 1620 493 1632 527
rect 1574 459 1632 493
rect 1574 425 1586 459
rect 1620 425 1632 459
rect 1574 391 1632 425
rect 1574 357 1586 391
rect 1620 357 1632 391
rect 1574 323 1632 357
rect 1574 289 1586 323
rect 1620 289 1632 323
rect 1574 255 1632 289
rect 1574 221 1586 255
rect 1620 221 1632 255
rect 1574 187 1632 221
rect 1574 153 1586 187
rect 1620 153 1632 187
rect 1574 119 1632 153
rect 1574 85 1586 119
rect 1620 85 1632 119
rect 1574 51 1632 85
rect 1574 17 1586 51
rect 1620 17 1632 51
rect 1574 -17 1632 17
rect 1574 -51 1586 -17
rect 1620 -51 1632 -17
rect 1574 -85 1632 -51
rect 1574 -119 1586 -85
rect 1620 -119 1632 -85
rect 1574 -153 1632 -119
rect 1574 -187 1586 -153
rect 1620 -187 1632 -153
rect 1574 -221 1632 -187
rect 1574 -255 1586 -221
rect 1620 -255 1632 -221
rect 1574 -289 1632 -255
rect 1574 -323 1586 -289
rect 1620 -323 1632 -289
rect 1574 -357 1632 -323
rect 1574 -391 1586 -357
rect 1620 -391 1632 -357
rect 1574 -425 1632 -391
rect 1574 -459 1586 -425
rect 1620 -459 1632 -425
rect 1574 -493 1632 -459
rect 1574 -527 1586 -493
rect 1620 -527 1632 -493
rect 1574 -561 1632 -527
rect 1574 -595 1586 -561
rect 1620 -595 1632 -561
rect 1574 -629 1632 -595
rect 1574 -663 1586 -629
rect 1620 -663 1632 -629
rect 1574 -700 1632 -663
<< ndiffc >>
rect -1620 629 -1586 663
rect -1620 561 -1586 595
rect -1620 493 -1586 527
rect -1620 425 -1586 459
rect -1620 357 -1586 391
rect -1620 289 -1586 323
rect -1620 221 -1586 255
rect -1620 153 -1586 187
rect -1620 85 -1586 119
rect -1620 17 -1586 51
rect -1620 -51 -1586 -17
rect -1620 -119 -1586 -85
rect -1620 -187 -1586 -153
rect -1620 -255 -1586 -221
rect -1620 -323 -1586 -289
rect -1620 -391 -1586 -357
rect -1620 -459 -1586 -425
rect -1620 -527 -1586 -493
rect -1620 -595 -1586 -561
rect -1620 -663 -1586 -629
rect -1162 629 -1128 663
rect -1162 561 -1128 595
rect -1162 493 -1128 527
rect -1162 425 -1128 459
rect -1162 357 -1128 391
rect -1162 289 -1128 323
rect -1162 221 -1128 255
rect -1162 153 -1128 187
rect -1162 85 -1128 119
rect -1162 17 -1128 51
rect -1162 -51 -1128 -17
rect -1162 -119 -1128 -85
rect -1162 -187 -1128 -153
rect -1162 -255 -1128 -221
rect -1162 -323 -1128 -289
rect -1162 -391 -1128 -357
rect -1162 -459 -1128 -425
rect -1162 -527 -1128 -493
rect -1162 -595 -1128 -561
rect -1162 -663 -1128 -629
rect -704 629 -670 663
rect -704 561 -670 595
rect -704 493 -670 527
rect -704 425 -670 459
rect -704 357 -670 391
rect -704 289 -670 323
rect -704 221 -670 255
rect -704 153 -670 187
rect -704 85 -670 119
rect -704 17 -670 51
rect -704 -51 -670 -17
rect -704 -119 -670 -85
rect -704 -187 -670 -153
rect -704 -255 -670 -221
rect -704 -323 -670 -289
rect -704 -391 -670 -357
rect -704 -459 -670 -425
rect -704 -527 -670 -493
rect -704 -595 -670 -561
rect -704 -663 -670 -629
rect -246 629 -212 663
rect -246 561 -212 595
rect -246 493 -212 527
rect -246 425 -212 459
rect -246 357 -212 391
rect -246 289 -212 323
rect -246 221 -212 255
rect -246 153 -212 187
rect -246 85 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -85
rect -246 -187 -212 -153
rect -246 -255 -212 -221
rect -246 -323 -212 -289
rect -246 -391 -212 -357
rect -246 -459 -212 -425
rect -246 -527 -212 -493
rect -246 -595 -212 -561
rect -246 -663 -212 -629
rect 212 629 246 663
rect 212 561 246 595
rect 212 493 246 527
rect 212 425 246 459
rect 212 357 246 391
rect 212 289 246 323
rect 212 221 246 255
rect 212 153 246 187
rect 212 85 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -85
rect 212 -187 246 -153
rect 212 -255 246 -221
rect 212 -323 246 -289
rect 212 -391 246 -357
rect 212 -459 246 -425
rect 212 -527 246 -493
rect 212 -595 246 -561
rect 212 -663 246 -629
rect 670 629 704 663
rect 670 561 704 595
rect 670 493 704 527
rect 670 425 704 459
rect 670 357 704 391
rect 670 289 704 323
rect 670 221 704 255
rect 670 153 704 187
rect 670 85 704 119
rect 670 17 704 51
rect 670 -51 704 -17
rect 670 -119 704 -85
rect 670 -187 704 -153
rect 670 -255 704 -221
rect 670 -323 704 -289
rect 670 -391 704 -357
rect 670 -459 704 -425
rect 670 -527 704 -493
rect 670 -595 704 -561
rect 670 -663 704 -629
rect 1128 629 1162 663
rect 1128 561 1162 595
rect 1128 493 1162 527
rect 1128 425 1162 459
rect 1128 357 1162 391
rect 1128 289 1162 323
rect 1128 221 1162 255
rect 1128 153 1162 187
rect 1128 85 1162 119
rect 1128 17 1162 51
rect 1128 -51 1162 -17
rect 1128 -119 1162 -85
rect 1128 -187 1162 -153
rect 1128 -255 1162 -221
rect 1128 -323 1162 -289
rect 1128 -391 1162 -357
rect 1128 -459 1162 -425
rect 1128 -527 1162 -493
rect 1128 -595 1162 -561
rect 1128 -663 1162 -629
rect 1586 629 1620 663
rect 1586 561 1620 595
rect 1586 493 1620 527
rect 1586 425 1620 459
rect 1586 357 1620 391
rect 1586 289 1620 323
rect 1586 221 1620 255
rect 1586 153 1620 187
rect 1586 85 1620 119
rect 1586 17 1620 51
rect 1586 -51 1620 -17
rect 1586 -119 1620 -85
rect 1586 -187 1620 -153
rect 1586 -255 1620 -221
rect 1586 -323 1620 -289
rect 1586 -391 1620 -357
rect 1586 -459 1620 -425
rect 1586 -527 1620 -493
rect 1586 -595 1620 -561
rect 1586 -663 1620 -629
<< psubdiff >>
rect -1734 840 -1615 874
rect -1581 840 -1547 874
rect -1513 840 -1479 874
rect -1445 840 -1411 874
rect -1377 840 -1343 874
rect -1309 840 -1275 874
rect -1241 840 -1207 874
rect -1173 840 -1139 874
rect -1105 840 -1071 874
rect -1037 840 -1003 874
rect -969 840 -935 874
rect -901 840 -867 874
rect -833 840 -799 874
rect -765 840 -731 874
rect -697 840 -663 874
rect -629 840 -595 874
rect -561 840 -527 874
rect -493 840 -459 874
rect -425 840 -391 874
rect -357 840 -323 874
rect -289 840 -255 874
rect -221 840 -187 874
rect -153 840 -119 874
rect -85 840 -51 874
rect -17 840 17 874
rect 51 840 85 874
rect 119 840 153 874
rect 187 840 221 874
rect 255 840 289 874
rect 323 840 357 874
rect 391 840 425 874
rect 459 840 493 874
rect 527 840 561 874
rect 595 840 629 874
rect 663 840 697 874
rect 731 840 765 874
rect 799 840 833 874
rect 867 840 901 874
rect 935 840 969 874
rect 1003 840 1037 874
rect 1071 840 1105 874
rect 1139 840 1173 874
rect 1207 840 1241 874
rect 1275 840 1309 874
rect 1343 840 1377 874
rect 1411 840 1445 874
rect 1479 840 1513 874
rect 1547 840 1581 874
rect 1615 840 1734 874
rect -1734 765 -1700 840
rect -1734 697 -1700 731
rect 1700 765 1734 840
rect -1734 629 -1700 663
rect -1734 561 -1700 595
rect -1734 493 -1700 527
rect -1734 425 -1700 459
rect -1734 357 -1700 391
rect -1734 289 -1700 323
rect -1734 221 -1700 255
rect -1734 153 -1700 187
rect -1734 85 -1700 119
rect -1734 17 -1700 51
rect -1734 -51 -1700 -17
rect -1734 -119 -1700 -85
rect -1734 -187 -1700 -153
rect -1734 -255 -1700 -221
rect -1734 -323 -1700 -289
rect -1734 -391 -1700 -357
rect -1734 -459 -1700 -425
rect -1734 -527 -1700 -493
rect -1734 -595 -1700 -561
rect -1734 -663 -1700 -629
rect -1734 -731 -1700 -697
rect 1700 697 1734 731
rect 1700 629 1734 663
rect 1700 561 1734 595
rect 1700 493 1734 527
rect 1700 425 1734 459
rect 1700 357 1734 391
rect 1700 289 1734 323
rect 1700 221 1734 255
rect 1700 153 1734 187
rect 1700 85 1734 119
rect 1700 17 1734 51
rect 1700 -51 1734 -17
rect 1700 -119 1734 -85
rect 1700 -187 1734 -153
rect 1700 -255 1734 -221
rect 1700 -323 1734 -289
rect 1700 -391 1734 -357
rect 1700 -459 1734 -425
rect 1700 -527 1734 -493
rect 1700 -595 1734 -561
rect 1700 -663 1734 -629
rect -1734 -840 -1700 -765
rect 1700 -731 1734 -697
rect 1700 -840 1734 -765
rect -1734 -874 -1615 -840
rect -1581 -874 -1547 -840
rect -1513 -874 -1479 -840
rect -1445 -874 -1411 -840
rect -1377 -874 -1343 -840
rect -1309 -874 -1275 -840
rect -1241 -874 -1207 -840
rect -1173 -874 -1139 -840
rect -1105 -874 -1071 -840
rect -1037 -874 -1003 -840
rect -969 -874 -935 -840
rect -901 -874 -867 -840
rect -833 -874 -799 -840
rect -765 -874 -731 -840
rect -697 -874 -663 -840
rect -629 -874 -595 -840
rect -561 -874 -527 -840
rect -493 -874 -459 -840
rect -425 -874 -391 -840
rect -357 -874 -323 -840
rect -289 -874 -255 -840
rect -221 -874 -187 -840
rect -153 -874 -119 -840
rect -85 -874 -51 -840
rect -17 -874 17 -840
rect 51 -874 85 -840
rect 119 -874 153 -840
rect 187 -874 221 -840
rect 255 -874 289 -840
rect 323 -874 357 -840
rect 391 -874 425 -840
rect 459 -874 493 -840
rect 527 -874 561 -840
rect 595 -874 629 -840
rect 663 -874 697 -840
rect 731 -874 765 -840
rect 799 -874 833 -840
rect 867 -874 901 -840
rect 935 -874 969 -840
rect 1003 -874 1037 -840
rect 1071 -874 1105 -840
rect 1139 -874 1173 -840
rect 1207 -874 1241 -840
rect 1275 -874 1309 -840
rect 1343 -874 1377 -840
rect 1411 -874 1445 -840
rect 1479 -874 1513 -840
rect 1547 -874 1581 -840
rect 1615 -874 1734 -840
<< psubdiffcont >>
rect -1615 840 -1581 874
rect -1547 840 -1513 874
rect -1479 840 -1445 874
rect -1411 840 -1377 874
rect -1343 840 -1309 874
rect -1275 840 -1241 874
rect -1207 840 -1173 874
rect -1139 840 -1105 874
rect -1071 840 -1037 874
rect -1003 840 -969 874
rect -935 840 -901 874
rect -867 840 -833 874
rect -799 840 -765 874
rect -731 840 -697 874
rect -663 840 -629 874
rect -595 840 -561 874
rect -527 840 -493 874
rect -459 840 -425 874
rect -391 840 -357 874
rect -323 840 -289 874
rect -255 840 -221 874
rect -187 840 -153 874
rect -119 840 -85 874
rect -51 840 -17 874
rect 17 840 51 874
rect 85 840 119 874
rect 153 840 187 874
rect 221 840 255 874
rect 289 840 323 874
rect 357 840 391 874
rect 425 840 459 874
rect 493 840 527 874
rect 561 840 595 874
rect 629 840 663 874
rect 697 840 731 874
rect 765 840 799 874
rect 833 840 867 874
rect 901 840 935 874
rect 969 840 1003 874
rect 1037 840 1071 874
rect 1105 840 1139 874
rect 1173 840 1207 874
rect 1241 840 1275 874
rect 1309 840 1343 874
rect 1377 840 1411 874
rect 1445 840 1479 874
rect 1513 840 1547 874
rect 1581 840 1615 874
rect -1734 731 -1700 765
rect 1700 731 1734 765
rect -1734 663 -1700 697
rect -1734 595 -1700 629
rect -1734 527 -1700 561
rect -1734 459 -1700 493
rect -1734 391 -1700 425
rect -1734 323 -1700 357
rect -1734 255 -1700 289
rect -1734 187 -1700 221
rect -1734 119 -1700 153
rect -1734 51 -1700 85
rect -1734 -17 -1700 17
rect -1734 -85 -1700 -51
rect -1734 -153 -1700 -119
rect -1734 -221 -1700 -187
rect -1734 -289 -1700 -255
rect -1734 -357 -1700 -323
rect -1734 -425 -1700 -391
rect -1734 -493 -1700 -459
rect -1734 -561 -1700 -527
rect -1734 -629 -1700 -595
rect -1734 -697 -1700 -663
rect 1700 663 1734 697
rect 1700 595 1734 629
rect 1700 527 1734 561
rect 1700 459 1734 493
rect 1700 391 1734 425
rect 1700 323 1734 357
rect 1700 255 1734 289
rect 1700 187 1734 221
rect 1700 119 1734 153
rect 1700 51 1734 85
rect 1700 -17 1734 17
rect 1700 -85 1734 -51
rect 1700 -153 1734 -119
rect 1700 -221 1734 -187
rect 1700 -289 1734 -255
rect 1700 -357 1734 -323
rect 1700 -425 1734 -391
rect 1700 -493 1734 -459
rect 1700 -561 1734 -527
rect 1700 -629 1734 -595
rect 1700 -697 1734 -663
rect -1734 -765 -1700 -731
rect 1700 -765 1734 -731
rect -1615 -874 -1581 -840
rect -1547 -874 -1513 -840
rect -1479 -874 -1445 -840
rect -1411 -874 -1377 -840
rect -1343 -874 -1309 -840
rect -1275 -874 -1241 -840
rect -1207 -874 -1173 -840
rect -1139 -874 -1105 -840
rect -1071 -874 -1037 -840
rect -1003 -874 -969 -840
rect -935 -874 -901 -840
rect -867 -874 -833 -840
rect -799 -874 -765 -840
rect -731 -874 -697 -840
rect -663 -874 -629 -840
rect -595 -874 -561 -840
rect -527 -874 -493 -840
rect -459 -874 -425 -840
rect -391 -874 -357 -840
rect -323 -874 -289 -840
rect -255 -874 -221 -840
rect -187 -874 -153 -840
rect -119 -874 -85 -840
rect -51 -874 -17 -840
rect 17 -874 51 -840
rect 85 -874 119 -840
rect 153 -874 187 -840
rect 221 -874 255 -840
rect 289 -874 323 -840
rect 357 -874 391 -840
rect 425 -874 459 -840
rect 493 -874 527 -840
rect 561 -874 595 -840
rect 629 -874 663 -840
rect 697 -874 731 -840
rect 765 -874 799 -840
rect 833 -874 867 -840
rect 901 -874 935 -840
rect 969 -874 1003 -840
rect 1037 -874 1071 -840
rect 1105 -874 1139 -840
rect 1173 -874 1207 -840
rect 1241 -874 1275 -840
rect 1309 -874 1343 -840
rect 1377 -874 1411 -840
rect 1445 -874 1479 -840
rect 1513 -874 1547 -840
rect 1581 -874 1615 -840
<< poly >>
rect -1574 772 -1174 788
rect -1574 738 -1527 772
rect -1493 738 -1459 772
rect -1425 738 -1391 772
rect -1357 738 -1323 772
rect -1289 738 -1255 772
rect -1221 738 -1174 772
rect -1574 700 -1174 738
rect -1116 772 -716 788
rect -1116 738 -1069 772
rect -1035 738 -1001 772
rect -967 738 -933 772
rect -899 738 -865 772
rect -831 738 -797 772
rect -763 738 -716 772
rect -1116 700 -716 738
rect -658 772 -258 788
rect -658 738 -611 772
rect -577 738 -543 772
rect -509 738 -475 772
rect -441 738 -407 772
rect -373 738 -339 772
rect -305 738 -258 772
rect -658 700 -258 738
rect -200 772 200 788
rect -200 738 -153 772
rect -119 738 -85 772
rect -51 738 -17 772
rect 17 738 51 772
rect 85 738 119 772
rect 153 738 200 772
rect -200 700 200 738
rect 258 772 658 788
rect 258 738 305 772
rect 339 738 373 772
rect 407 738 441 772
rect 475 738 509 772
rect 543 738 577 772
rect 611 738 658 772
rect 258 700 658 738
rect 716 772 1116 788
rect 716 738 763 772
rect 797 738 831 772
rect 865 738 899 772
rect 933 738 967 772
rect 1001 738 1035 772
rect 1069 738 1116 772
rect 716 700 1116 738
rect 1174 772 1574 788
rect 1174 738 1221 772
rect 1255 738 1289 772
rect 1323 738 1357 772
rect 1391 738 1425 772
rect 1459 738 1493 772
rect 1527 738 1574 772
rect 1174 700 1574 738
rect -1574 -738 -1174 -700
rect -1574 -772 -1527 -738
rect -1493 -772 -1459 -738
rect -1425 -772 -1391 -738
rect -1357 -772 -1323 -738
rect -1289 -772 -1255 -738
rect -1221 -772 -1174 -738
rect -1574 -788 -1174 -772
rect -1116 -738 -716 -700
rect -1116 -772 -1069 -738
rect -1035 -772 -1001 -738
rect -967 -772 -933 -738
rect -899 -772 -865 -738
rect -831 -772 -797 -738
rect -763 -772 -716 -738
rect -1116 -788 -716 -772
rect -658 -738 -258 -700
rect -658 -772 -611 -738
rect -577 -772 -543 -738
rect -509 -772 -475 -738
rect -441 -772 -407 -738
rect -373 -772 -339 -738
rect -305 -772 -258 -738
rect -658 -788 -258 -772
rect -200 -738 200 -700
rect -200 -772 -153 -738
rect -119 -772 -85 -738
rect -51 -772 -17 -738
rect 17 -772 51 -738
rect 85 -772 119 -738
rect 153 -772 200 -738
rect -200 -788 200 -772
rect 258 -738 658 -700
rect 258 -772 305 -738
rect 339 -772 373 -738
rect 407 -772 441 -738
rect 475 -772 509 -738
rect 543 -772 577 -738
rect 611 -772 658 -738
rect 258 -788 658 -772
rect 716 -738 1116 -700
rect 716 -772 763 -738
rect 797 -772 831 -738
rect 865 -772 899 -738
rect 933 -772 967 -738
rect 1001 -772 1035 -738
rect 1069 -772 1116 -738
rect 716 -788 1116 -772
rect 1174 -738 1574 -700
rect 1174 -772 1221 -738
rect 1255 -772 1289 -738
rect 1323 -772 1357 -738
rect 1391 -772 1425 -738
rect 1459 -772 1493 -738
rect 1527 -772 1574 -738
rect 1174 -788 1574 -772
<< polycont >>
rect -1527 738 -1493 772
rect -1459 738 -1425 772
rect -1391 738 -1357 772
rect -1323 738 -1289 772
rect -1255 738 -1221 772
rect -1069 738 -1035 772
rect -1001 738 -967 772
rect -933 738 -899 772
rect -865 738 -831 772
rect -797 738 -763 772
rect -611 738 -577 772
rect -543 738 -509 772
rect -475 738 -441 772
rect -407 738 -373 772
rect -339 738 -305 772
rect -153 738 -119 772
rect -85 738 -51 772
rect -17 738 17 772
rect 51 738 85 772
rect 119 738 153 772
rect 305 738 339 772
rect 373 738 407 772
rect 441 738 475 772
rect 509 738 543 772
rect 577 738 611 772
rect 763 738 797 772
rect 831 738 865 772
rect 899 738 933 772
rect 967 738 1001 772
rect 1035 738 1069 772
rect 1221 738 1255 772
rect 1289 738 1323 772
rect 1357 738 1391 772
rect 1425 738 1459 772
rect 1493 738 1527 772
rect -1527 -772 -1493 -738
rect -1459 -772 -1425 -738
rect -1391 -772 -1357 -738
rect -1323 -772 -1289 -738
rect -1255 -772 -1221 -738
rect -1069 -772 -1035 -738
rect -1001 -772 -967 -738
rect -933 -772 -899 -738
rect -865 -772 -831 -738
rect -797 -772 -763 -738
rect -611 -772 -577 -738
rect -543 -772 -509 -738
rect -475 -772 -441 -738
rect -407 -772 -373 -738
rect -339 -772 -305 -738
rect -153 -772 -119 -738
rect -85 -772 -51 -738
rect -17 -772 17 -738
rect 51 -772 85 -738
rect 119 -772 153 -738
rect 305 -772 339 -738
rect 373 -772 407 -738
rect 441 -772 475 -738
rect 509 -772 543 -738
rect 577 -772 611 -738
rect 763 -772 797 -738
rect 831 -772 865 -738
rect 899 -772 933 -738
rect 967 -772 1001 -738
rect 1035 -772 1069 -738
rect 1221 -772 1255 -738
rect 1289 -772 1323 -738
rect 1357 -772 1391 -738
rect 1425 -772 1459 -738
rect 1493 -772 1527 -738
<< locali >>
rect -1734 840 -1615 874
rect -1581 840 -1547 874
rect -1513 840 -1479 874
rect -1445 840 -1411 874
rect -1377 840 -1343 874
rect -1309 840 -1275 874
rect -1241 840 -1207 874
rect -1173 840 -1139 874
rect -1105 840 -1071 874
rect -1037 840 -1003 874
rect -969 840 -935 874
rect -901 840 -867 874
rect -833 840 -799 874
rect -765 840 -731 874
rect -697 840 -663 874
rect -629 840 -595 874
rect -561 840 -527 874
rect -493 840 -459 874
rect -425 840 -391 874
rect -357 840 -323 874
rect -289 840 -255 874
rect -221 840 -187 874
rect -153 840 -119 874
rect -85 840 -51 874
rect -17 840 17 874
rect 51 840 85 874
rect 119 840 153 874
rect 187 840 221 874
rect 255 840 289 874
rect 323 840 357 874
rect 391 840 425 874
rect 459 840 493 874
rect 527 840 561 874
rect 595 840 629 874
rect 663 840 697 874
rect 731 840 765 874
rect 799 840 833 874
rect 867 840 901 874
rect 935 840 969 874
rect 1003 840 1037 874
rect 1071 840 1105 874
rect 1139 840 1173 874
rect 1207 840 1241 874
rect 1275 840 1309 874
rect 1343 840 1377 874
rect 1411 840 1445 874
rect 1479 840 1513 874
rect 1547 840 1581 874
rect 1615 840 1734 874
rect -1734 765 -1700 840
rect -1574 738 -1527 772
rect -1493 738 -1459 772
rect -1425 738 -1391 772
rect -1357 738 -1323 772
rect -1289 738 -1255 772
rect -1221 738 -1174 772
rect -1116 738 -1069 772
rect -1035 738 -1001 772
rect -967 738 -933 772
rect -899 738 -865 772
rect -831 738 -797 772
rect -763 738 -716 772
rect -658 738 -611 772
rect -577 738 -543 772
rect -509 738 -475 772
rect -441 738 -407 772
rect -373 738 -339 772
rect -305 738 -258 772
rect -200 738 -153 772
rect -119 738 -85 772
rect -51 738 -17 772
rect 17 738 51 772
rect 85 738 119 772
rect 153 738 200 772
rect 258 738 305 772
rect 339 738 373 772
rect 407 738 441 772
rect 475 738 509 772
rect 543 738 577 772
rect 611 738 658 772
rect 716 738 763 772
rect 797 738 831 772
rect 865 738 899 772
rect 933 738 967 772
rect 1001 738 1035 772
rect 1069 738 1116 772
rect 1174 738 1221 772
rect 1255 738 1289 772
rect 1323 738 1357 772
rect 1391 738 1425 772
rect 1459 738 1493 772
rect 1527 738 1574 772
rect 1700 765 1734 840
rect -1734 697 -1700 731
rect -1734 629 -1700 663
rect -1734 561 -1700 595
rect -1734 493 -1700 527
rect -1734 425 -1700 459
rect -1734 357 -1700 391
rect -1734 289 -1700 323
rect -1734 221 -1700 255
rect -1734 153 -1700 187
rect -1734 85 -1700 119
rect -1734 17 -1700 51
rect -1734 -51 -1700 -17
rect -1734 -119 -1700 -85
rect -1734 -187 -1700 -153
rect -1734 -255 -1700 -221
rect -1734 -323 -1700 -289
rect -1734 -391 -1700 -357
rect -1734 -459 -1700 -425
rect -1734 -527 -1700 -493
rect -1734 -595 -1700 -561
rect -1734 -663 -1700 -629
rect -1734 -731 -1700 -697
rect -1620 663 -1586 704
rect -1620 595 -1586 629
rect -1620 527 -1586 561
rect -1620 459 -1586 493
rect -1620 391 -1586 425
rect -1620 323 -1586 357
rect -1620 255 -1586 289
rect -1620 187 -1586 221
rect -1620 119 -1586 153
rect -1620 51 -1586 85
rect -1620 -17 -1586 17
rect -1620 -85 -1586 -51
rect -1620 -153 -1586 -119
rect -1620 -221 -1586 -187
rect -1620 -289 -1586 -255
rect -1620 -357 -1586 -323
rect -1620 -425 -1586 -391
rect -1620 -493 -1586 -459
rect -1620 -561 -1586 -527
rect -1620 -629 -1586 -595
rect -1620 -704 -1586 -663
rect -1162 663 -1128 704
rect -1162 595 -1128 629
rect -1162 527 -1128 561
rect -1162 459 -1128 493
rect -1162 391 -1128 425
rect -1162 323 -1128 357
rect -1162 255 -1128 289
rect -1162 187 -1128 221
rect -1162 119 -1128 153
rect -1162 51 -1128 85
rect -1162 -17 -1128 17
rect -1162 -85 -1128 -51
rect -1162 -153 -1128 -119
rect -1162 -221 -1128 -187
rect -1162 -289 -1128 -255
rect -1162 -357 -1128 -323
rect -1162 -425 -1128 -391
rect -1162 -493 -1128 -459
rect -1162 -561 -1128 -527
rect -1162 -629 -1128 -595
rect -1162 -704 -1128 -663
rect -704 663 -670 704
rect -704 595 -670 629
rect -704 527 -670 561
rect -704 459 -670 493
rect -704 391 -670 425
rect -704 323 -670 357
rect -704 255 -670 289
rect -704 187 -670 221
rect -704 119 -670 153
rect -704 51 -670 85
rect -704 -17 -670 17
rect -704 -85 -670 -51
rect -704 -153 -670 -119
rect -704 -221 -670 -187
rect -704 -289 -670 -255
rect -704 -357 -670 -323
rect -704 -425 -670 -391
rect -704 -493 -670 -459
rect -704 -561 -670 -527
rect -704 -629 -670 -595
rect -704 -704 -670 -663
rect -246 663 -212 704
rect -246 595 -212 629
rect -246 527 -212 561
rect -246 459 -212 493
rect -246 391 -212 425
rect -246 323 -212 357
rect -246 255 -212 289
rect -246 187 -212 221
rect -246 119 -212 153
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect -246 -153 -212 -119
rect -246 -221 -212 -187
rect -246 -289 -212 -255
rect -246 -357 -212 -323
rect -246 -425 -212 -391
rect -246 -493 -212 -459
rect -246 -561 -212 -527
rect -246 -629 -212 -595
rect -246 -704 -212 -663
rect 212 663 246 704
rect 212 595 246 629
rect 212 527 246 561
rect 212 459 246 493
rect 212 391 246 425
rect 212 323 246 357
rect 212 255 246 289
rect 212 187 246 221
rect 212 119 246 153
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
rect 212 -153 246 -119
rect 212 -221 246 -187
rect 212 -289 246 -255
rect 212 -357 246 -323
rect 212 -425 246 -391
rect 212 -493 246 -459
rect 212 -561 246 -527
rect 212 -629 246 -595
rect 212 -704 246 -663
rect 670 663 704 704
rect 670 595 704 629
rect 670 527 704 561
rect 670 459 704 493
rect 670 391 704 425
rect 670 323 704 357
rect 670 255 704 289
rect 670 187 704 221
rect 670 119 704 153
rect 670 51 704 85
rect 670 -17 704 17
rect 670 -85 704 -51
rect 670 -153 704 -119
rect 670 -221 704 -187
rect 670 -289 704 -255
rect 670 -357 704 -323
rect 670 -425 704 -391
rect 670 -493 704 -459
rect 670 -561 704 -527
rect 670 -629 704 -595
rect 670 -704 704 -663
rect 1128 663 1162 704
rect 1128 595 1162 629
rect 1128 527 1162 561
rect 1128 459 1162 493
rect 1128 391 1162 425
rect 1128 323 1162 357
rect 1128 255 1162 289
rect 1128 187 1162 221
rect 1128 119 1162 153
rect 1128 51 1162 85
rect 1128 -17 1162 17
rect 1128 -85 1162 -51
rect 1128 -153 1162 -119
rect 1128 -221 1162 -187
rect 1128 -289 1162 -255
rect 1128 -357 1162 -323
rect 1128 -425 1162 -391
rect 1128 -493 1162 -459
rect 1128 -561 1162 -527
rect 1128 -629 1162 -595
rect 1128 -704 1162 -663
rect 1586 663 1620 704
rect 1586 595 1620 629
rect 1586 527 1620 561
rect 1586 459 1620 493
rect 1586 391 1620 425
rect 1586 323 1620 357
rect 1586 255 1620 289
rect 1586 187 1620 221
rect 1586 119 1620 153
rect 1586 51 1620 85
rect 1586 -17 1620 17
rect 1586 -85 1620 -51
rect 1586 -153 1620 -119
rect 1586 -221 1620 -187
rect 1586 -289 1620 -255
rect 1586 -357 1620 -323
rect 1586 -425 1620 -391
rect 1586 -493 1620 -459
rect 1586 -561 1620 -527
rect 1586 -629 1620 -595
rect 1586 -704 1620 -663
rect 1700 697 1734 731
rect 1700 629 1734 663
rect 1700 561 1734 595
rect 1700 493 1734 527
rect 1700 425 1734 459
rect 1700 357 1734 391
rect 1700 289 1734 323
rect 1700 221 1734 255
rect 1700 153 1734 187
rect 1700 85 1734 119
rect 1700 17 1734 51
rect 1700 -51 1734 -17
rect 1700 -119 1734 -85
rect 1700 -187 1734 -153
rect 1700 -255 1734 -221
rect 1700 -323 1734 -289
rect 1700 -391 1734 -357
rect 1700 -459 1734 -425
rect 1700 -527 1734 -493
rect 1700 -595 1734 -561
rect 1700 -663 1734 -629
rect 1700 -731 1734 -697
rect -1734 -840 -1700 -765
rect -1574 -772 -1527 -738
rect -1493 -772 -1459 -738
rect -1425 -772 -1391 -738
rect -1357 -772 -1323 -738
rect -1289 -772 -1255 -738
rect -1221 -772 -1174 -738
rect -1116 -772 -1069 -738
rect -1035 -772 -1001 -738
rect -967 -772 -933 -738
rect -899 -772 -865 -738
rect -831 -772 -797 -738
rect -763 -772 -716 -738
rect -658 -772 -611 -738
rect -577 -772 -543 -738
rect -509 -772 -475 -738
rect -441 -772 -407 -738
rect -373 -772 -339 -738
rect -305 -772 -258 -738
rect -200 -772 -153 -738
rect -119 -772 -85 -738
rect -51 -772 -17 -738
rect 17 -772 51 -738
rect 85 -772 119 -738
rect 153 -772 200 -738
rect 258 -772 305 -738
rect 339 -772 373 -738
rect 407 -772 441 -738
rect 475 -772 509 -738
rect 543 -772 577 -738
rect 611 -772 658 -738
rect 716 -772 763 -738
rect 797 -772 831 -738
rect 865 -772 899 -738
rect 933 -772 967 -738
rect 1001 -772 1035 -738
rect 1069 -772 1116 -738
rect 1174 -772 1221 -738
rect 1255 -772 1289 -738
rect 1323 -772 1357 -738
rect 1391 -772 1425 -738
rect 1459 -772 1493 -738
rect 1527 -772 1574 -738
rect 1700 -840 1734 -765
rect -1734 -874 -1615 -840
rect -1581 -874 -1547 -840
rect -1513 -874 -1479 -840
rect -1445 -874 -1411 -840
rect -1377 -874 -1343 -840
rect -1309 -874 -1275 -840
rect -1241 -874 -1207 -840
rect -1173 -874 -1139 -840
rect -1105 -874 -1071 -840
rect -1037 -874 -1003 -840
rect -969 -874 -935 -840
rect -901 -874 -867 -840
rect -833 -874 -799 -840
rect -765 -874 -731 -840
rect -697 -874 -663 -840
rect -629 -874 -595 -840
rect -561 -874 -527 -840
rect -493 -874 -459 -840
rect -425 -874 -391 -840
rect -357 -874 -323 -840
rect -289 -874 -255 -840
rect -221 -874 -187 -840
rect -153 -874 -119 -840
rect -85 -874 -51 -840
rect -17 -874 17 -840
rect 51 -874 85 -840
rect 119 -874 153 -840
rect 187 -874 221 -840
rect 255 -874 289 -840
rect 323 -874 357 -840
rect 391 -874 425 -840
rect 459 -874 493 -840
rect 527 -874 561 -840
rect 595 -874 629 -840
rect 663 -874 697 -840
rect 731 -874 765 -840
rect 799 -874 833 -840
rect 867 -874 901 -840
rect 935 -874 969 -840
rect 1003 -874 1037 -840
rect 1071 -874 1105 -840
rect 1139 -874 1173 -840
rect 1207 -874 1241 -840
rect 1275 -874 1309 -840
rect 1343 -874 1377 -840
rect 1411 -874 1445 -840
rect 1479 -874 1513 -840
rect 1547 -874 1581 -840
rect 1615 -874 1734 -840
<< properties >>
string FIXED_BBOX -1716 -856 1716 856
<< end >>
