magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -611 190 611 224
rect -611 -190 -577 190
rect 577 -190 611 190
rect -611 -224 611 -190
<< nmoslvt >>
rect -447 -50 -417 50
rect -351 -50 -321 50
rect -255 -50 -225 50
rect -159 -50 -129 50
rect -63 -50 -33 50
rect 33 -50 63 50
rect 129 -50 159 50
rect 225 -50 255 50
rect 321 -50 351 50
rect 417 -50 447 50
<< ndiff >>
rect -509 17 -447 50
rect -509 -17 -497 17
rect -463 -17 -447 17
rect -509 -50 -447 -17
rect -417 17 -351 50
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -50 -351 -17
rect -321 17 -255 50
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -50 -255 -17
rect -225 17 -159 50
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -50 -159 -17
rect -129 17 -63 50
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -50 -63 -17
rect -33 17 33 50
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -50 33 -17
rect 63 17 129 50
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -50 129 -17
rect 159 17 225 50
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -50 225 -17
rect 255 17 321 50
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -50 321 -17
rect 351 17 417 50
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -50 417 -17
rect 447 17 509 50
rect 447 -17 463 17
rect 497 -17 509 17
rect 447 -50 509 -17
<< ndiffc >>
rect -497 -17 -463 17
rect -401 -17 -367 17
rect -305 -17 -271 17
rect -209 -17 -175 17
rect -113 -17 -79 17
rect -17 -17 17 17
rect 79 -17 113 17
rect 175 -17 209 17
rect 271 -17 305 17
rect 367 -17 401 17
rect 463 -17 497 17
<< psubdiff >>
rect -611 190 -493 224
rect -459 190 -425 224
rect -391 190 -357 224
rect -323 190 -289 224
rect -255 190 -221 224
rect -187 190 -153 224
rect -119 190 -85 224
rect -51 190 -17 224
rect 17 190 51 224
rect 85 190 119 224
rect 153 190 187 224
rect 221 190 255 224
rect 289 190 323 224
rect 357 190 391 224
rect 425 190 459 224
rect 493 190 611 224
rect -611 119 -577 190
rect -611 51 -577 85
rect 577 119 611 190
rect 577 51 611 85
rect -611 -17 -577 17
rect 577 -17 611 17
rect -611 -85 -577 -51
rect -611 -190 -577 -119
rect 577 -85 611 -51
rect 577 -190 611 -119
rect -611 -224 -493 -190
rect -459 -224 -425 -190
rect -391 -224 -357 -190
rect -323 -224 -289 -190
rect -255 -224 -221 -190
rect -187 -224 -153 -190
rect -119 -224 -85 -190
rect -51 -224 -17 -190
rect 17 -224 51 -190
rect 85 -224 119 -190
rect 153 -224 187 -190
rect 221 -224 255 -190
rect 289 -224 323 -190
rect 357 -224 391 -190
rect 425 -224 459 -190
rect 493 -224 611 -190
<< psubdiffcont >>
rect -493 190 -459 224
rect -425 190 -391 224
rect -357 190 -323 224
rect -289 190 -255 224
rect -221 190 -187 224
rect -153 190 -119 224
rect -85 190 -51 224
rect -17 190 17 224
rect 51 190 85 224
rect 119 190 153 224
rect 187 190 221 224
rect 255 190 289 224
rect 323 190 357 224
rect 391 190 425 224
rect 459 190 493 224
rect -611 85 -577 119
rect -611 17 -577 51
rect 577 85 611 119
rect -611 -51 -577 -17
rect 577 17 611 51
rect -611 -119 -577 -85
rect 577 -51 611 -17
rect 577 -119 611 -85
rect -493 -224 -459 -190
rect -425 -224 -391 -190
rect -357 -224 -323 -190
rect -289 -224 -255 -190
rect -221 -224 -187 -190
rect -153 -224 -119 -190
rect -85 -224 -51 -190
rect -17 -224 17 -190
rect 51 -224 85 -190
rect 119 -224 153 -190
rect 187 -224 221 -190
rect 255 -224 289 -190
rect 323 -224 357 -190
rect 391 -224 425 -190
rect 459 -224 493 -190
<< poly >>
rect -369 122 -303 138
rect -369 88 -353 122
rect -319 88 -303 122
rect -447 50 -417 76
rect -369 72 -303 88
rect -177 122 -111 138
rect -177 88 -161 122
rect -127 88 -111 122
rect -351 50 -321 72
rect -255 50 -225 76
rect -177 72 -111 88
rect 15 122 81 138
rect 15 88 31 122
rect 65 88 81 122
rect -159 50 -129 72
rect -63 50 -33 76
rect 15 72 81 88
rect 207 122 273 138
rect 207 88 223 122
rect 257 88 273 122
rect 33 50 63 72
rect 129 50 159 76
rect 207 72 273 88
rect 399 122 465 138
rect 399 88 415 122
rect 449 88 465 122
rect 225 50 255 72
rect 321 50 351 76
rect 399 72 465 88
rect 417 50 447 72
rect -447 -72 -417 -50
rect -465 -88 -399 -72
rect -351 -76 -321 -50
rect -255 -72 -225 -50
rect -465 -122 -449 -88
rect -415 -122 -399 -88
rect -465 -138 -399 -122
rect -273 -88 -207 -72
rect -159 -76 -129 -50
rect -63 -72 -33 -50
rect -273 -122 -257 -88
rect -223 -122 -207 -88
rect -273 -138 -207 -122
rect -81 -88 -15 -72
rect 33 -76 63 -50
rect 129 -72 159 -50
rect -81 -122 -65 -88
rect -31 -122 -15 -88
rect -81 -138 -15 -122
rect 111 -88 177 -72
rect 225 -76 255 -50
rect 321 -72 351 -50
rect 111 -122 127 -88
rect 161 -122 177 -88
rect 111 -138 177 -122
rect 303 -88 369 -72
rect 417 -76 447 -50
rect 303 -122 319 -88
rect 353 -122 369 -88
rect 303 -138 369 -122
<< polycont >>
rect -353 88 -319 122
rect -161 88 -127 122
rect 31 88 65 122
rect 223 88 257 122
rect 415 88 449 122
rect -449 -122 -415 -88
rect -257 -122 -223 -88
rect -65 -122 -31 -88
rect 127 -122 161 -88
rect 319 -122 353 -88
<< locali >>
rect -611 190 -493 224
rect -459 190 -425 224
rect -391 190 -357 224
rect -323 190 -289 224
rect -255 190 -221 224
rect -187 190 -153 224
rect -119 190 -85 224
rect -51 190 -17 224
rect 17 190 51 224
rect 85 190 119 224
rect 153 190 187 224
rect 221 190 255 224
rect 289 190 323 224
rect 357 190 391 224
rect 425 190 459 224
rect 493 190 611 224
rect -611 119 -577 190
rect -369 88 -353 122
rect -319 88 -303 122
rect -177 88 -161 122
rect -127 88 -111 122
rect 15 88 31 122
rect 65 88 81 122
rect 207 88 223 122
rect 257 88 273 122
rect 399 88 415 122
rect 449 88 465 122
rect 577 119 611 190
rect -611 51 -577 85
rect -611 -17 -577 17
rect -611 -85 -577 -51
rect -497 17 -463 54
rect -497 -54 -463 -17
rect -401 17 -367 54
rect -401 -54 -367 -17
rect -305 17 -271 54
rect -305 -54 -271 -17
rect -209 17 -175 54
rect -209 -54 -175 -17
rect -113 17 -79 54
rect -113 -54 -79 -17
rect -17 17 17 54
rect -17 -54 17 -17
rect 79 17 113 54
rect 79 -54 113 -17
rect 175 17 209 54
rect 175 -54 209 -17
rect 271 17 305 54
rect 271 -54 305 -17
rect 367 17 401 54
rect 367 -54 401 -17
rect 463 17 497 54
rect 463 -54 497 -17
rect 577 51 611 85
rect 577 -17 611 17
rect 577 -85 611 -51
rect -611 -190 -577 -119
rect -465 -122 -449 -88
rect -415 -122 -399 -88
rect -273 -122 -257 -88
rect -223 -122 -207 -88
rect -81 -122 -65 -88
rect -31 -122 -15 -88
rect 111 -122 127 -88
rect 161 -122 177 -88
rect 303 -122 319 -88
rect 353 -122 369 -88
rect 577 -190 611 -119
rect -611 -224 -493 -190
rect -459 -224 -425 -190
rect -391 -224 -357 -190
rect -323 -224 -289 -190
rect -255 -224 -221 -190
rect -187 -224 -153 -190
rect -119 -224 -85 -190
rect -51 -224 -17 -190
rect 17 -224 51 -190
rect 85 -224 119 -190
rect 153 -224 187 -190
rect 221 -224 255 -190
rect 289 -224 323 -190
rect 357 -224 391 -190
rect 425 -224 459 -190
rect 493 -224 611 -190
<< viali >>
rect -497 -17 -463 17
rect -401 -17 -367 17
rect -305 -17 -271 17
rect -209 -17 -175 17
rect -113 -17 -79 17
rect -17 -17 17 17
rect 79 -17 113 17
rect 175 -17 209 17
rect 271 -17 305 17
rect 367 -17 401 17
rect 463 -17 497 17
<< metal1 >>
rect -503 17 -457 50
rect -503 -17 -497 17
rect -463 -17 -457 17
rect -503 -50 -457 -17
rect -407 17 -361 50
rect -407 -17 -401 17
rect -367 -17 -361 17
rect -407 -50 -361 -17
rect -311 17 -265 50
rect -311 -17 -305 17
rect -271 -17 -265 17
rect -311 -50 -265 -17
rect -215 17 -169 50
rect -215 -17 -209 17
rect -175 -17 -169 17
rect -215 -50 -169 -17
rect -119 17 -73 50
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -50 -73 -17
rect -23 17 23 50
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -50 23 -17
rect 73 17 119 50
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -50 119 -17
rect 169 17 215 50
rect 169 -17 175 17
rect 209 -17 215 17
rect 169 -50 215 -17
rect 265 17 311 50
rect 265 -17 271 17
rect 305 -17 311 17
rect 265 -50 311 -17
rect 361 17 407 50
rect 361 -17 367 17
rect 401 -17 407 17
rect 361 -50 407 -17
rect 457 17 503 50
rect 457 -17 463 17
rect 497 -17 503 17
rect 457 -50 503 -17
<< properties >>
string FIXED_BBOX -594 -207 594 207
<< end >>
