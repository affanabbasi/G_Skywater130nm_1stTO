magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< locali >>
rect 165785 -25054 166173 -24622
rect 166421 -25054 166809 -24622
rect 167057 -25054 167445 -24622
rect 167693 -25054 168081 -24622
rect 168329 -25054 168717 -24622
rect 160358 -26118 160381 -26084
rect 160415 -26118 160453 -26084
rect 160487 -26118 160525 -26084
rect 160559 -26118 160597 -26084
rect 160631 -26118 160669 -26084
rect 160703 -26118 160741 -26084
rect 160775 -26118 160813 -26084
rect 160847 -26118 160885 -26084
rect 160919 -26118 160957 -26084
rect 160991 -26118 161029 -26084
rect 161063 -26118 161101 -26084
rect 161135 -26118 161173 -26084
rect 161207 -26118 161245 -26084
rect 161279 -26118 161317 -26084
rect 161351 -26118 161389 -26084
rect 161423 -26118 161461 -26084
rect 161495 -26118 161533 -26084
rect 161567 -26118 161605 -26084
rect 161639 -26118 161677 -26084
rect 161711 -26118 161749 -26084
rect 161783 -26118 161821 -26084
rect 161855 -26118 161893 -26084
rect 161927 -26118 161965 -26084
rect 161999 -26118 162037 -26084
rect 162071 -26118 162109 -26084
rect 162143 -26118 162181 -26084
rect 162215 -26118 162253 -26084
rect 162287 -26118 162325 -26084
rect 162359 -26118 162397 -26084
rect 162431 -26118 162469 -26084
rect 162503 -26118 162541 -26084
rect 162575 -26118 162613 -26084
rect 162647 -26118 162685 -26084
rect 162719 -26118 162757 -26084
rect 162791 -26118 162829 -26084
rect 162863 -26118 162901 -26084
rect 162935 -26118 162973 -26084
rect 163007 -26118 163045 -26084
rect 163079 -26118 163117 -26084
rect 163151 -26118 163189 -26084
rect 163223 -26118 163261 -26084
rect 163295 -26118 163333 -26084
rect 163367 -26118 163405 -26084
rect 163439 -26118 163477 -26084
rect 163511 -26118 163549 -26084
rect 163583 -26118 163621 -26084
rect 163655 -26118 163693 -26084
rect 163727 -26118 163765 -26084
rect 163799 -26118 163837 -26084
rect 163871 -26118 163909 -26084
rect 163943 -26118 163981 -26084
rect 164015 -26118 164053 -26084
rect 164087 -26118 164125 -26084
rect 164159 -26118 164197 -26084
rect 164231 -26118 164269 -26084
rect 164303 -26118 164326 -26084
rect 160358 -26528 160381 -26494
rect 160415 -26528 160453 -26494
rect 160487 -26528 160525 -26494
rect 160559 -26528 160597 -26494
rect 160631 -26528 160669 -26494
rect 160703 -26528 160741 -26494
rect 160775 -26528 160813 -26494
rect 160847 -26528 160885 -26494
rect 160919 -26528 160957 -26494
rect 160991 -26528 161029 -26494
rect 161063 -26528 161101 -26494
rect 161135 -26528 161173 -26494
rect 161207 -26528 161245 -26494
rect 161279 -26528 161317 -26494
rect 161351 -26528 161389 -26494
rect 161423 -26528 161461 -26494
rect 161495 -26528 161533 -26494
rect 161567 -26528 161605 -26494
rect 161639 -26528 161677 -26494
rect 161711 -26528 161749 -26494
rect 161783 -26528 161821 -26494
rect 161855 -26528 161893 -26494
rect 161927 -26528 161965 -26494
rect 161999 -26528 162037 -26494
rect 162071 -26528 162109 -26494
rect 162143 -26528 162181 -26494
rect 162215 -26528 162253 -26494
rect 162287 -26528 162325 -26494
rect 162359 -26528 162397 -26494
rect 162431 -26528 162469 -26494
rect 162503 -26528 162541 -26494
rect 162575 -26528 162613 -26494
rect 162647 -26528 162685 -26494
rect 162719 -26528 162757 -26494
rect 162791 -26528 162829 -26494
rect 162863 -26528 162901 -26494
rect 162935 -26528 162973 -26494
rect 163007 -26528 163045 -26494
rect 163079 -26528 163117 -26494
rect 163151 -26528 163189 -26494
rect 163223 -26528 163261 -26494
rect 163295 -26528 163333 -26494
rect 163367 -26528 163405 -26494
rect 163439 -26528 163477 -26494
rect 163511 -26528 163549 -26494
rect 163583 -26528 163621 -26494
rect 163655 -26528 163693 -26494
rect 163727 -26528 163765 -26494
rect 163799 -26528 163837 -26494
rect 163871 -26528 163909 -26494
rect 163943 -26528 163981 -26494
rect 164015 -26528 164053 -26494
rect 164087 -26528 164125 -26494
rect 164159 -26528 164197 -26494
rect 164231 -26528 164269 -26494
rect 164303 -26528 164326 -26494
rect 164438 -26674 165689 -25938
rect 165785 -27073 165855 -27054
rect 165785 -27107 165803 -27073
rect 165837 -27107 165855 -27073
rect 165785 -27145 165855 -27107
rect 165785 -27179 165803 -27145
rect 165837 -27179 165855 -27145
rect 165785 -27217 165855 -27179
rect 165785 -27251 165803 -27217
rect 165837 -27251 165855 -27217
rect 146718 -27412 156544 -27258
rect 165785 -27289 165855 -27251
rect 165785 -27323 165803 -27289
rect 165837 -27323 165855 -27289
rect 165785 -27361 165855 -27323
rect 165785 -27395 165803 -27361
rect 165837 -27395 165855 -27361
rect 146718 -28390 156580 -27412
rect 165785 -27433 165855 -27395
rect 165785 -27467 165803 -27433
rect 165837 -27467 165855 -27433
rect 165785 -27486 165855 -27467
rect 166103 -27486 166491 -27054
rect 166739 -27486 167127 -27054
rect 167375 -27486 167763 -27054
rect 168011 -27486 168399 -27054
rect 168647 -27073 168717 -27054
rect 168647 -27107 168665 -27073
rect 168699 -27107 168717 -27073
rect 168647 -27145 168717 -27107
rect 168647 -27179 168665 -27145
rect 168699 -27179 168717 -27145
rect 168647 -27217 168717 -27179
rect 168647 -27251 168665 -27217
rect 168699 -27251 168717 -27217
rect 168647 -27289 168717 -27251
rect 168647 -27323 168665 -27289
rect 168699 -27323 168717 -27289
rect 168647 -27361 168717 -27323
rect 168647 -27395 168665 -27361
rect 168699 -27395 168717 -27361
rect 168647 -27433 168717 -27395
rect 168647 -27467 168665 -27433
rect 168699 -27467 168717 -27433
rect 168647 -27486 168717 -27467
rect 165655 -28392 166532 -27614
rect 146820 -30688 156480 -30684
rect 146820 -30698 146845 -30688
rect 146718 -30722 146845 -30698
rect 146879 -30722 146917 -30688
rect 146951 -30722 146989 -30688
rect 147023 -30722 147061 -30688
rect 147095 -30722 147133 -30688
rect 147167 -30722 147205 -30688
rect 147239 -30722 147277 -30688
rect 147311 -30722 147349 -30688
rect 147383 -30722 147421 -30688
rect 147455 -30722 147493 -30688
rect 147527 -30722 147565 -30688
rect 147599 -30722 147637 -30688
rect 147671 -30722 147709 -30688
rect 147743 -30722 147781 -30688
rect 147815 -30722 147853 -30688
rect 147887 -30722 147925 -30688
rect 147959 -30722 147997 -30688
rect 148031 -30722 148069 -30688
rect 148103 -30722 148141 -30688
rect 148175 -30722 148213 -30688
rect 148247 -30722 148285 -30688
rect 148319 -30722 148357 -30688
rect 148391 -30722 148429 -30688
rect 148463 -30722 148501 -30688
rect 148535 -30722 148573 -30688
rect 148607 -30722 148645 -30688
rect 148679 -30722 148717 -30688
rect 148751 -30722 148789 -30688
rect 148823 -30722 148861 -30688
rect 148895 -30722 148933 -30688
rect 148967 -30722 149005 -30688
rect 149039 -30722 149077 -30688
rect 149111 -30722 149149 -30688
rect 149183 -30722 149221 -30688
rect 149255 -30722 149293 -30688
rect 149327 -30722 149365 -30688
rect 149399 -30722 149437 -30688
rect 149471 -30722 149509 -30688
rect 149543 -30722 149581 -30688
rect 149615 -30722 149653 -30688
rect 149687 -30722 149725 -30688
rect 149759 -30722 149797 -30688
rect 149831 -30722 149869 -30688
rect 149903 -30722 149941 -30688
rect 149975 -30722 150013 -30688
rect 150047 -30722 150085 -30688
rect 150119 -30722 150157 -30688
rect 150191 -30722 150229 -30688
rect 150263 -30722 150301 -30688
rect 150335 -30722 150373 -30688
rect 150407 -30722 150445 -30688
rect 150479 -30722 150517 -30688
rect 150551 -30722 150589 -30688
rect 150623 -30722 150661 -30688
rect 150695 -30722 150733 -30688
rect 150767 -30722 150805 -30688
rect 150839 -30722 150877 -30688
rect 150911 -30722 150949 -30688
rect 150983 -30722 151021 -30688
rect 151055 -30722 151093 -30688
rect 151127 -30722 151165 -30688
rect 151199 -30722 151237 -30688
rect 151271 -30722 151309 -30688
rect 151343 -30722 151381 -30688
rect 151415 -30722 151453 -30688
rect 151487 -30722 151525 -30688
rect 151559 -30722 151597 -30688
rect 151631 -30722 151669 -30688
rect 151703 -30722 151741 -30688
rect 151775 -30722 151813 -30688
rect 151847 -30722 151885 -30688
rect 151919 -30722 151957 -30688
rect 151991 -30722 152029 -30688
rect 152063 -30722 152101 -30688
rect 152135 -30722 152173 -30688
rect 152207 -30722 152245 -30688
rect 152279 -30722 152317 -30688
rect 152351 -30722 152389 -30688
rect 152423 -30722 152461 -30688
rect 152495 -30722 152533 -30688
rect 152567 -30722 152605 -30688
rect 152639 -30722 152677 -30688
rect 152711 -30722 152749 -30688
rect 152783 -30722 152821 -30688
rect 152855 -30722 152893 -30688
rect 152927 -30722 152965 -30688
rect 152999 -30722 153037 -30688
rect 153071 -30722 153109 -30688
rect 153143 -30722 153181 -30688
rect 153215 -30722 153253 -30688
rect 153287 -30722 153325 -30688
rect 153359 -30722 153397 -30688
rect 153431 -30722 153469 -30688
rect 153503 -30722 153541 -30688
rect 153575 -30722 153613 -30688
rect 153647 -30722 153685 -30688
rect 153719 -30722 153757 -30688
rect 153791 -30722 153829 -30688
rect 153863 -30722 153901 -30688
rect 153935 -30722 153973 -30688
rect 154007 -30722 154045 -30688
rect 154079 -30722 154117 -30688
rect 154151 -30722 154189 -30688
rect 154223 -30722 154261 -30688
rect 154295 -30722 154333 -30688
rect 154367 -30722 154405 -30688
rect 154439 -30722 154477 -30688
rect 154511 -30722 154549 -30688
rect 154583 -30722 154621 -30688
rect 154655 -30722 154693 -30688
rect 154727 -30722 154765 -30688
rect 154799 -30722 154837 -30688
rect 154871 -30722 154909 -30688
rect 154943 -30722 154981 -30688
rect 155015 -30722 155053 -30688
rect 155087 -30722 155125 -30688
rect 155159 -30722 155197 -30688
rect 155231 -30722 155269 -30688
rect 155303 -30722 155341 -30688
rect 155375 -30722 155413 -30688
rect 155447 -30722 155485 -30688
rect 155519 -30722 155557 -30688
rect 155591 -30722 155629 -30688
rect 155663 -30722 155701 -30688
rect 155735 -30722 155773 -30688
rect 155807 -30722 155845 -30688
rect 155879 -30722 155917 -30688
rect 155951 -30722 155989 -30688
rect 156023 -30722 156061 -30688
rect 156095 -30722 156133 -30688
rect 156167 -30722 156205 -30688
rect 156239 -30722 156277 -30688
rect 156311 -30722 156349 -30688
rect 156383 -30722 156421 -30688
rect 156455 -30698 156480 -30688
rect 157854 -30688 167514 -30684
rect 156455 -30722 156580 -30698
rect 146718 -30732 156580 -30722
rect 157854 -30722 157879 -30688
rect 157913 -30722 157951 -30688
rect 157985 -30722 158023 -30688
rect 158057 -30722 158095 -30688
rect 158129 -30722 158167 -30688
rect 158201 -30722 158239 -30688
rect 158273 -30722 158311 -30688
rect 158345 -30722 158383 -30688
rect 158417 -30722 158455 -30688
rect 158489 -30722 158527 -30688
rect 158561 -30722 158599 -30688
rect 158633 -30722 158671 -30688
rect 158705 -30722 158743 -30688
rect 158777 -30722 158815 -30688
rect 158849 -30722 158887 -30688
rect 158921 -30722 158959 -30688
rect 158993 -30722 159031 -30688
rect 159065 -30722 159103 -30688
rect 159137 -30722 159175 -30688
rect 159209 -30722 159247 -30688
rect 159281 -30722 159319 -30688
rect 159353 -30722 159391 -30688
rect 159425 -30722 159463 -30688
rect 159497 -30722 159535 -30688
rect 159569 -30722 159607 -30688
rect 159641 -30722 159679 -30688
rect 159713 -30722 159751 -30688
rect 159785 -30722 159823 -30688
rect 159857 -30722 159895 -30688
rect 159929 -30722 159967 -30688
rect 160001 -30722 160039 -30688
rect 160073 -30722 160111 -30688
rect 160145 -30722 160183 -30688
rect 160217 -30722 160255 -30688
rect 160289 -30722 160327 -30688
rect 160361 -30722 160399 -30688
rect 160433 -30722 160471 -30688
rect 160505 -30722 160543 -30688
rect 160577 -30722 160615 -30688
rect 160649 -30722 160687 -30688
rect 160721 -30722 160759 -30688
rect 160793 -30722 160831 -30688
rect 160865 -30722 160903 -30688
rect 160937 -30722 160975 -30688
rect 161009 -30722 161047 -30688
rect 161081 -30722 161119 -30688
rect 161153 -30722 161191 -30688
rect 161225 -30722 161263 -30688
rect 161297 -30722 161335 -30688
rect 161369 -30722 161407 -30688
rect 161441 -30722 161479 -30688
rect 161513 -30722 161551 -30688
rect 161585 -30722 161623 -30688
rect 161657 -30722 161695 -30688
rect 161729 -30722 161767 -30688
rect 161801 -30722 161839 -30688
rect 161873 -30722 161911 -30688
rect 161945 -30722 161983 -30688
rect 162017 -30722 162055 -30688
rect 162089 -30722 162127 -30688
rect 162161 -30722 162199 -30688
rect 162233 -30722 162271 -30688
rect 162305 -30722 162343 -30688
rect 162377 -30722 162415 -30688
rect 162449 -30722 162487 -30688
rect 162521 -30722 162559 -30688
rect 162593 -30722 162631 -30688
rect 162665 -30722 162703 -30688
rect 162737 -30722 162775 -30688
rect 162809 -30722 162847 -30688
rect 162881 -30722 162919 -30688
rect 162953 -30722 162991 -30688
rect 163025 -30722 163063 -30688
rect 163097 -30722 163135 -30688
rect 163169 -30722 163207 -30688
rect 163241 -30722 163279 -30688
rect 163313 -30722 163351 -30688
rect 163385 -30722 163423 -30688
rect 163457 -30722 163495 -30688
rect 163529 -30722 163567 -30688
rect 163601 -30722 163639 -30688
rect 163673 -30722 163711 -30688
rect 163745 -30722 163783 -30688
rect 163817 -30722 163855 -30688
rect 163889 -30722 163927 -30688
rect 163961 -30722 163999 -30688
rect 164033 -30722 164071 -30688
rect 164105 -30722 164143 -30688
rect 164177 -30722 164215 -30688
rect 164249 -30722 164287 -30688
rect 164321 -30722 164359 -30688
rect 164393 -30722 164431 -30688
rect 164465 -30722 164503 -30688
rect 164537 -30722 164575 -30688
rect 164609 -30722 164647 -30688
rect 164681 -30722 164719 -30688
rect 164753 -30722 164791 -30688
rect 164825 -30722 164863 -30688
rect 164897 -30722 164935 -30688
rect 164969 -30722 165007 -30688
rect 165041 -30722 165079 -30688
rect 165113 -30722 165151 -30688
rect 165185 -30722 165223 -30688
rect 165257 -30722 165295 -30688
rect 165329 -30722 165367 -30688
rect 165401 -30722 165439 -30688
rect 165473 -30722 165511 -30688
rect 165545 -30722 165583 -30688
rect 165617 -30722 165655 -30688
rect 165689 -30722 165727 -30688
rect 165761 -30722 165799 -30688
rect 165833 -30722 165871 -30688
rect 165905 -30722 165943 -30688
rect 165977 -30722 166015 -30688
rect 166049 -30722 166087 -30688
rect 166121 -30722 166159 -30688
rect 166193 -30722 166231 -30688
rect 166265 -30722 166303 -30688
rect 166337 -30722 166375 -30688
rect 166409 -30722 166447 -30688
rect 166481 -30722 166519 -30688
rect 166553 -30722 166591 -30688
rect 166625 -30722 166663 -30688
rect 166697 -30722 166735 -30688
rect 166769 -30722 166807 -30688
rect 166841 -30722 166879 -30688
rect 166913 -30722 166951 -30688
rect 166985 -30722 167023 -30688
rect 167057 -30722 167095 -30688
rect 167129 -30722 167167 -30688
rect 167201 -30722 167239 -30688
rect 167273 -30722 167311 -30688
rect 167345 -30722 167383 -30688
rect 167417 -30722 167455 -30688
rect 167489 -30722 167514 -30688
rect 157854 -30726 167514 -30722
<< viali >>
rect 160381 -26118 160415 -26084
rect 160453 -26118 160487 -26084
rect 160525 -26118 160559 -26084
rect 160597 -26118 160631 -26084
rect 160669 -26118 160703 -26084
rect 160741 -26118 160775 -26084
rect 160813 -26118 160847 -26084
rect 160885 -26118 160919 -26084
rect 160957 -26118 160991 -26084
rect 161029 -26118 161063 -26084
rect 161101 -26118 161135 -26084
rect 161173 -26118 161207 -26084
rect 161245 -26118 161279 -26084
rect 161317 -26118 161351 -26084
rect 161389 -26118 161423 -26084
rect 161461 -26118 161495 -26084
rect 161533 -26118 161567 -26084
rect 161605 -26118 161639 -26084
rect 161677 -26118 161711 -26084
rect 161749 -26118 161783 -26084
rect 161821 -26118 161855 -26084
rect 161893 -26118 161927 -26084
rect 161965 -26118 161999 -26084
rect 162037 -26118 162071 -26084
rect 162109 -26118 162143 -26084
rect 162181 -26118 162215 -26084
rect 162253 -26118 162287 -26084
rect 162325 -26118 162359 -26084
rect 162397 -26118 162431 -26084
rect 162469 -26118 162503 -26084
rect 162541 -26118 162575 -26084
rect 162613 -26118 162647 -26084
rect 162685 -26118 162719 -26084
rect 162757 -26118 162791 -26084
rect 162829 -26118 162863 -26084
rect 162901 -26118 162935 -26084
rect 162973 -26118 163007 -26084
rect 163045 -26118 163079 -26084
rect 163117 -26118 163151 -26084
rect 163189 -26118 163223 -26084
rect 163261 -26118 163295 -26084
rect 163333 -26118 163367 -26084
rect 163405 -26118 163439 -26084
rect 163477 -26118 163511 -26084
rect 163549 -26118 163583 -26084
rect 163621 -26118 163655 -26084
rect 163693 -26118 163727 -26084
rect 163765 -26118 163799 -26084
rect 163837 -26118 163871 -26084
rect 163909 -26118 163943 -26084
rect 163981 -26118 164015 -26084
rect 164053 -26118 164087 -26084
rect 164125 -26118 164159 -26084
rect 164197 -26118 164231 -26084
rect 164269 -26118 164303 -26084
rect 160381 -26528 160415 -26494
rect 160453 -26528 160487 -26494
rect 160525 -26528 160559 -26494
rect 160597 -26528 160631 -26494
rect 160669 -26528 160703 -26494
rect 160741 -26528 160775 -26494
rect 160813 -26528 160847 -26494
rect 160885 -26528 160919 -26494
rect 160957 -26528 160991 -26494
rect 161029 -26528 161063 -26494
rect 161101 -26528 161135 -26494
rect 161173 -26528 161207 -26494
rect 161245 -26528 161279 -26494
rect 161317 -26528 161351 -26494
rect 161389 -26528 161423 -26494
rect 161461 -26528 161495 -26494
rect 161533 -26528 161567 -26494
rect 161605 -26528 161639 -26494
rect 161677 -26528 161711 -26494
rect 161749 -26528 161783 -26494
rect 161821 -26528 161855 -26494
rect 161893 -26528 161927 -26494
rect 161965 -26528 161999 -26494
rect 162037 -26528 162071 -26494
rect 162109 -26528 162143 -26494
rect 162181 -26528 162215 -26494
rect 162253 -26528 162287 -26494
rect 162325 -26528 162359 -26494
rect 162397 -26528 162431 -26494
rect 162469 -26528 162503 -26494
rect 162541 -26528 162575 -26494
rect 162613 -26528 162647 -26494
rect 162685 -26528 162719 -26494
rect 162757 -26528 162791 -26494
rect 162829 -26528 162863 -26494
rect 162901 -26528 162935 -26494
rect 162973 -26528 163007 -26494
rect 163045 -26528 163079 -26494
rect 163117 -26528 163151 -26494
rect 163189 -26528 163223 -26494
rect 163261 -26528 163295 -26494
rect 163333 -26528 163367 -26494
rect 163405 -26528 163439 -26494
rect 163477 -26528 163511 -26494
rect 163549 -26528 163583 -26494
rect 163621 -26528 163655 -26494
rect 163693 -26528 163727 -26494
rect 163765 -26528 163799 -26494
rect 163837 -26528 163871 -26494
rect 163909 -26528 163943 -26494
rect 163981 -26528 164015 -26494
rect 164053 -26528 164087 -26494
rect 164125 -26528 164159 -26494
rect 164197 -26528 164231 -26494
rect 164269 -26528 164303 -26494
rect 165803 -27107 165837 -27073
rect 165803 -27179 165837 -27145
rect 165803 -27251 165837 -27217
rect 165803 -27323 165837 -27289
rect 165803 -27395 165837 -27361
rect 165803 -27467 165837 -27433
rect 168665 -27107 168699 -27073
rect 168665 -27179 168699 -27145
rect 168665 -27251 168699 -27217
rect 168665 -27323 168699 -27289
rect 168665 -27395 168699 -27361
rect 168665 -27467 168699 -27433
rect 146845 -30722 146879 -30688
rect 146917 -30722 146951 -30688
rect 146989 -30722 147023 -30688
rect 147061 -30722 147095 -30688
rect 147133 -30722 147167 -30688
rect 147205 -30722 147239 -30688
rect 147277 -30722 147311 -30688
rect 147349 -30722 147383 -30688
rect 147421 -30722 147455 -30688
rect 147493 -30722 147527 -30688
rect 147565 -30722 147599 -30688
rect 147637 -30722 147671 -30688
rect 147709 -30722 147743 -30688
rect 147781 -30722 147815 -30688
rect 147853 -30722 147887 -30688
rect 147925 -30722 147959 -30688
rect 147997 -30722 148031 -30688
rect 148069 -30722 148103 -30688
rect 148141 -30722 148175 -30688
rect 148213 -30722 148247 -30688
rect 148285 -30722 148319 -30688
rect 148357 -30722 148391 -30688
rect 148429 -30722 148463 -30688
rect 148501 -30722 148535 -30688
rect 148573 -30722 148607 -30688
rect 148645 -30722 148679 -30688
rect 148717 -30722 148751 -30688
rect 148789 -30722 148823 -30688
rect 148861 -30722 148895 -30688
rect 148933 -30722 148967 -30688
rect 149005 -30722 149039 -30688
rect 149077 -30722 149111 -30688
rect 149149 -30722 149183 -30688
rect 149221 -30722 149255 -30688
rect 149293 -30722 149327 -30688
rect 149365 -30722 149399 -30688
rect 149437 -30722 149471 -30688
rect 149509 -30722 149543 -30688
rect 149581 -30722 149615 -30688
rect 149653 -30722 149687 -30688
rect 149725 -30722 149759 -30688
rect 149797 -30722 149831 -30688
rect 149869 -30722 149903 -30688
rect 149941 -30722 149975 -30688
rect 150013 -30722 150047 -30688
rect 150085 -30722 150119 -30688
rect 150157 -30722 150191 -30688
rect 150229 -30722 150263 -30688
rect 150301 -30722 150335 -30688
rect 150373 -30722 150407 -30688
rect 150445 -30722 150479 -30688
rect 150517 -30722 150551 -30688
rect 150589 -30722 150623 -30688
rect 150661 -30722 150695 -30688
rect 150733 -30722 150767 -30688
rect 150805 -30722 150839 -30688
rect 150877 -30722 150911 -30688
rect 150949 -30722 150983 -30688
rect 151021 -30722 151055 -30688
rect 151093 -30722 151127 -30688
rect 151165 -30722 151199 -30688
rect 151237 -30722 151271 -30688
rect 151309 -30722 151343 -30688
rect 151381 -30722 151415 -30688
rect 151453 -30722 151487 -30688
rect 151525 -30722 151559 -30688
rect 151597 -30722 151631 -30688
rect 151669 -30722 151703 -30688
rect 151741 -30722 151775 -30688
rect 151813 -30722 151847 -30688
rect 151885 -30722 151919 -30688
rect 151957 -30722 151991 -30688
rect 152029 -30722 152063 -30688
rect 152101 -30722 152135 -30688
rect 152173 -30722 152207 -30688
rect 152245 -30722 152279 -30688
rect 152317 -30722 152351 -30688
rect 152389 -30722 152423 -30688
rect 152461 -30722 152495 -30688
rect 152533 -30722 152567 -30688
rect 152605 -30722 152639 -30688
rect 152677 -30722 152711 -30688
rect 152749 -30722 152783 -30688
rect 152821 -30722 152855 -30688
rect 152893 -30722 152927 -30688
rect 152965 -30722 152999 -30688
rect 153037 -30722 153071 -30688
rect 153109 -30722 153143 -30688
rect 153181 -30722 153215 -30688
rect 153253 -30722 153287 -30688
rect 153325 -30722 153359 -30688
rect 153397 -30722 153431 -30688
rect 153469 -30722 153503 -30688
rect 153541 -30722 153575 -30688
rect 153613 -30722 153647 -30688
rect 153685 -30722 153719 -30688
rect 153757 -30722 153791 -30688
rect 153829 -30722 153863 -30688
rect 153901 -30722 153935 -30688
rect 153973 -30722 154007 -30688
rect 154045 -30722 154079 -30688
rect 154117 -30722 154151 -30688
rect 154189 -30722 154223 -30688
rect 154261 -30722 154295 -30688
rect 154333 -30722 154367 -30688
rect 154405 -30722 154439 -30688
rect 154477 -30722 154511 -30688
rect 154549 -30722 154583 -30688
rect 154621 -30722 154655 -30688
rect 154693 -30722 154727 -30688
rect 154765 -30722 154799 -30688
rect 154837 -30722 154871 -30688
rect 154909 -30722 154943 -30688
rect 154981 -30722 155015 -30688
rect 155053 -30722 155087 -30688
rect 155125 -30722 155159 -30688
rect 155197 -30722 155231 -30688
rect 155269 -30722 155303 -30688
rect 155341 -30722 155375 -30688
rect 155413 -30722 155447 -30688
rect 155485 -30722 155519 -30688
rect 155557 -30722 155591 -30688
rect 155629 -30722 155663 -30688
rect 155701 -30722 155735 -30688
rect 155773 -30722 155807 -30688
rect 155845 -30722 155879 -30688
rect 155917 -30722 155951 -30688
rect 155989 -30722 156023 -30688
rect 156061 -30722 156095 -30688
rect 156133 -30722 156167 -30688
rect 156205 -30722 156239 -30688
rect 156277 -30722 156311 -30688
rect 156349 -30722 156383 -30688
rect 156421 -30722 156455 -30688
rect 157879 -30722 157913 -30688
rect 157951 -30722 157985 -30688
rect 158023 -30722 158057 -30688
rect 158095 -30722 158129 -30688
rect 158167 -30722 158201 -30688
rect 158239 -30722 158273 -30688
rect 158311 -30722 158345 -30688
rect 158383 -30722 158417 -30688
rect 158455 -30722 158489 -30688
rect 158527 -30722 158561 -30688
rect 158599 -30722 158633 -30688
rect 158671 -30722 158705 -30688
rect 158743 -30722 158777 -30688
rect 158815 -30722 158849 -30688
rect 158887 -30722 158921 -30688
rect 158959 -30722 158993 -30688
rect 159031 -30722 159065 -30688
rect 159103 -30722 159137 -30688
rect 159175 -30722 159209 -30688
rect 159247 -30722 159281 -30688
rect 159319 -30722 159353 -30688
rect 159391 -30722 159425 -30688
rect 159463 -30722 159497 -30688
rect 159535 -30722 159569 -30688
rect 159607 -30722 159641 -30688
rect 159679 -30722 159713 -30688
rect 159751 -30722 159785 -30688
rect 159823 -30722 159857 -30688
rect 159895 -30722 159929 -30688
rect 159967 -30722 160001 -30688
rect 160039 -30722 160073 -30688
rect 160111 -30722 160145 -30688
rect 160183 -30722 160217 -30688
rect 160255 -30722 160289 -30688
rect 160327 -30722 160361 -30688
rect 160399 -30722 160433 -30688
rect 160471 -30722 160505 -30688
rect 160543 -30722 160577 -30688
rect 160615 -30722 160649 -30688
rect 160687 -30722 160721 -30688
rect 160759 -30722 160793 -30688
rect 160831 -30722 160865 -30688
rect 160903 -30722 160937 -30688
rect 160975 -30722 161009 -30688
rect 161047 -30722 161081 -30688
rect 161119 -30722 161153 -30688
rect 161191 -30722 161225 -30688
rect 161263 -30722 161297 -30688
rect 161335 -30722 161369 -30688
rect 161407 -30722 161441 -30688
rect 161479 -30722 161513 -30688
rect 161551 -30722 161585 -30688
rect 161623 -30722 161657 -30688
rect 161695 -30722 161729 -30688
rect 161767 -30722 161801 -30688
rect 161839 -30722 161873 -30688
rect 161911 -30722 161945 -30688
rect 161983 -30722 162017 -30688
rect 162055 -30722 162089 -30688
rect 162127 -30722 162161 -30688
rect 162199 -30722 162233 -30688
rect 162271 -30722 162305 -30688
rect 162343 -30722 162377 -30688
rect 162415 -30722 162449 -30688
rect 162487 -30722 162521 -30688
rect 162559 -30722 162593 -30688
rect 162631 -30722 162665 -30688
rect 162703 -30722 162737 -30688
rect 162775 -30722 162809 -30688
rect 162847 -30722 162881 -30688
rect 162919 -30722 162953 -30688
rect 162991 -30722 163025 -30688
rect 163063 -30722 163097 -30688
rect 163135 -30722 163169 -30688
rect 163207 -30722 163241 -30688
rect 163279 -30722 163313 -30688
rect 163351 -30722 163385 -30688
rect 163423 -30722 163457 -30688
rect 163495 -30722 163529 -30688
rect 163567 -30722 163601 -30688
rect 163639 -30722 163673 -30688
rect 163711 -30722 163745 -30688
rect 163783 -30722 163817 -30688
rect 163855 -30722 163889 -30688
rect 163927 -30722 163961 -30688
rect 163999 -30722 164033 -30688
rect 164071 -30722 164105 -30688
rect 164143 -30722 164177 -30688
rect 164215 -30722 164249 -30688
rect 164287 -30722 164321 -30688
rect 164359 -30722 164393 -30688
rect 164431 -30722 164465 -30688
rect 164503 -30722 164537 -30688
rect 164575 -30722 164609 -30688
rect 164647 -30722 164681 -30688
rect 164719 -30722 164753 -30688
rect 164791 -30722 164825 -30688
rect 164863 -30722 164897 -30688
rect 164935 -30722 164969 -30688
rect 165007 -30722 165041 -30688
rect 165079 -30722 165113 -30688
rect 165151 -30722 165185 -30688
rect 165223 -30722 165257 -30688
rect 165295 -30722 165329 -30688
rect 165367 -30722 165401 -30688
rect 165439 -30722 165473 -30688
rect 165511 -30722 165545 -30688
rect 165583 -30722 165617 -30688
rect 165655 -30722 165689 -30688
rect 165727 -30722 165761 -30688
rect 165799 -30722 165833 -30688
rect 165871 -30722 165905 -30688
rect 165943 -30722 165977 -30688
rect 166015 -30722 166049 -30688
rect 166087 -30722 166121 -30688
rect 166159 -30722 166193 -30688
rect 166231 -30722 166265 -30688
rect 166303 -30722 166337 -30688
rect 166375 -30722 166409 -30688
rect 166447 -30722 166481 -30688
rect 166519 -30722 166553 -30688
rect 166591 -30722 166625 -30688
rect 166663 -30722 166697 -30688
rect 166735 -30722 166769 -30688
rect 166807 -30722 166841 -30688
rect 166879 -30722 166913 -30688
rect 166951 -30722 166985 -30688
rect 167023 -30722 167057 -30688
rect 167095 -30722 167129 -30688
rect 167167 -30722 167201 -30688
rect 167239 -30722 167273 -30688
rect 167311 -30722 167345 -30688
rect 167383 -30722 167417 -30688
rect 167455 -30722 167489 -30688
<< metal1 >>
rect 156671 -25063 156781 -25001
rect 156671 -25115 156695 -25063
rect 156747 -25115 156781 -25063
rect 156671 -25127 156781 -25115
rect 156671 -25179 156695 -25127
rect 156747 -25179 156781 -25127
rect 156671 -25191 156781 -25179
rect 156671 -25243 156695 -25191
rect 156747 -25243 156781 -25191
rect 156671 -25255 156781 -25243
rect 156671 -25307 156695 -25255
rect 156747 -25307 156781 -25255
rect 156671 -25319 156781 -25307
rect 156671 -25371 156695 -25319
rect 156747 -25371 156781 -25319
rect 156671 -25383 156781 -25371
rect 156671 -25435 156695 -25383
rect 156747 -25435 156781 -25383
rect 156671 -25447 156781 -25435
rect 156671 -25499 156695 -25447
rect 156747 -25499 156781 -25447
rect 156671 -25511 156781 -25499
rect 156671 -25563 156695 -25511
rect 156747 -25563 156781 -25511
rect 156671 -25575 156781 -25563
rect 156671 -25627 156695 -25575
rect 156747 -25627 156781 -25575
rect 156671 -25639 156781 -25627
rect 156671 -25691 156695 -25639
rect 156747 -25691 156781 -25639
rect 156671 -25703 156781 -25691
rect 156671 -25755 156695 -25703
rect 156747 -25755 156781 -25703
rect 156671 -25767 156781 -25755
rect 156671 -25819 156695 -25767
rect 156747 -25819 156781 -25767
rect 156671 -25831 156781 -25819
rect 156671 -25883 156695 -25831
rect 156747 -25883 156781 -25831
rect 156671 -25895 156781 -25883
rect 156671 -25947 156695 -25895
rect 156747 -25947 156781 -25895
rect 156671 -25959 156781 -25947
rect 156671 -26011 156695 -25959
rect 156747 -26011 156781 -25959
rect 156671 -26023 156781 -26011
rect 156671 -26075 156695 -26023
rect 156747 -26075 156781 -26023
rect 156671 -26087 156781 -26075
rect 156671 -26139 156695 -26087
rect 156747 -26139 156781 -26087
rect 160343 -25464 164348 -25419
rect 160343 -25580 160383 -25464
rect 164275 -25580 164348 -25464
rect 160343 -26084 164348 -25580
rect 160343 -26118 160381 -26084
rect 160415 -26118 160453 -26084
rect 160487 -26118 160525 -26084
rect 160559 -26118 160597 -26084
rect 160631 -26118 160669 -26084
rect 160703 -26118 160741 -26084
rect 160775 -26118 160813 -26084
rect 160847 -26118 160885 -26084
rect 160919 -26118 160957 -26084
rect 160991 -26118 161029 -26084
rect 161063 -26118 161101 -26084
rect 161135 -26118 161173 -26084
rect 161207 -26118 161245 -26084
rect 161279 -26118 161317 -26084
rect 161351 -26118 161389 -26084
rect 161423 -26118 161461 -26084
rect 161495 -26118 161533 -26084
rect 161567 -26118 161605 -26084
rect 161639 -26118 161677 -26084
rect 161711 -26118 161749 -26084
rect 161783 -26118 161821 -26084
rect 161855 -26118 161893 -26084
rect 161927 -26118 161965 -26084
rect 161999 -26118 162037 -26084
rect 162071 -26118 162109 -26084
rect 162143 -26118 162181 -26084
rect 162215 -26118 162253 -26084
rect 162287 -26118 162325 -26084
rect 162359 -26118 162397 -26084
rect 162431 -26118 162469 -26084
rect 162503 -26118 162541 -26084
rect 162575 -26118 162613 -26084
rect 162647 -26118 162685 -26084
rect 162719 -26118 162757 -26084
rect 162791 -26118 162829 -26084
rect 162863 -26118 162901 -26084
rect 162935 -26118 162973 -26084
rect 163007 -26118 163045 -26084
rect 163079 -26118 163117 -26084
rect 163151 -26118 163189 -26084
rect 163223 -26118 163261 -26084
rect 163295 -26118 163333 -26084
rect 163367 -26118 163405 -26084
rect 163439 -26118 163477 -26084
rect 163511 -26118 163549 -26084
rect 163583 -26118 163621 -26084
rect 163655 -26118 163693 -26084
rect 163727 -26118 163765 -26084
rect 163799 -26118 163837 -26084
rect 163871 -26118 163909 -26084
rect 163943 -26118 163981 -26084
rect 164015 -26118 164053 -26084
rect 164087 -26118 164125 -26084
rect 164159 -26118 164197 -26084
rect 164231 -26118 164269 -26084
rect 164303 -26118 164348 -26084
rect 160343 -26134 164348 -26118
rect 156671 -26151 156781 -26139
rect 156671 -26203 156695 -26151
rect 156747 -26203 156781 -26151
rect 156671 -26215 156781 -26203
rect 156671 -26267 156695 -26215
rect 156747 -26267 156781 -26215
rect 156671 -26279 156781 -26267
rect 156671 -26331 156695 -26279
rect 156747 -26331 156781 -26279
rect 156671 -26343 156781 -26331
rect 156671 -26395 156695 -26343
rect 156747 -26395 156781 -26343
rect 156671 -26407 156781 -26395
rect 156671 -26459 156695 -26407
rect 156747 -26459 156781 -26407
rect 156671 -26471 156781 -26459
rect 156671 -26523 156695 -26471
rect 156747 -26523 156781 -26471
rect 156671 -26535 156781 -26523
rect 156671 -26587 156695 -26535
rect 156747 -26587 156781 -26535
rect 156671 -26599 156781 -26587
rect 156671 -26651 156695 -26599
rect 156747 -26651 156781 -26599
rect 156671 -26663 156781 -26651
rect 156671 -26715 156695 -26663
rect 156747 -26715 156781 -26663
rect 156671 -26727 156781 -26715
rect 156671 -26779 156695 -26727
rect 156747 -26779 156781 -26727
rect 156671 -26791 156781 -26779
rect 156671 -26843 156695 -26791
rect 156747 -26843 156781 -26791
rect 156671 -26855 156781 -26843
rect 156671 -26907 156695 -26855
rect 156747 -26907 156781 -26855
rect 156671 -26919 156781 -26907
rect 156671 -26971 156695 -26919
rect 156747 -26971 156781 -26919
rect 156671 -26983 156781 -26971
rect 156671 -27035 156695 -26983
rect 156747 -27035 156781 -26983
rect 156671 -27047 156781 -27035
rect 156671 -27099 156695 -27047
rect 156747 -27099 156781 -27047
rect 156671 -27111 156781 -27099
rect 156671 -27139 156695 -27111
rect 156691 -27163 156695 -27139
rect 156747 -27163 156781 -27111
rect 156691 -27179 156781 -27163
rect 156737 -27209 156781 -27179
rect 159452 -26494 164356 -26457
rect 159452 -26528 160381 -26494
rect 160415 -26528 160453 -26494
rect 160487 -26528 160525 -26494
rect 160559 -26528 160597 -26494
rect 160631 -26528 160669 -26494
rect 160703 -26528 160741 -26494
rect 160775 -26528 160813 -26494
rect 160847 -26528 160885 -26494
rect 160919 -26528 160957 -26494
rect 160991 -26528 161029 -26494
rect 161063 -26528 161101 -26494
rect 161135 -26528 161173 -26494
rect 161207 -26528 161245 -26494
rect 161279 -26528 161317 -26494
rect 161351 -26528 161389 -26494
rect 161423 -26528 161461 -26494
rect 161495 -26528 161533 -26494
rect 161567 -26528 161605 -26494
rect 161639 -26528 161677 -26494
rect 161711 -26528 161749 -26494
rect 161783 -26528 161821 -26494
rect 161855 -26528 161893 -26494
rect 161927 -26528 161965 -26494
rect 161999 -26528 162037 -26494
rect 162071 -26528 162109 -26494
rect 162143 -26528 162181 -26494
rect 162215 -26528 162253 -26494
rect 162287 -26528 162325 -26494
rect 162359 -26528 162397 -26494
rect 162431 -26528 162469 -26494
rect 162503 -26528 162541 -26494
rect 162575 -26528 162613 -26494
rect 162647 -26528 162685 -26494
rect 162719 -26528 162757 -26494
rect 162791 -26528 162829 -26494
rect 162863 -26528 162901 -26494
rect 162935 -26528 162973 -26494
rect 163007 -26528 163045 -26494
rect 163079 -26528 163117 -26494
rect 163151 -26528 163189 -26494
rect 163223 -26528 163261 -26494
rect 163295 -26528 163333 -26494
rect 163367 -26528 163405 -26494
rect 163439 -26528 163477 -26494
rect 163511 -26528 163549 -26494
rect 163583 -26528 163621 -26494
rect 163655 -26528 163693 -26494
rect 163727 -26528 163765 -26494
rect 163799 -26528 163837 -26494
rect 163871 -26528 163909 -26494
rect 163943 -26528 163981 -26494
rect 164015 -26528 164053 -26494
rect 164087 -26528 164125 -26494
rect 164159 -26528 164197 -26494
rect 164231 -26528 164269 -26494
rect 164303 -26528 164356 -26494
rect 159452 -27008 164356 -26528
rect 159452 -27073 165892 -27008
rect 159452 -27107 165803 -27073
rect 165837 -27107 165892 -27073
rect 159452 -27145 165892 -27107
rect 159452 -27179 165803 -27145
rect 165837 -27179 165892 -27145
rect 159452 -27217 165892 -27179
rect 159452 -27251 165803 -27217
rect 165837 -27251 165892 -27217
rect 159452 -27289 165892 -27251
rect 159452 -27323 165803 -27289
rect 165837 -27323 165892 -27289
rect 159452 -27361 165892 -27323
rect 159452 -27395 165803 -27361
rect 165837 -27395 165892 -27361
rect 159452 -27433 165892 -27395
rect 159452 -27461 165803 -27433
rect 157051 -27462 165803 -27461
rect 156707 -27467 165803 -27462
rect 165837 -27467 165892 -27433
rect 156707 -27567 165892 -27467
rect 168611 -27073 168750 -27022
rect 168611 -27107 168665 -27073
rect 168699 -27107 168750 -27073
rect 168611 -27145 168750 -27107
rect 168611 -27179 168665 -27145
rect 168699 -27179 168750 -27145
rect 168611 -27217 168750 -27179
rect 168611 -27251 168665 -27217
rect 168699 -27251 168750 -27217
rect 168611 -27289 168750 -27251
rect 168611 -27323 168665 -27289
rect 168699 -27323 168750 -27289
rect 168611 -27361 168750 -27323
rect 168611 -27395 168665 -27361
rect 168699 -27395 168750 -27361
rect 168611 -27433 168750 -27395
rect 168611 -27467 168665 -27433
rect 168699 -27467 168750 -27433
rect 156707 -27951 164356 -27567
rect 168611 -27925 168750 -27467
rect 156707 -29795 157450 -27951
rect 166918 -27981 169100 -27925
rect 166918 -28088 168806 -27981
rect 166918 -28140 166962 -28088
rect 167014 -28140 167026 -28088
rect 167078 -28140 167090 -28088
rect 167142 -28140 167154 -28088
rect 167206 -28140 167218 -28088
rect 167270 -28140 167282 -28088
rect 167334 -28140 167346 -28088
rect 167398 -28140 167410 -28088
rect 167462 -28140 167474 -28088
rect 167526 -28140 167538 -28088
rect 167590 -28140 168806 -28088
rect 166918 -28161 168806 -28140
rect 169050 -28161 169100 -27981
rect 166918 -28213 169100 -28161
rect 166918 -28506 167630 -28213
rect 146808 -30688 156508 -30672
rect 146808 -30722 146845 -30688
rect 146879 -30722 146917 -30688
rect 146951 -30722 146989 -30688
rect 147023 -30722 147061 -30688
rect 147095 -30722 147133 -30688
rect 147167 -30722 147205 -30688
rect 147239 -30722 147277 -30688
rect 147311 -30722 147349 -30688
rect 147383 -30722 147421 -30688
rect 147455 -30722 147493 -30688
rect 147527 -30722 147565 -30688
rect 147599 -30722 147637 -30688
rect 147671 -30722 147709 -30688
rect 147743 -30722 147781 -30688
rect 147815 -30722 147853 -30688
rect 147887 -30722 147925 -30688
rect 147959 -30722 147997 -30688
rect 148031 -30722 148069 -30688
rect 148103 -30722 148141 -30688
rect 148175 -30722 148213 -30688
rect 148247 -30722 148285 -30688
rect 148319 -30722 148357 -30688
rect 148391 -30722 148429 -30688
rect 148463 -30722 148501 -30688
rect 148535 -30722 148573 -30688
rect 148607 -30722 148645 -30688
rect 148679 -30722 148717 -30688
rect 148751 -30722 148789 -30688
rect 148823 -30722 148861 -30688
rect 148895 -30722 148933 -30688
rect 148967 -30722 149005 -30688
rect 149039 -30722 149077 -30688
rect 149111 -30722 149149 -30688
rect 149183 -30722 149221 -30688
rect 149255 -30722 149293 -30688
rect 149327 -30722 149365 -30688
rect 149399 -30722 149437 -30688
rect 149471 -30722 149509 -30688
rect 149543 -30722 149581 -30688
rect 149615 -30722 149653 -30688
rect 149687 -30722 149725 -30688
rect 149759 -30722 149797 -30688
rect 149831 -30722 149869 -30688
rect 149903 -30722 149941 -30688
rect 149975 -30722 150013 -30688
rect 150047 -30722 150085 -30688
rect 150119 -30722 150157 -30688
rect 150191 -30722 150229 -30688
rect 150263 -30722 150301 -30688
rect 150335 -30722 150373 -30688
rect 150407 -30722 150445 -30688
rect 150479 -30722 150517 -30688
rect 150551 -30722 150589 -30688
rect 150623 -30722 150661 -30688
rect 150695 -30722 150733 -30688
rect 150767 -30722 150805 -30688
rect 150839 -30722 150877 -30688
rect 150911 -30722 150949 -30688
rect 150983 -30722 151021 -30688
rect 151055 -30722 151093 -30688
rect 151127 -30722 151165 -30688
rect 151199 -30722 151237 -30688
rect 151271 -30722 151309 -30688
rect 151343 -30722 151381 -30688
rect 151415 -30722 151453 -30688
rect 151487 -30722 151525 -30688
rect 151559 -30722 151597 -30688
rect 151631 -30722 151669 -30688
rect 151703 -30722 151741 -30688
rect 151775 -30722 151813 -30688
rect 151847 -30722 151885 -30688
rect 151919 -30722 151957 -30688
rect 151991 -30722 152029 -30688
rect 152063 -30722 152101 -30688
rect 152135 -30722 152173 -30688
rect 152207 -30722 152245 -30688
rect 152279 -30722 152317 -30688
rect 152351 -30722 152389 -30688
rect 152423 -30722 152461 -30688
rect 152495 -30722 152533 -30688
rect 152567 -30722 152605 -30688
rect 152639 -30722 152677 -30688
rect 152711 -30722 152749 -30688
rect 152783 -30722 152821 -30688
rect 152855 -30722 152893 -30688
rect 152927 -30722 152965 -30688
rect 152999 -30722 153037 -30688
rect 153071 -30722 153109 -30688
rect 153143 -30722 153181 -30688
rect 153215 -30722 153253 -30688
rect 153287 -30722 153325 -30688
rect 153359 -30722 153397 -30688
rect 153431 -30722 153469 -30688
rect 153503 -30722 153541 -30688
rect 153575 -30722 153613 -30688
rect 153647 -30722 153685 -30688
rect 153719 -30722 153757 -30688
rect 153791 -30722 153829 -30688
rect 153863 -30722 153901 -30688
rect 153935 -30722 153973 -30688
rect 154007 -30722 154045 -30688
rect 154079 -30722 154117 -30688
rect 154151 -30722 154189 -30688
rect 154223 -30722 154261 -30688
rect 154295 -30722 154333 -30688
rect 154367 -30722 154405 -30688
rect 154439 -30722 154477 -30688
rect 154511 -30722 154549 -30688
rect 154583 -30722 154621 -30688
rect 154655 -30722 154693 -30688
rect 154727 -30722 154765 -30688
rect 154799 -30722 154837 -30688
rect 154871 -30722 154909 -30688
rect 154943 -30722 154981 -30688
rect 155015 -30722 155053 -30688
rect 155087 -30722 155125 -30688
rect 155159 -30722 155197 -30688
rect 155231 -30722 155269 -30688
rect 155303 -30722 155341 -30688
rect 155375 -30722 155413 -30688
rect 155447 -30722 155485 -30688
rect 155519 -30722 155557 -30688
rect 155591 -30722 155629 -30688
rect 155663 -30722 155701 -30688
rect 155735 -30722 155773 -30688
rect 155807 -30722 155845 -30688
rect 155879 -30722 155917 -30688
rect 155951 -30722 155989 -30688
rect 156023 -30722 156061 -30688
rect 156095 -30722 156133 -30688
rect 156167 -30722 156205 -30688
rect 156239 -30722 156277 -30688
rect 156311 -30722 156349 -30688
rect 156383 -30722 156421 -30688
rect 156455 -30722 156508 -30688
rect 146808 -30732 156508 -30722
rect 146802 -30748 156508 -30732
rect 157842 -30688 167562 -30674
rect 157842 -30722 157879 -30688
rect 157913 -30722 157951 -30688
rect 157985 -30722 158023 -30688
rect 158057 -30722 158095 -30688
rect 158129 -30722 158167 -30688
rect 158201 -30722 158239 -30688
rect 158273 -30722 158311 -30688
rect 158345 -30722 158383 -30688
rect 158417 -30722 158455 -30688
rect 158489 -30722 158527 -30688
rect 158561 -30722 158599 -30688
rect 158633 -30722 158671 -30688
rect 158705 -30722 158743 -30688
rect 158777 -30722 158815 -30688
rect 158849 -30722 158887 -30688
rect 158921 -30722 158959 -30688
rect 158993 -30722 159031 -30688
rect 159065 -30722 159103 -30688
rect 159137 -30722 159175 -30688
rect 159209 -30722 159247 -30688
rect 159281 -30722 159319 -30688
rect 159353 -30722 159391 -30688
rect 159425 -30722 159463 -30688
rect 159497 -30722 159535 -30688
rect 159569 -30722 159607 -30688
rect 159641 -30722 159679 -30688
rect 159713 -30722 159751 -30688
rect 159785 -30722 159823 -30688
rect 159857 -30722 159895 -30688
rect 159929 -30722 159967 -30688
rect 160001 -30722 160039 -30688
rect 160073 -30722 160111 -30688
rect 160145 -30722 160183 -30688
rect 160217 -30722 160255 -30688
rect 160289 -30722 160327 -30688
rect 160361 -30722 160399 -30688
rect 160433 -30722 160471 -30688
rect 160505 -30722 160543 -30688
rect 160577 -30722 160615 -30688
rect 160649 -30722 160687 -30688
rect 160721 -30722 160759 -30688
rect 160793 -30722 160831 -30688
rect 160865 -30722 160903 -30688
rect 160937 -30722 160975 -30688
rect 161009 -30722 161047 -30688
rect 161081 -30722 161119 -30688
rect 161153 -30722 161191 -30688
rect 161225 -30722 161263 -30688
rect 161297 -30722 161335 -30688
rect 161369 -30722 161407 -30688
rect 161441 -30722 161479 -30688
rect 161513 -30722 161551 -30688
rect 161585 -30722 161623 -30688
rect 161657 -30722 161695 -30688
rect 161729 -30722 161767 -30688
rect 161801 -30722 161839 -30688
rect 161873 -30722 161911 -30688
rect 161945 -30722 161983 -30688
rect 162017 -30722 162055 -30688
rect 162089 -30722 162127 -30688
rect 162161 -30722 162199 -30688
rect 162233 -30722 162271 -30688
rect 162305 -30722 162343 -30688
rect 162377 -30722 162415 -30688
rect 162449 -30722 162487 -30688
rect 162521 -30722 162559 -30688
rect 162593 -30722 162631 -30688
rect 162665 -30722 162703 -30688
rect 162737 -30722 162775 -30688
rect 162809 -30722 162847 -30688
rect 162881 -30722 162919 -30688
rect 162953 -30722 162991 -30688
rect 163025 -30722 163063 -30688
rect 163097 -30722 163135 -30688
rect 163169 -30722 163207 -30688
rect 163241 -30722 163279 -30688
rect 163313 -30722 163351 -30688
rect 163385 -30722 163423 -30688
rect 163457 -30722 163495 -30688
rect 163529 -30722 163567 -30688
rect 163601 -30722 163639 -30688
rect 163673 -30722 163711 -30688
rect 163745 -30722 163783 -30688
rect 163817 -30722 163855 -30688
rect 163889 -30722 163927 -30688
rect 163961 -30722 163999 -30688
rect 164033 -30722 164071 -30688
rect 164105 -30722 164143 -30688
rect 164177 -30722 164215 -30688
rect 164249 -30722 164287 -30688
rect 164321 -30722 164359 -30688
rect 164393 -30722 164431 -30688
rect 164465 -30722 164503 -30688
rect 164537 -30722 164575 -30688
rect 164609 -30722 164647 -30688
rect 164681 -30722 164719 -30688
rect 164753 -30722 164791 -30688
rect 164825 -30722 164863 -30688
rect 164897 -30722 164935 -30688
rect 164969 -30722 165007 -30688
rect 165041 -30722 165079 -30688
rect 165113 -30722 165151 -30688
rect 165185 -30722 165223 -30688
rect 165257 -30722 165295 -30688
rect 165329 -30722 165367 -30688
rect 165401 -30722 165439 -30688
rect 165473 -30722 165511 -30688
rect 165545 -30722 165583 -30688
rect 165617 -30722 165655 -30688
rect 165689 -30722 165727 -30688
rect 165761 -30722 165799 -30688
rect 165833 -30722 165871 -30688
rect 165905 -30722 165943 -30688
rect 165977 -30722 166015 -30688
rect 166049 -30722 166087 -30688
rect 166121 -30722 166159 -30688
rect 166193 -30722 166231 -30688
rect 166265 -30722 166303 -30688
rect 166337 -30722 166375 -30688
rect 166409 -30722 166447 -30688
rect 166481 -30722 166519 -30688
rect 166553 -30722 166591 -30688
rect 166625 -30722 166663 -30688
rect 166697 -30722 166735 -30688
rect 166769 -30722 166807 -30688
rect 166841 -30722 166879 -30688
rect 166913 -30722 166951 -30688
rect 166985 -30722 167023 -30688
rect 167057 -30722 167095 -30688
rect 167129 -30722 167167 -30688
rect 167201 -30722 167239 -30688
rect 167273 -30722 167311 -30688
rect 167345 -30722 167383 -30688
rect 167417 -30722 167455 -30688
rect 167489 -30722 167562 -30688
rect 157842 -30748 167562 -30722
rect 146802 -30868 167562 -30748
rect 146802 -30876 157897 -30868
rect 146802 -30928 146843 -30876
rect 146895 -30928 146907 -30876
rect 146959 -30928 146971 -30876
rect 147023 -30928 147035 -30876
rect 147087 -30928 147099 -30876
rect 147151 -30928 147163 -30876
rect 147215 -30928 147227 -30876
rect 147279 -30928 147291 -30876
rect 147343 -30928 147355 -30876
rect 147407 -30928 147419 -30876
rect 147471 -30928 147483 -30876
rect 147535 -30928 147547 -30876
rect 147599 -30928 147611 -30876
rect 147663 -30928 147675 -30876
rect 147727 -30928 147739 -30876
rect 147791 -30928 147803 -30876
rect 147855 -30928 147867 -30876
rect 147919 -30928 147931 -30876
rect 147983 -30928 147995 -30876
rect 148047 -30928 148059 -30876
rect 148111 -30928 148123 -30876
rect 148175 -30928 148187 -30876
rect 148239 -30928 148251 -30876
rect 148303 -30928 148315 -30876
rect 148367 -30928 148379 -30876
rect 148431 -30928 148443 -30876
rect 148495 -30928 148507 -30876
rect 148559 -30928 148571 -30876
rect 148623 -30928 148635 -30876
rect 148687 -30928 148699 -30876
rect 148751 -30928 148763 -30876
rect 148815 -30928 148827 -30876
rect 148879 -30928 148891 -30876
rect 148943 -30928 148955 -30876
rect 149007 -30928 149019 -30876
rect 149071 -30928 149083 -30876
rect 149135 -30928 149147 -30876
rect 149199 -30928 149211 -30876
rect 149263 -30928 149275 -30876
rect 149327 -30928 149339 -30876
rect 149391 -30928 149403 -30876
rect 149455 -30928 149467 -30876
rect 149519 -30928 149531 -30876
rect 149583 -30928 149595 -30876
rect 149647 -30928 149659 -30876
rect 149711 -30928 149723 -30876
rect 149775 -30928 149787 -30876
rect 149839 -30928 149851 -30876
rect 149903 -30928 149915 -30876
rect 149967 -30928 149979 -30876
rect 150031 -30928 150043 -30876
rect 150095 -30928 150107 -30876
rect 150159 -30928 150171 -30876
rect 150223 -30928 150235 -30876
rect 150287 -30928 150299 -30876
rect 150351 -30928 150363 -30876
rect 150415 -30928 150427 -30876
rect 150479 -30928 150491 -30876
rect 150543 -30928 150555 -30876
rect 150607 -30928 150619 -30876
rect 150671 -30928 150683 -30876
rect 150735 -30928 150747 -30876
rect 150799 -30928 150811 -30876
rect 150863 -30928 150875 -30876
rect 150927 -30928 150939 -30876
rect 150991 -30928 151003 -30876
rect 151055 -30928 151067 -30876
rect 151119 -30928 151131 -30876
rect 151183 -30928 151195 -30876
rect 151247 -30928 151259 -30876
rect 151311 -30928 151323 -30876
rect 151375 -30928 151387 -30876
rect 151439 -30928 151451 -30876
rect 151503 -30928 151515 -30876
rect 151567 -30928 151579 -30876
rect 151631 -30928 151643 -30876
rect 151695 -30928 151707 -30876
rect 151759 -30928 151771 -30876
rect 151823 -30928 151835 -30876
rect 151887 -30928 151899 -30876
rect 151951 -30928 151963 -30876
rect 152015 -30928 152027 -30876
rect 152079 -30928 152091 -30876
rect 152143 -30928 152155 -30876
rect 152207 -30928 152219 -30876
rect 152271 -30928 152283 -30876
rect 152335 -30928 152347 -30876
rect 152399 -30928 152411 -30876
rect 152463 -30928 152475 -30876
rect 152527 -30928 152539 -30876
rect 152591 -30928 152603 -30876
rect 152655 -30928 152667 -30876
rect 152719 -30928 152731 -30876
rect 152783 -30928 152795 -30876
rect 152847 -30928 152859 -30876
rect 152911 -30928 152923 -30876
rect 152975 -30928 152987 -30876
rect 153039 -30928 153051 -30876
rect 153103 -30928 153115 -30876
rect 153167 -30928 153179 -30876
rect 153231 -30928 153243 -30876
rect 153295 -30928 153307 -30876
rect 153359 -30928 153371 -30876
rect 153423 -30928 153435 -30876
rect 153487 -30928 153499 -30876
rect 153551 -30928 153563 -30876
rect 153615 -30928 153627 -30876
rect 153679 -30928 153691 -30876
rect 153743 -30928 153755 -30876
rect 153807 -30928 153819 -30876
rect 153871 -30928 153883 -30876
rect 153935 -30928 153947 -30876
rect 153999 -30928 154011 -30876
rect 154063 -30928 154075 -30876
rect 154127 -30928 154139 -30876
rect 154191 -30928 154203 -30876
rect 154255 -30928 154267 -30876
rect 154319 -30928 154331 -30876
rect 154383 -30928 154395 -30876
rect 154447 -30928 154459 -30876
rect 154511 -30928 154523 -30876
rect 154575 -30928 154587 -30876
rect 154639 -30928 154651 -30876
rect 154703 -30928 154715 -30876
rect 154767 -30928 154779 -30876
rect 154831 -30928 154843 -30876
rect 154895 -30928 154907 -30876
rect 154959 -30928 154971 -30876
rect 155023 -30928 155035 -30876
rect 155087 -30928 155099 -30876
rect 155151 -30928 155163 -30876
rect 155215 -30928 155227 -30876
rect 155279 -30928 155291 -30876
rect 155343 -30928 155355 -30876
rect 155407 -30928 155419 -30876
rect 155471 -30928 155483 -30876
rect 155535 -30928 155547 -30876
rect 155599 -30928 155611 -30876
rect 155663 -30928 155675 -30876
rect 155727 -30928 155739 -30876
rect 155791 -30928 155803 -30876
rect 155855 -30928 155867 -30876
rect 155919 -30928 155931 -30876
rect 155983 -30928 155995 -30876
rect 156047 -30928 156059 -30876
rect 156111 -30928 156123 -30876
rect 156175 -30928 156187 -30876
rect 156239 -30928 156251 -30876
rect 156303 -30928 156315 -30876
rect 156367 -30928 156379 -30876
rect 156431 -30920 157897 -30876
rect 157949 -30920 157961 -30868
rect 158013 -30920 158025 -30868
rect 158077 -30920 158089 -30868
rect 158141 -30920 158153 -30868
rect 158205 -30920 158217 -30868
rect 158269 -30920 158281 -30868
rect 158333 -30920 158345 -30868
rect 158397 -30920 158409 -30868
rect 158461 -30920 158473 -30868
rect 158525 -30920 158537 -30868
rect 158589 -30920 158601 -30868
rect 158653 -30920 158665 -30868
rect 158717 -30920 158729 -30868
rect 158781 -30920 158793 -30868
rect 158845 -30920 158857 -30868
rect 158909 -30920 158921 -30868
rect 158973 -30920 158985 -30868
rect 159037 -30920 159049 -30868
rect 159101 -30920 159113 -30868
rect 159165 -30920 159177 -30868
rect 159229 -30920 159241 -30868
rect 159293 -30920 159305 -30868
rect 159357 -30920 159369 -30868
rect 159421 -30920 159433 -30868
rect 159485 -30920 159497 -30868
rect 159549 -30920 159561 -30868
rect 159613 -30920 159625 -30868
rect 159677 -30920 159689 -30868
rect 159741 -30920 159753 -30868
rect 159805 -30920 159817 -30868
rect 159869 -30920 159881 -30868
rect 159933 -30920 159945 -30868
rect 159997 -30920 160009 -30868
rect 160061 -30920 160073 -30868
rect 160125 -30920 160137 -30868
rect 160189 -30920 160201 -30868
rect 160253 -30920 160265 -30868
rect 160317 -30920 160329 -30868
rect 160381 -30920 160393 -30868
rect 160445 -30920 160457 -30868
rect 160509 -30920 160521 -30868
rect 160573 -30920 160585 -30868
rect 160637 -30920 160649 -30868
rect 160701 -30920 160713 -30868
rect 160765 -30920 160777 -30868
rect 160829 -30920 160841 -30868
rect 160893 -30920 160905 -30868
rect 160957 -30920 160969 -30868
rect 161021 -30920 161033 -30868
rect 161085 -30920 161097 -30868
rect 161149 -30920 161161 -30868
rect 161213 -30920 161225 -30868
rect 161277 -30920 161289 -30868
rect 161341 -30920 161353 -30868
rect 161405 -30920 161417 -30868
rect 161469 -30920 161481 -30868
rect 161533 -30920 161545 -30868
rect 161597 -30920 161609 -30868
rect 161661 -30920 161673 -30868
rect 161725 -30920 161737 -30868
rect 161789 -30920 161801 -30868
rect 161853 -30920 161865 -30868
rect 161917 -30920 161929 -30868
rect 161981 -30920 161993 -30868
rect 162045 -30920 162057 -30868
rect 162109 -30920 162121 -30868
rect 162173 -30920 162185 -30868
rect 162237 -30920 162249 -30868
rect 162301 -30920 162313 -30868
rect 162365 -30920 162377 -30868
rect 162429 -30920 162441 -30868
rect 162493 -30920 162505 -30868
rect 162557 -30920 162569 -30868
rect 162621 -30920 162633 -30868
rect 162685 -30920 162697 -30868
rect 162749 -30920 162761 -30868
rect 162813 -30920 162825 -30868
rect 162877 -30920 162889 -30868
rect 162941 -30920 162953 -30868
rect 163005 -30920 163017 -30868
rect 163069 -30920 163081 -30868
rect 163133 -30920 163145 -30868
rect 163197 -30920 163209 -30868
rect 163261 -30920 163273 -30868
rect 163325 -30920 163337 -30868
rect 163389 -30920 163401 -30868
rect 163453 -30920 163465 -30868
rect 163517 -30920 163529 -30868
rect 163581 -30920 163593 -30868
rect 163645 -30920 163657 -30868
rect 163709 -30920 163721 -30868
rect 163773 -30920 163785 -30868
rect 163837 -30920 163849 -30868
rect 163901 -30920 163913 -30868
rect 163965 -30920 163977 -30868
rect 164029 -30920 164041 -30868
rect 164093 -30920 164105 -30868
rect 164157 -30920 164169 -30868
rect 164221 -30920 164233 -30868
rect 164285 -30920 164297 -30868
rect 164349 -30920 164361 -30868
rect 164413 -30920 164425 -30868
rect 164477 -30920 164489 -30868
rect 164541 -30920 164553 -30868
rect 164605 -30920 164617 -30868
rect 164669 -30920 164681 -30868
rect 164733 -30920 164745 -30868
rect 164797 -30920 164809 -30868
rect 164861 -30920 164873 -30868
rect 164925 -30920 164937 -30868
rect 164989 -30920 165001 -30868
rect 165053 -30920 165065 -30868
rect 165117 -30920 165129 -30868
rect 165181 -30920 165193 -30868
rect 165245 -30920 165257 -30868
rect 165309 -30920 165321 -30868
rect 165373 -30920 165385 -30868
rect 165437 -30920 165449 -30868
rect 165501 -30920 165513 -30868
rect 165565 -30920 165577 -30868
rect 165629 -30920 165641 -30868
rect 165693 -30920 165705 -30868
rect 165757 -30920 165769 -30868
rect 165821 -30920 165833 -30868
rect 165885 -30920 165897 -30868
rect 165949 -30920 165961 -30868
rect 166013 -30920 166025 -30868
rect 166077 -30920 166089 -30868
rect 166141 -30920 166153 -30868
rect 166205 -30920 166217 -30868
rect 166269 -30920 166281 -30868
rect 166333 -30920 166345 -30868
rect 166397 -30920 166409 -30868
rect 166461 -30920 166473 -30868
rect 166525 -30920 166537 -30868
rect 166589 -30920 166601 -30868
rect 166653 -30920 166665 -30868
rect 166717 -30920 166729 -30868
rect 166781 -30920 166793 -30868
rect 166845 -30920 166857 -30868
rect 166909 -30920 166921 -30868
rect 166973 -30920 166985 -30868
rect 167037 -30920 167049 -30868
rect 167101 -30920 167113 -30868
rect 167165 -30920 167177 -30868
rect 167229 -30920 167241 -30868
rect 167293 -30920 167305 -30868
rect 167357 -30920 167369 -30868
rect 167421 -30920 167433 -30868
rect 167485 -30920 167562 -30868
rect 156431 -30928 167562 -30920
rect 146802 -30944 167562 -30928
rect 146802 -30952 157862 -30944
<< via1 >>
rect 156695 -25115 156747 -25063
rect 156695 -25179 156747 -25127
rect 156695 -25243 156747 -25191
rect 156695 -25307 156747 -25255
rect 156695 -25371 156747 -25319
rect 156695 -25435 156747 -25383
rect 156695 -25499 156747 -25447
rect 156695 -25563 156747 -25511
rect 156695 -25627 156747 -25575
rect 156695 -25691 156747 -25639
rect 156695 -25755 156747 -25703
rect 156695 -25819 156747 -25767
rect 156695 -25883 156747 -25831
rect 156695 -25947 156747 -25895
rect 156695 -26011 156747 -25959
rect 156695 -26075 156747 -26023
rect 156695 -26139 156747 -26087
rect 160383 -25580 164275 -25464
rect 156695 -26203 156747 -26151
rect 156695 -26267 156747 -26215
rect 156695 -26331 156747 -26279
rect 156695 -26395 156747 -26343
rect 156695 -26459 156747 -26407
rect 156695 -26523 156747 -26471
rect 156695 -26587 156747 -26535
rect 156695 -26651 156747 -26599
rect 156695 -26715 156747 -26663
rect 156695 -26779 156747 -26727
rect 156695 -26843 156747 -26791
rect 156695 -26907 156747 -26855
rect 156695 -26971 156747 -26919
rect 156695 -27035 156747 -26983
rect 156695 -27099 156747 -27047
rect 156695 -27163 156747 -27111
rect 166962 -28140 167014 -28088
rect 167026 -28140 167078 -28088
rect 167090 -28140 167142 -28088
rect 167154 -28140 167206 -28088
rect 167218 -28140 167270 -28088
rect 167282 -28140 167334 -28088
rect 167346 -28140 167398 -28088
rect 167410 -28140 167462 -28088
rect 167474 -28140 167526 -28088
rect 167538 -28140 167590 -28088
rect 168806 -28161 169050 -27981
rect 146843 -30928 146895 -30876
rect 146907 -30928 146959 -30876
rect 146971 -30928 147023 -30876
rect 147035 -30928 147087 -30876
rect 147099 -30928 147151 -30876
rect 147163 -30928 147215 -30876
rect 147227 -30928 147279 -30876
rect 147291 -30928 147343 -30876
rect 147355 -30928 147407 -30876
rect 147419 -30928 147471 -30876
rect 147483 -30928 147535 -30876
rect 147547 -30928 147599 -30876
rect 147611 -30928 147663 -30876
rect 147675 -30928 147727 -30876
rect 147739 -30928 147791 -30876
rect 147803 -30928 147855 -30876
rect 147867 -30928 147919 -30876
rect 147931 -30928 147983 -30876
rect 147995 -30928 148047 -30876
rect 148059 -30928 148111 -30876
rect 148123 -30928 148175 -30876
rect 148187 -30928 148239 -30876
rect 148251 -30928 148303 -30876
rect 148315 -30928 148367 -30876
rect 148379 -30928 148431 -30876
rect 148443 -30928 148495 -30876
rect 148507 -30928 148559 -30876
rect 148571 -30928 148623 -30876
rect 148635 -30928 148687 -30876
rect 148699 -30928 148751 -30876
rect 148763 -30928 148815 -30876
rect 148827 -30928 148879 -30876
rect 148891 -30928 148943 -30876
rect 148955 -30928 149007 -30876
rect 149019 -30928 149071 -30876
rect 149083 -30928 149135 -30876
rect 149147 -30928 149199 -30876
rect 149211 -30928 149263 -30876
rect 149275 -30928 149327 -30876
rect 149339 -30928 149391 -30876
rect 149403 -30928 149455 -30876
rect 149467 -30928 149519 -30876
rect 149531 -30928 149583 -30876
rect 149595 -30928 149647 -30876
rect 149659 -30928 149711 -30876
rect 149723 -30928 149775 -30876
rect 149787 -30928 149839 -30876
rect 149851 -30928 149903 -30876
rect 149915 -30928 149967 -30876
rect 149979 -30928 150031 -30876
rect 150043 -30928 150095 -30876
rect 150107 -30928 150159 -30876
rect 150171 -30928 150223 -30876
rect 150235 -30928 150287 -30876
rect 150299 -30928 150351 -30876
rect 150363 -30928 150415 -30876
rect 150427 -30928 150479 -30876
rect 150491 -30928 150543 -30876
rect 150555 -30928 150607 -30876
rect 150619 -30928 150671 -30876
rect 150683 -30928 150735 -30876
rect 150747 -30928 150799 -30876
rect 150811 -30928 150863 -30876
rect 150875 -30928 150927 -30876
rect 150939 -30928 150991 -30876
rect 151003 -30928 151055 -30876
rect 151067 -30928 151119 -30876
rect 151131 -30928 151183 -30876
rect 151195 -30928 151247 -30876
rect 151259 -30928 151311 -30876
rect 151323 -30928 151375 -30876
rect 151387 -30928 151439 -30876
rect 151451 -30928 151503 -30876
rect 151515 -30928 151567 -30876
rect 151579 -30928 151631 -30876
rect 151643 -30928 151695 -30876
rect 151707 -30928 151759 -30876
rect 151771 -30928 151823 -30876
rect 151835 -30928 151887 -30876
rect 151899 -30928 151951 -30876
rect 151963 -30928 152015 -30876
rect 152027 -30928 152079 -30876
rect 152091 -30928 152143 -30876
rect 152155 -30928 152207 -30876
rect 152219 -30928 152271 -30876
rect 152283 -30928 152335 -30876
rect 152347 -30928 152399 -30876
rect 152411 -30928 152463 -30876
rect 152475 -30928 152527 -30876
rect 152539 -30928 152591 -30876
rect 152603 -30928 152655 -30876
rect 152667 -30928 152719 -30876
rect 152731 -30928 152783 -30876
rect 152795 -30928 152847 -30876
rect 152859 -30928 152911 -30876
rect 152923 -30928 152975 -30876
rect 152987 -30928 153039 -30876
rect 153051 -30928 153103 -30876
rect 153115 -30928 153167 -30876
rect 153179 -30928 153231 -30876
rect 153243 -30928 153295 -30876
rect 153307 -30928 153359 -30876
rect 153371 -30928 153423 -30876
rect 153435 -30928 153487 -30876
rect 153499 -30928 153551 -30876
rect 153563 -30928 153615 -30876
rect 153627 -30928 153679 -30876
rect 153691 -30928 153743 -30876
rect 153755 -30928 153807 -30876
rect 153819 -30928 153871 -30876
rect 153883 -30928 153935 -30876
rect 153947 -30928 153999 -30876
rect 154011 -30928 154063 -30876
rect 154075 -30928 154127 -30876
rect 154139 -30928 154191 -30876
rect 154203 -30928 154255 -30876
rect 154267 -30928 154319 -30876
rect 154331 -30928 154383 -30876
rect 154395 -30928 154447 -30876
rect 154459 -30928 154511 -30876
rect 154523 -30928 154575 -30876
rect 154587 -30928 154639 -30876
rect 154651 -30928 154703 -30876
rect 154715 -30928 154767 -30876
rect 154779 -30928 154831 -30876
rect 154843 -30928 154895 -30876
rect 154907 -30928 154959 -30876
rect 154971 -30928 155023 -30876
rect 155035 -30928 155087 -30876
rect 155099 -30928 155151 -30876
rect 155163 -30928 155215 -30876
rect 155227 -30928 155279 -30876
rect 155291 -30928 155343 -30876
rect 155355 -30928 155407 -30876
rect 155419 -30928 155471 -30876
rect 155483 -30928 155535 -30876
rect 155547 -30928 155599 -30876
rect 155611 -30928 155663 -30876
rect 155675 -30928 155727 -30876
rect 155739 -30928 155791 -30876
rect 155803 -30928 155855 -30876
rect 155867 -30928 155919 -30876
rect 155931 -30928 155983 -30876
rect 155995 -30928 156047 -30876
rect 156059 -30928 156111 -30876
rect 156123 -30928 156175 -30876
rect 156187 -30928 156239 -30876
rect 156251 -30928 156303 -30876
rect 156315 -30928 156367 -30876
rect 156379 -30928 156431 -30876
rect 157897 -30920 157949 -30868
rect 157961 -30920 158013 -30868
rect 158025 -30920 158077 -30868
rect 158089 -30920 158141 -30868
rect 158153 -30920 158205 -30868
rect 158217 -30920 158269 -30868
rect 158281 -30920 158333 -30868
rect 158345 -30920 158397 -30868
rect 158409 -30920 158461 -30868
rect 158473 -30920 158525 -30868
rect 158537 -30920 158589 -30868
rect 158601 -30920 158653 -30868
rect 158665 -30920 158717 -30868
rect 158729 -30920 158781 -30868
rect 158793 -30920 158845 -30868
rect 158857 -30920 158909 -30868
rect 158921 -30920 158973 -30868
rect 158985 -30920 159037 -30868
rect 159049 -30920 159101 -30868
rect 159113 -30920 159165 -30868
rect 159177 -30920 159229 -30868
rect 159241 -30920 159293 -30868
rect 159305 -30920 159357 -30868
rect 159369 -30920 159421 -30868
rect 159433 -30920 159485 -30868
rect 159497 -30920 159549 -30868
rect 159561 -30920 159613 -30868
rect 159625 -30920 159677 -30868
rect 159689 -30920 159741 -30868
rect 159753 -30920 159805 -30868
rect 159817 -30920 159869 -30868
rect 159881 -30920 159933 -30868
rect 159945 -30920 159997 -30868
rect 160009 -30920 160061 -30868
rect 160073 -30920 160125 -30868
rect 160137 -30920 160189 -30868
rect 160201 -30920 160253 -30868
rect 160265 -30920 160317 -30868
rect 160329 -30920 160381 -30868
rect 160393 -30920 160445 -30868
rect 160457 -30920 160509 -30868
rect 160521 -30920 160573 -30868
rect 160585 -30920 160637 -30868
rect 160649 -30920 160701 -30868
rect 160713 -30920 160765 -30868
rect 160777 -30920 160829 -30868
rect 160841 -30920 160893 -30868
rect 160905 -30920 160957 -30868
rect 160969 -30920 161021 -30868
rect 161033 -30920 161085 -30868
rect 161097 -30920 161149 -30868
rect 161161 -30920 161213 -30868
rect 161225 -30920 161277 -30868
rect 161289 -30920 161341 -30868
rect 161353 -30920 161405 -30868
rect 161417 -30920 161469 -30868
rect 161481 -30920 161533 -30868
rect 161545 -30920 161597 -30868
rect 161609 -30920 161661 -30868
rect 161673 -30920 161725 -30868
rect 161737 -30920 161789 -30868
rect 161801 -30920 161853 -30868
rect 161865 -30920 161917 -30868
rect 161929 -30920 161981 -30868
rect 161993 -30920 162045 -30868
rect 162057 -30920 162109 -30868
rect 162121 -30920 162173 -30868
rect 162185 -30920 162237 -30868
rect 162249 -30920 162301 -30868
rect 162313 -30920 162365 -30868
rect 162377 -30920 162429 -30868
rect 162441 -30920 162493 -30868
rect 162505 -30920 162557 -30868
rect 162569 -30920 162621 -30868
rect 162633 -30920 162685 -30868
rect 162697 -30920 162749 -30868
rect 162761 -30920 162813 -30868
rect 162825 -30920 162877 -30868
rect 162889 -30920 162941 -30868
rect 162953 -30920 163005 -30868
rect 163017 -30920 163069 -30868
rect 163081 -30920 163133 -30868
rect 163145 -30920 163197 -30868
rect 163209 -30920 163261 -30868
rect 163273 -30920 163325 -30868
rect 163337 -30920 163389 -30868
rect 163401 -30920 163453 -30868
rect 163465 -30920 163517 -30868
rect 163529 -30920 163581 -30868
rect 163593 -30920 163645 -30868
rect 163657 -30920 163709 -30868
rect 163721 -30920 163773 -30868
rect 163785 -30920 163837 -30868
rect 163849 -30920 163901 -30868
rect 163913 -30920 163965 -30868
rect 163977 -30920 164029 -30868
rect 164041 -30920 164093 -30868
rect 164105 -30920 164157 -30868
rect 164169 -30920 164221 -30868
rect 164233 -30920 164285 -30868
rect 164297 -30920 164349 -30868
rect 164361 -30920 164413 -30868
rect 164425 -30920 164477 -30868
rect 164489 -30920 164541 -30868
rect 164553 -30920 164605 -30868
rect 164617 -30920 164669 -30868
rect 164681 -30920 164733 -30868
rect 164745 -30920 164797 -30868
rect 164809 -30920 164861 -30868
rect 164873 -30920 164925 -30868
rect 164937 -30920 164989 -30868
rect 165001 -30920 165053 -30868
rect 165065 -30920 165117 -30868
rect 165129 -30920 165181 -30868
rect 165193 -30920 165245 -30868
rect 165257 -30920 165309 -30868
rect 165321 -30920 165373 -30868
rect 165385 -30920 165437 -30868
rect 165449 -30920 165501 -30868
rect 165513 -30920 165565 -30868
rect 165577 -30920 165629 -30868
rect 165641 -30920 165693 -30868
rect 165705 -30920 165757 -30868
rect 165769 -30920 165821 -30868
rect 165833 -30920 165885 -30868
rect 165897 -30920 165949 -30868
rect 165961 -30920 166013 -30868
rect 166025 -30920 166077 -30868
rect 166089 -30920 166141 -30868
rect 166153 -30920 166205 -30868
rect 166217 -30920 166269 -30868
rect 166281 -30920 166333 -30868
rect 166345 -30920 166397 -30868
rect 166409 -30920 166461 -30868
rect 166473 -30920 166525 -30868
rect 166537 -30920 166589 -30868
rect 166601 -30920 166653 -30868
rect 166665 -30920 166717 -30868
rect 166729 -30920 166781 -30868
rect 166793 -30920 166845 -30868
rect 166857 -30920 166909 -30868
rect 166921 -30920 166973 -30868
rect 166985 -30920 167037 -30868
rect 167049 -30920 167101 -30868
rect 167113 -30920 167165 -30868
rect 167177 -30920 167229 -30868
rect 167241 -30920 167293 -30868
rect 167305 -30920 167357 -30868
rect 167369 -30920 167421 -30868
rect 167433 -30920 167485 -30868
<< metal2 >>
rect 156671 -20655 158155 -20476
rect 156671 -21591 156793 -20655
rect 158049 -21591 158155 -20655
rect 156671 -25063 158155 -21591
rect 156671 -25115 156695 -25063
rect 156747 -25115 158155 -25063
rect 156671 -25127 158155 -25115
rect 156671 -25179 156695 -25127
rect 156747 -25179 158155 -25127
rect 156671 -25191 158155 -25179
rect 156671 -25243 156695 -25191
rect 156747 -25243 158155 -25191
rect 156671 -25255 158155 -25243
rect 156671 -25307 156695 -25255
rect 156747 -25307 158155 -25255
rect 156671 -25319 158155 -25307
rect 156671 -25371 156695 -25319
rect 156747 -25371 158155 -25319
rect 156671 -25383 158155 -25371
rect 156671 -25435 156695 -25383
rect 156747 -25435 158155 -25383
rect 156671 -25447 158155 -25435
rect 156671 -25499 156695 -25447
rect 156747 -25499 158155 -25447
rect 156671 -25511 158155 -25499
rect 156671 -25563 156695 -25511
rect 156747 -25563 158155 -25511
rect 156671 -25575 158155 -25563
rect 156671 -25627 156695 -25575
rect 156747 -25627 158155 -25575
rect 160343 -25029 164348 -24939
rect 160343 -25085 160442 -25029
rect 160498 -25085 160522 -25029
rect 160578 -25085 160602 -25029
rect 160658 -25085 160682 -25029
rect 160738 -25085 160762 -25029
rect 160818 -25085 160842 -25029
rect 160898 -25085 160922 -25029
rect 160978 -25085 161002 -25029
rect 161058 -25085 161082 -25029
rect 161138 -25085 161162 -25029
rect 161218 -25085 161242 -25029
rect 161298 -25085 161322 -25029
rect 161378 -25085 161402 -25029
rect 161458 -25085 161482 -25029
rect 161538 -25085 161562 -25029
rect 161618 -25085 161642 -25029
rect 161698 -25085 161722 -25029
rect 161778 -25085 161802 -25029
rect 161858 -25085 161882 -25029
rect 161938 -25085 161962 -25029
rect 162018 -25085 162042 -25029
rect 162098 -25085 162122 -25029
rect 162178 -25085 162202 -25029
rect 162258 -25085 162282 -25029
rect 162338 -25085 162362 -25029
rect 162418 -25085 162442 -25029
rect 162498 -25085 162522 -25029
rect 162578 -25085 162602 -25029
rect 162658 -25085 162682 -25029
rect 162738 -25085 162762 -25029
rect 162818 -25085 162842 -25029
rect 162898 -25085 162922 -25029
rect 162978 -25085 163002 -25029
rect 163058 -25085 163082 -25029
rect 163138 -25085 163162 -25029
rect 163218 -25085 163242 -25029
rect 163298 -25085 163322 -25029
rect 163378 -25085 163402 -25029
rect 163458 -25085 163482 -25029
rect 163538 -25085 163562 -25029
rect 163618 -25085 163642 -25029
rect 163698 -25085 163722 -25029
rect 163778 -25085 163802 -25029
rect 163858 -25085 163882 -25029
rect 163938 -25085 163962 -25029
rect 164018 -25085 164042 -25029
rect 164098 -25085 164122 -25029
rect 164178 -25085 164202 -25029
rect 164258 -25085 164348 -25029
rect 160343 -25464 164348 -25085
rect 160343 -25580 160383 -25464
rect 164275 -25580 164348 -25464
rect 160343 -25604 164348 -25580
rect 156671 -25639 158155 -25627
rect 156671 -25691 156695 -25639
rect 156747 -25691 158155 -25639
rect 156671 -25703 158155 -25691
rect 156671 -25755 156695 -25703
rect 156747 -25755 158155 -25703
rect 156671 -25767 158155 -25755
rect 156671 -25819 156695 -25767
rect 156747 -25819 158155 -25767
rect 156671 -25831 158155 -25819
rect 156671 -25883 156695 -25831
rect 156747 -25883 158155 -25831
rect 156671 -25895 158155 -25883
rect 156671 -25947 156695 -25895
rect 156747 -25947 158155 -25895
rect 156671 -25959 158155 -25947
rect 156671 -26011 156695 -25959
rect 156747 -26011 158155 -25959
rect 156671 -26023 158155 -26011
rect 156671 -26075 156695 -26023
rect 156747 -26075 158155 -26023
rect 156671 -26087 158155 -26075
rect 156671 -26139 156695 -26087
rect 156747 -26139 158155 -26087
rect 156671 -26151 158155 -26139
rect 156671 -26203 156695 -26151
rect 156747 -26203 158155 -26151
rect 156671 -26215 158155 -26203
rect 156671 -26267 156695 -26215
rect 156747 -26267 158155 -26215
rect 156671 -26279 158155 -26267
rect 156671 -26331 156695 -26279
rect 156747 -26331 158155 -26279
rect 156671 -26343 158155 -26331
rect 156671 -26395 156695 -26343
rect 156747 -26395 158155 -26343
rect 156671 -26407 158155 -26395
rect 156671 -26459 156695 -26407
rect 156747 -26459 158155 -26407
rect 156671 -26471 158155 -26459
rect 156671 -26523 156695 -26471
rect 156747 -26523 158155 -26471
rect 156671 -26535 158155 -26523
rect 156671 -26587 156695 -26535
rect 156747 -26587 158155 -26535
rect 156671 -26599 158155 -26587
rect 156671 -26651 156695 -26599
rect 156747 -26651 158155 -26599
rect 156671 -26663 158155 -26651
rect 156671 -26715 156695 -26663
rect 156747 -26715 158155 -26663
rect 156671 -26727 158155 -26715
rect 156671 -26779 156695 -26727
rect 156747 -26779 158155 -26727
rect 156671 -26791 158155 -26779
rect 156671 -26843 156695 -26791
rect 156747 -26843 158155 -26791
rect 156671 -26855 158155 -26843
rect 156671 -26907 156695 -26855
rect 156747 -26907 158155 -26855
rect 156671 -26919 158155 -26907
rect 156671 -26971 156695 -26919
rect 156747 -26971 158155 -26919
rect 156671 -26983 158155 -26971
rect 156671 -27035 156695 -26983
rect 156747 -27035 158155 -26983
rect 156671 -27047 158155 -27035
rect 156671 -27099 156695 -27047
rect 156747 -27099 158155 -27047
rect 156671 -27111 158155 -27099
rect 156671 -27163 156695 -27111
rect 156747 -27163 158155 -27111
rect 156671 -27209 158155 -27163
rect 146934 -27441 156410 -27440
rect 146934 -27497 146964 -27441
rect 147020 -27497 147044 -27441
rect 147100 -27497 147124 -27441
rect 147180 -27497 147204 -27441
rect 147260 -27497 147284 -27441
rect 147340 -27497 147364 -27441
rect 147420 -27497 147444 -27441
rect 147500 -27497 147524 -27441
rect 147580 -27497 147604 -27441
rect 147660 -27497 147684 -27441
rect 147740 -27497 147764 -27441
rect 147820 -27497 147844 -27441
rect 147900 -27497 147924 -27441
rect 147980 -27497 148004 -27441
rect 148060 -27497 148084 -27441
rect 148140 -27497 148164 -27441
rect 148220 -27497 148244 -27441
rect 148300 -27497 148324 -27441
rect 148380 -27497 148404 -27441
rect 148460 -27497 148484 -27441
rect 148540 -27497 148564 -27441
rect 148620 -27497 148644 -27441
rect 148700 -27497 148724 -27441
rect 148780 -27497 148804 -27441
rect 148860 -27497 148884 -27441
rect 148940 -27497 148964 -27441
rect 149020 -27497 149044 -27441
rect 149100 -27497 149124 -27441
rect 149180 -27497 149204 -27441
rect 149260 -27497 149284 -27441
rect 149340 -27497 149364 -27441
rect 149420 -27497 149444 -27441
rect 149500 -27497 149524 -27441
rect 149580 -27497 149604 -27441
rect 149660 -27497 149684 -27441
rect 149740 -27497 149764 -27441
rect 149820 -27497 149844 -27441
rect 149900 -27497 149924 -27441
rect 149980 -27497 150004 -27441
rect 150060 -27497 150084 -27441
rect 150140 -27497 150164 -27441
rect 150220 -27497 150244 -27441
rect 150300 -27497 150324 -27441
rect 150380 -27497 150404 -27441
rect 150460 -27497 150484 -27441
rect 150540 -27497 150564 -27441
rect 150620 -27497 150644 -27441
rect 150700 -27497 150724 -27441
rect 150780 -27497 150804 -27441
rect 150860 -27497 150884 -27441
rect 150940 -27497 150964 -27441
rect 151020 -27497 151044 -27441
rect 151100 -27497 151124 -27441
rect 151180 -27497 151204 -27441
rect 151260 -27497 151284 -27441
rect 151340 -27497 151364 -27441
rect 151420 -27497 151444 -27441
rect 151500 -27497 151524 -27441
rect 151580 -27497 151604 -27441
rect 151660 -27497 151684 -27441
rect 151740 -27497 151764 -27441
rect 151820 -27497 151844 -27441
rect 151900 -27497 151924 -27441
rect 151980 -27497 152004 -27441
rect 152060 -27497 152084 -27441
rect 152140 -27497 152164 -27441
rect 152220 -27497 152244 -27441
rect 152300 -27497 152324 -27441
rect 152380 -27497 152404 -27441
rect 152460 -27497 152484 -27441
rect 152540 -27497 152564 -27441
rect 152620 -27497 152644 -27441
rect 152700 -27497 152724 -27441
rect 152780 -27497 152804 -27441
rect 152860 -27497 152884 -27441
rect 152940 -27497 152964 -27441
rect 153020 -27497 153044 -27441
rect 153100 -27497 153124 -27441
rect 153180 -27497 153204 -27441
rect 153260 -27497 153284 -27441
rect 153340 -27497 153364 -27441
rect 153420 -27497 153444 -27441
rect 153500 -27497 153524 -27441
rect 153580 -27497 153604 -27441
rect 153660 -27497 153684 -27441
rect 153740 -27497 153764 -27441
rect 153820 -27497 153844 -27441
rect 153900 -27497 153924 -27441
rect 153980 -27497 154004 -27441
rect 154060 -27497 154084 -27441
rect 154140 -27497 154164 -27441
rect 154220 -27497 154244 -27441
rect 154300 -27497 154324 -27441
rect 154380 -27497 154404 -27441
rect 154460 -27497 154484 -27441
rect 154540 -27497 154564 -27441
rect 154620 -27497 154644 -27441
rect 154700 -27497 154724 -27441
rect 154780 -27497 154804 -27441
rect 154860 -27497 154884 -27441
rect 154940 -27497 154964 -27441
rect 155020 -27497 155044 -27441
rect 155100 -27497 155124 -27441
rect 155180 -27497 155204 -27441
rect 155260 -27497 155284 -27441
rect 155340 -27497 155364 -27441
rect 155420 -27497 155444 -27441
rect 155500 -27497 155524 -27441
rect 155580 -27497 155604 -27441
rect 155660 -27497 155684 -27441
rect 155740 -27497 155764 -27441
rect 155820 -27497 155844 -27441
rect 155900 -27497 155924 -27441
rect 155980 -27497 156004 -27441
rect 156060 -27497 156084 -27441
rect 156140 -27497 156164 -27441
rect 156220 -27497 156244 -27441
rect 156300 -27497 156324 -27441
rect 156380 -27497 156410 -27441
rect 146934 -27498 156410 -27497
rect 168769 -27961 169780 -27925
rect 168769 -27981 169494 -27961
rect 166901 -28088 167652 -28062
rect 166901 -28140 166962 -28088
rect 167014 -28096 167026 -28088
rect 167078 -28096 167090 -28088
rect 167142 -28096 167154 -28088
rect 167206 -28096 167218 -28088
rect 167023 -28140 167026 -28096
rect 167206 -28140 167207 -28096
rect 167270 -28140 167282 -28088
rect 167334 -28096 167346 -28088
rect 167398 -28096 167410 -28088
rect 167462 -28096 167474 -28088
rect 167526 -28096 167538 -28088
rect 167343 -28140 167346 -28096
rect 167526 -28140 167527 -28096
rect 167590 -28140 167652 -28088
rect 166901 -28152 166967 -28140
rect 167023 -28152 167047 -28140
rect 167103 -28152 167127 -28140
rect 167183 -28152 167207 -28140
rect 167263 -28152 167287 -28140
rect 167343 -28152 167367 -28140
rect 167423 -28152 167447 -28140
rect 167503 -28152 167527 -28140
rect 167583 -28152 167652 -28140
rect 166901 -28196 167652 -28152
rect 168769 -28161 168806 -27981
rect 169050 -28161 169494 -27981
rect 168769 -28177 169494 -28161
rect 169710 -28177 169780 -27961
rect 168769 -28213 169780 -28177
rect 146820 -30868 167519 -30855
rect 146820 -30876 157897 -30868
rect 146820 -30928 146843 -30876
rect 146895 -30928 146907 -30876
rect 146959 -30928 146971 -30876
rect 147023 -30928 147035 -30876
rect 147087 -30928 147099 -30876
rect 147151 -30928 147163 -30876
rect 147215 -30928 147227 -30876
rect 147279 -30928 147291 -30876
rect 147343 -30928 147355 -30876
rect 147407 -30928 147419 -30876
rect 147471 -30928 147483 -30876
rect 147535 -30928 147547 -30876
rect 147599 -30928 147611 -30876
rect 147663 -30928 147675 -30876
rect 147727 -30928 147739 -30876
rect 147791 -30928 147803 -30876
rect 147855 -30928 147867 -30876
rect 147919 -30928 147931 -30876
rect 147983 -30928 147995 -30876
rect 148047 -30928 148059 -30876
rect 148111 -30928 148123 -30876
rect 148175 -30928 148187 -30876
rect 148239 -30928 148251 -30876
rect 148303 -30928 148315 -30876
rect 148367 -30928 148379 -30876
rect 148431 -30928 148443 -30876
rect 148495 -30928 148507 -30876
rect 148559 -30928 148571 -30876
rect 148623 -30928 148635 -30876
rect 148687 -30928 148699 -30876
rect 148751 -30928 148763 -30876
rect 148815 -30928 148827 -30876
rect 148879 -30928 148891 -30876
rect 148943 -30928 148955 -30876
rect 149007 -30928 149019 -30876
rect 149071 -30928 149083 -30876
rect 149135 -30928 149147 -30876
rect 149199 -30928 149211 -30876
rect 149263 -30928 149275 -30876
rect 149327 -30928 149339 -30876
rect 149391 -30928 149403 -30876
rect 149455 -30928 149467 -30876
rect 149519 -30928 149531 -30876
rect 149583 -30928 149595 -30876
rect 149647 -30928 149659 -30876
rect 149711 -30928 149723 -30876
rect 149775 -30928 149787 -30876
rect 149839 -30928 149851 -30876
rect 149903 -30928 149915 -30876
rect 149967 -30928 149979 -30876
rect 150031 -30928 150043 -30876
rect 150095 -30928 150107 -30876
rect 150159 -30928 150171 -30876
rect 150223 -30928 150235 -30876
rect 150287 -30928 150299 -30876
rect 150351 -30928 150363 -30876
rect 150415 -30928 150427 -30876
rect 150479 -30928 150491 -30876
rect 150543 -30928 150555 -30876
rect 150607 -30928 150619 -30876
rect 150671 -30928 150683 -30876
rect 150735 -30928 150747 -30876
rect 150799 -30928 150811 -30876
rect 150863 -30928 150875 -30876
rect 150927 -30928 150939 -30876
rect 150991 -30928 151003 -30876
rect 151055 -30928 151067 -30876
rect 151119 -30928 151131 -30876
rect 151183 -30928 151195 -30876
rect 151247 -30928 151259 -30876
rect 151311 -30928 151323 -30876
rect 151375 -30928 151387 -30876
rect 151439 -30928 151451 -30876
rect 151503 -30928 151515 -30876
rect 151567 -30928 151579 -30876
rect 151631 -30928 151643 -30876
rect 151695 -30928 151707 -30876
rect 151759 -30928 151771 -30876
rect 151823 -30928 151835 -30876
rect 151887 -30928 151899 -30876
rect 151951 -30928 151963 -30876
rect 152015 -30928 152027 -30876
rect 152079 -30928 152091 -30876
rect 152143 -30928 152155 -30876
rect 152207 -30928 152219 -30876
rect 152271 -30928 152283 -30876
rect 152335 -30928 152347 -30876
rect 152399 -30928 152411 -30876
rect 152463 -30928 152475 -30876
rect 152527 -30928 152539 -30876
rect 152591 -30928 152603 -30876
rect 152655 -30928 152667 -30876
rect 152719 -30928 152731 -30876
rect 152783 -30928 152795 -30876
rect 152847 -30928 152859 -30876
rect 152911 -30928 152923 -30876
rect 152975 -30928 152987 -30876
rect 153039 -30928 153051 -30876
rect 153103 -30928 153115 -30876
rect 153167 -30928 153179 -30876
rect 153231 -30928 153243 -30876
rect 153295 -30928 153307 -30876
rect 153359 -30928 153371 -30876
rect 153423 -30928 153435 -30876
rect 153487 -30928 153499 -30876
rect 153551 -30928 153563 -30876
rect 153615 -30928 153627 -30876
rect 153679 -30928 153691 -30876
rect 153743 -30928 153755 -30876
rect 153807 -30928 153819 -30876
rect 153871 -30928 153883 -30876
rect 153935 -30928 153947 -30876
rect 153999 -30928 154011 -30876
rect 154063 -30928 154075 -30876
rect 154127 -30928 154139 -30876
rect 154191 -30928 154203 -30876
rect 154255 -30928 154267 -30876
rect 154319 -30928 154331 -30876
rect 154383 -30928 154395 -30876
rect 154447 -30928 154459 -30876
rect 154511 -30928 154523 -30876
rect 154575 -30928 154587 -30876
rect 154639 -30928 154651 -30876
rect 154703 -30928 154715 -30876
rect 154767 -30928 154779 -30876
rect 154831 -30928 154843 -30876
rect 154895 -30928 154907 -30876
rect 154959 -30928 154971 -30876
rect 155023 -30928 155035 -30876
rect 155087 -30928 155099 -30876
rect 155151 -30928 155163 -30876
rect 155215 -30928 155227 -30876
rect 155279 -30928 155291 -30876
rect 155343 -30928 155355 -30876
rect 155407 -30928 155419 -30876
rect 155471 -30928 155483 -30876
rect 155535 -30928 155547 -30876
rect 155599 -30928 155611 -30876
rect 155663 -30928 155675 -30876
rect 155727 -30928 155739 -30876
rect 155791 -30928 155803 -30876
rect 155855 -30928 155867 -30876
rect 155919 -30928 155931 -30876
rect 155983 -30928 155995 -30876
rect 156047 -30928 156059 -30876
rect 156111 -30928 156123 -30876
rect 156175 -30928 156187 -30876
rect 156239 -30928 156251 -30876
rect 156303 -30928 156315 -30876
rect 156367 -30928 156379 -30876
rect 156431 -30920 157897 -30876
rect 157949 -30920 157961 -30868
rect 158013 -30920 158025 -30868
rect 158077 -30920 158089 -30868
rect 158141 -30920 158153 -30868
rect 158205 -30920 158217 -30868
rect 158269 -30920 158281 -30868
rect 158333 -30920 158345 -30868
rect 158397 -30920 158409 -30868
rect 158461 -30920 158473 -30868
rect 158525 -30920 158537 -30868
rect 158589 -30920 158601 -30868
rect 158653 -30920 158665 -30868
rect 158717 -30920 158729 -30868
rect 158781 -30920 158793 -30868
rect 158845 -30920 158857 -30868
rect 158909 -30920 158921 -30868
rect 158973 -30920 158985 -30868
rect 159037 -30920 159049 -30868
rect 159101 -30920 159113 -30868
rect 159165 -30920 159177 -30868
rect 159229 -30920 159241 -30868
rect 159293 -30920 159305 -30868
rect 159357 -30920 159369 -30868
rect 159421 -30920 159433 -30868
rect 159485 -30920 159497 -30868
rect 159549 -30920 159561 -30868
rect 159613 -30920 159625 -30868
rect 159677 -30920 159689 -30868
rect 159741 -30920 159753 -30868
rect 159805 -30920 159817 -30868
rect 159869 -30920 159881 -30868
rect 159933 -30920 159945 -30868
rect 159997 -30920 160009 -30868
rect 160061 -30920 160073 -30868
rect 160125 -30920 160137 -30868
rect 160189 -30920 160201 -30868
rect 160253 -30920 160265 -30868
rect 160317 -30920 160329 -30868
rect 160381 -30920 160393 -30868
rect 160445 -30920 160457 -30868
rect 160509 -30920 160521 -30868
rect 160573 -30920 160585 -30868
rect 160637 -30920 160649 -30868
rect 160701 -30920 160713 -30868
rect 160765 -30920 160777 -30868
rect 160829 -30920 160841 -30868
rect 160893 -30920 160905 -30868
rect 160957 -30920 160969 -30868
rect 161021 -30920 161033 -30868
rect 161085 -30920 161097 -30868
rect 161149 -30920 161161 -30868
rect 161213 -30920 161225 -30868
rect 161277 -30920 161289 -30868
rect 161341 -30920 161353 -30868
rect 161405 -30920 161417 -30868
rect 161469 -30920 161481 -30868
rect 161533 -30920 161545 -30868
rect 161597 -30920 161609 -30868
rect 161661 -30920 161673 -30868
rect 161725 -30920 161737 -30868
rect 161789 -30920 161801 -30868
rect 161853 -30920 161865 -30868
rect 161917 -30920 161929 -30868
rect 161981 -30920 161993 -30868
rect 162045 -30920 162057 -30868
rect 162109 -30920 162121 -30868
rect 162173 -30920 162185 -30868
rect 162237 -30920 162249 -30868
rect 162301 -30920 162313 -30868
rect 162365 -30920 162377 -30868
rect 162429 -30920 162441 -30868
rect 162493 -30920 162505 -30868
rect 162557 -30920 162569 -30868
rect 162621 -30920 162633 -30868
rect 162685 -30920 162697 -30868
rect 162749 -30920 162761 -30868
rect 162813 -30920 162825 -30868
rect 162877 -30920 162889 -30868
rect 162941 -30920 162953 -30868
rect 163005 -30920 163017 -30868
rect 163069 -30920 163081 -30868
rect 163133 -30920 163145 -30868
rect 163197 -30920 163209 -30868
rect 163261 -30920 163273 -30868
rect 163325 -30920 163337 -30868
rect 163389 -30920 163401 -30868
rect 163453 -30920 163465 -30868
rect 163517 -30920 163529 -30868
rect 163581 -30920 163593 -30868
rect 163645 -30920 163657 -30868
rect 163709 -30920 163721 -30868
rect 163773 -30920 163785 -30868
rect 163837 -30920 163849 -30868
rect 163901 -30920 163913 -30868
rect 163965 -30920 163977 -30868
rect 164029 -30920 164041 -30868
rect 164093 -30920 164105 -30868
rect 164157 -30920 164169 -30868
rect 164221 -30920 164233 -30868
rect 164285 -30920 164297 -30868
rect 164349 -30920 164361 -30868
rect 164413 -30920 164425 -30868
rect 164477 -30920 164489 -30868
rect 164541 -30920 164553 -30868
rect 164605 -30920 164617 -30868
rect 164669 -30920 164681 -30868
rect 164733 -30920 164745 -30868
rect 164797 -30920 164809 -30868
rect 164861 -30920 164873 -30868
rect 164925 -30920 164937 -30868
rect 164989 -30920 165001 -30868
rect 165053 -30920 165065 -30868
rect 165117 -30920 165129 -30868
rect 165181 -30920 165193 -30868
rect 165245 -30920 165257 -30868
rect 165309 -30920 165321 -30868
rect 165373 -30920 165385 -30868
rect 165437 -30920 165449 -30868
rect 165501 -30920 165513 -30868
rect 165565 -30920 165577 -30868
rect 165629 -30920 165641 -30868
rect 165693 -30920 165705 -30868
rect 165757 -30920 165769 -30868
rect 165821 -30920 165833 -30868
rect 165885 -30920 165897 -30868
rect 165949 -30920 165961 -30868
rect 166013 -30920 166025 -30868
rect 166077 -30920 166089 -30868
rect 166141 -30920 166153 -30868
rect 166205 -30920 166217 -30868
rect 166269 -30920 166281 -30868
rect 166333 -30920 166345 -30868
rect 166397 -30920 166409 -30868
rect 166461 -30920 166473 -30868
rect 166525 -30920 166537 -30868
rect 166589 -30920 166601 -30868
rect 166653 -30920 166665 -30868
rect 166717 -30920 166729 -30868
rect 166781 -30920 166793 -30868
rect 166845 -30920 166857 -30868
rect 166909 -30920 166921 -30868
rect 166973 -30920 166985 -30868
rect 167037 -30920 167049 -30868
rect 167101 -30920 167113 -30868
rect 167165 -30920 167177 -30868
rect 167229 -30920 167241 -30868
rect 167293 -30920 167305 -30868
rect 167357 -30920 167369 -30868
rect 167421 -30920 167433 -30868
rect 167485 -30920 167519 -30868
rect 156431 -30928 167519 -30920
rect 146820 -31380 167519 -30928
rect 146820 -31516 146865 -31380
rect 167401 -31516 167519 -31380
rect 146820 -31558 167519 -31516
<< via2 >>
rect 156793 -21591 158049 -20655
rect 160442 -25085 160498 -25029
rect 160522 -25085 160578 -25029
rect 160602 -25085 160658 -25029
rect 160682 -25085 160738 -25029
rect 160762 -25085 160818 -25029
rect 160842 -25085 160898 -25029
rect 160922 -25085 160978 -25029
rect 161002 -25085 161058 -25029
rect 161082 -25085 161138 -25029
rect 161162 -25085 161218 -25029
rect 161242 -25085 161298 -25029
rect 161322 -25085 161378 -25029
rect 161402 -25085 161458 -25029
rect 161482 -25085 161538 -25029
rect 161562 -25085 161618 -25029
rect 161642 -25085 161698 -25029
rect 161722 -25085 161778 -25029
rect 161802 -25085 161858 -25029
rect 161882 -25085 161938 -25029
rect 161962 -25085 162018 -25029
rect 162042 -25085 162098 -25029
rect 162122 -25085 162178 -25029
rect 162202 -25085 162258 -25029
rect 162282 -25085 162338 -25029
rect 162362 -25085 162418 -25029
rect 162442 -25085 162498 -25029
rect 162522 -25085 162578 -25029
rect 162602 -25085 162658 -25029
rect 162682 -25085 162738 -25029
rect 162762 -25085 162818 -25029
rect 162842 -25085 162898 -25029
rect 162922 -25085 162978 -25029
rect 163002 -25085 163058 -25029
rect 163082 -25085 163138 -25029
rect 163162 -25085 163218 -25029
rect 163242 -25085 163298 -25029
rect 163322 -25085 163378 -25029
rect 163402 -25085 163458 -25029
rect 163482 -25085 163538 -25029
rect 163562 -25085 163618 -25029
rect 163642 -25085 163698 -25029
rect 163722 -25085 163778 -25029
rect 163802 -25085 163858 -25029
rect 163882 -25085 163938 -25029
rect 163962 -25085 164018 -25029
rect 164042 -25085 164098 -25029
rect 164122 -25085 164178 -25029
rect 164202 -25085 164258 -25029
rect 146964 -27497 147020 -27441
rect 147044 -27497 147100 -27441
rect 147124 -27497 147180 -27441
rect 147204 -27497 147260 -27441
rect 147284 -27497 147340 -27441
rect 147364 -27497 147420 -27441
rect 147444 -27497 147500 -27441
rect 147524 -27497 147580 -27441
rect 147604 -27497 147660 -27441
rect 147684 -27497 147740 -27441
rect 147764 -27497 147820 -27441
rect 147844 -27497 147900 -27441
rect 147924 -27497 147980 -27441
rect 148004 -27497 148060 -27441
rect 148084 -27497 148140 -27441
rect 148164 -27497 148220 -27441
rect 148244 -27497 148300 -27441
rect 148324 -27497 148380 -27441
rect 148404 -27497 148460 -27441
rect 148484 -27497 148540 -27441
rect 148564 -27497 148620 -27441
rect 148644 -27497 148700 -27441
rect 148724 -27497 148780 -27441
rect 148804 -27497 148860 -27441
rect 148884 -27497 148940 -27441
rect 148964 -27497 149020 -27441
rect 149044 -27497 149100 -27441
rect 149124 -27497 149180 -27441
rect 149204 -27497 149260 -27441
rect 149284 -27497 149340 -27441
rect 149364 -27497 149420 -27441
rect 149444 -27497 149500 -27441
rect 149524 -27497 149580 -27441
rect 149604 -27497 149660 -27441
rect 149684 -27497 149740 -27441
rect 149764 -27497 149820 -27441
rect 149844 -27497 149900 -27441
rect 149924 -27497 149980 -27441
rect 150004 -27497 150060 -27441
rect 150084 -27497 150140 -27441
rect 150164 -27497 150220 -27441
rect 150244 -27497 150300 -27441
rect 150324 -27497 150380 -27441
rect 150404 -27497 150460 -27441
rect 150484 -27497 150540 -27441
rect 150564 -27497 150620 -27441
rect 150644 -27497 150700 -27441
rect 150724 -27497 150780 -27441
rect 150804 -27497 150860 -27441
rect 150884 -27497 150940 -27441
rect 150964 -27497 151020 -27441
rect 151044 -27497 151100 -27441
rect 151124 -27497 151180 -27441
rect 151204 -27497 151260 -27441
rect 151284 -27497 151340 -27441
rect 151364 -27497 151420 -27441
rect 151444 -27497 151500 -27441
rect 151524 -27497 151580 -27441
rect 151604 -27497 151660 -27441
rect 151684 -27497 151740 -27441
rect 151764 -27497 151820 -27441
rect 151844 -27497 151900 -27441
rect 151924 -27497 151980 -27441
rect 152004 -27497 152060 -27441
rect 152084 -27497 152140 -27441
rect 152164 -27497 152220 -27441
rect 152244 -27497 152300 -27441
rect 152324 -27497 152380 -27441
rect 152404 -27497 152460 -27441
rect 152484 -27497 152540 -27441
rect 152564 -27497 152620 -27441
rect 152644 -27497 152700 -27441
rect 152724 -27497 152780 -27441
rect 152804 -27497 152860 -27441
rect 152884 -27497 152940 -27441
rect 152964 -27497 153020 -27441
rect 153044 -27497 153100 -27441
rect 153124 -27497 153180 -27441
rect 153204 -27497 153260 -27441
rect 153284 -27497 153340 -27441
rect 153364 -27497 153420 -27441
rect 153444 -27497 153500 -27441
rect 153524 -27497 153580 -27441
rect 153604 -27497 153660 -27441
rect 153684 -27497 153740 -27441
rect 153764 -27497 153820 -27441
rect 153844 -27497 153900 -27441
rect 153924 -27497 153980 -27441
rect 154004 -27497 154060 -27441
rect 154084 -27497 154140 -27441
rect 154164 -27497 154220 -27441
rect 154244 -27497 154300 -27441
rect 154324 -27497 154380 -27441
rect 154404 -27497 154460 -27441
rect 154484 -27497 154540 -27441
rect 154564 -27497 154620 -27441
rect 154644 -27497 154700 -27441
rect 154724 -27497 154780 -27441
rect 154804 -27497 154860 -27441
rect 154884 -27497 154940 -27441
rect 154964 -27497 155020 -27441
rect 155044 -27497 155100 -27441
rect 155124 -27497 155180 -27441
rect 155204 -27497 155260 -27441
rect 155284 -27497 155340 -27441
rect 155364 -27497 155420 -27441
rect 155444 -27497 155500 -27441
rect 155524 -27497 155580 -27441
rect 155604 -27497 155660 -27441
rect 155684 -27497 155740 -27441
rect 155764 -27497 155820 -27441
rect 155844 -27497 155900 -27441
rect 155924 -27497 155980 -27441
rect 156004 -27497 156060 -27441
rect 156084 -27497 156140 -27441
rect 156164 -27497 156220 -27441
rect 156244 -27497 156300 -27441
rect 156324 -27497 156380 -27441
rect 166967 -28140 167014 -28096
rect 167014 -28140 167023 -28096
rect 167047 -28140 167078 -28096
rect 167078 -28140 167090 -28096
rect 167090 -28140 167103 -28096
rect 167127 -28140 167142 -28096
rect 167142 -28140 167154 -28096
rect 167154 -28140 167183 -28096
rect 167207 -28140 167218 -28096
rect 167218 -28140 167263 -28096
rect 167287 -28140 167334 -28096
rect 167334 -28140 167343 -28096
rect 167367 -28140 167398 -28096
rect 167398 -28140 167410 -28096
rect 167410 -28140 167423 -28096
rect 167447 -28140 167462 -28096
rect 167462 -28140 167474 -28096
rect 167474 -28140 167503 -28096
rect 167527 -28140 167538 -28096
rect 167538 -28140 167583 -28096
rect 166967 -28152 167023 -28140
rect 167047 -28152 167103 -28140
rect 167127 -28152 167183 -28140
rect 167207 -28152 167263 -28140
rect 167287 -28152 167343 -28140
rect 167367 -28152 167423 -28140
rect 167447 -28152 167503 -28140
rect 167527 -28152 167583 -28140
rect 169494 -28177 169710 -27961
rect 146865 -31516 167401 -31380
<< metal3 >>
rect 146874 14156 156352 16000
rect 146874 1932 148571 14156
rect 154635 1932 156352 14156
rect 146874 -24694 156352 1932
rect 156671 -20628 160881 -20476
rect 156671 -20655 160198 -20628
rect 156671 -21591 156793 -20655
rect 158049 -21572 160198 -20655
rect 160742 -21572 160881 -20628
rect 158049 -21591 160881 -21572
rect 156671 -21689 160881 -21591
rect 160343 -23179 164348 -23106
rect 160343 -23323 160467 -23179
rect 164211 -23323 164348 -23179
rect 160343 -25029 164348 -23323
rect 160343 -25085 160442 -25029
rect 160498 -25085 160522 -25029
rect 160578 -25085 160602 -25029
rect 160658 -25085 160682 -25029
rect 160738 -25085 160762 -25029
rect 160818 -25085 160842 -25029
rect 160898 -25085 160922 -25029
rect 160978 -25085 161002 -25029
rect 161058 -25085 161082 -25029
rect 161138 -25085 161162 -25029
rect 161218 -25085 161242 -25029
rect 161298 -25085 161322 -25029
rect 161378 -25085 161402 -25029
rect 161458 -25085 161482 -25029
rect 161538 -25085 161562 -25029
rect 161618 -25085 161642 -25029
rect 161698 -25085 161722 -25029
rect 161778 -25085 161802 -25029
rect 161858 -25085 161882 -25029
rect 161938 -25085 161962 -25029
rect 162018 -25085 162042 -25029
rect 162098 -25085 162122 -25029
rect 162178 -25085 162202 -25029
rect 162258 -25085 162282 -25029
rect 162338 -25085 162362 -25029
rect 162418 -25085 162442 -25029
rect 162498 -25085 162522 -25029
rect 162578 -25085 162602 -25029
rect 162658 -25085 162682 -25029
rect 162738 -25085 162762 -25029
rect 162818 -25085 162842 -25029
rect 162898 -25085 162922 -25029
rect 162978 -25085 163002 -25029
rect 163058 -25085 163082 -25029
rect 163138 -25085 163162 -25029
rect 163218 -25085 163242 -25029
rect 163298 -25085 163322 -25029
rect 163378 -25085 163402 -25029
rect 163458 -25085 163482 -25029
rect 163538 -25085 163562 -25029
rect 163618 -25085 163642 -25029
rect 163698 -25085 163722 -25029
rect 163778 -25085 163802 -25029
rect 163858 -25085 163882 -25029
rect 163938 -25085 163962 -25029
rect 164018 -25085 164042 -25029
rect 164098 -25085 164122 -25029
rect 164178 -25085 164202 -25029
rect 164258 -25085 164348 -25029
rect 160343 -25164 164348 -25085
rect 146912 -27441 156428 -27432
rect 146912 -27497 146964 -27441
rect 147020 -27497 147044 -27441
rect 147100 -27497 147124 -27441
rect 147180 -27497 147204 -27441
rect 147260 -27497 147284 -27441
rect 147340 -27497 147364 -27441
rect 147420 -27497 147444 -27441
rect 147500 -27497 147524 -27441
rect 147580 -27497 147604 -27441
rect 147660 -27497 147684 -27441
rect 147740 -27497 147764 -27441
rect 147820 -27497 147844 -27441
rect 147900 -27497 147924 -27441
rect 147980 -27497 148004 -27441
rect 148060 -27497 148084 -27441
rect 148140 -27497 148164 -27441
rect 148220 -27497 148244 -27441
rect 148300 -27497 148324 -27441
rect 148380 -27497 148404 -27441
rect 148460 -27497 148484 -27441
rect 148540 -27497 148564 -27441
rect 148620 -27497 148644 -27441
rect 148700 -27497 148724 -27441
rect 148780 -27497 148804 -27441
rect 148860 -27497 148884 -27441
rect 148940 -27497 148964 -27441
rect 149020 -27497 149044 -27441
rect 149100 -27497 149124 -27441
rect 149180 -27497 149204 -27441
rect 149260 -27497 149284 -27441
rect 149340 -27497 149364 -27441
rect 149420 -27497 149444 -27441
rect 149500 -27497 149524 -27441
rect 149580 -27497 149604 -27441
rect 149660 -27497 149684 -27441
rect 149740 -27497 149764 -27441
rect 149820 -27497 149844 -27441
rect 149900 -27497 149924 -27441
rect 149980 -27497 150004 -27441
rect 150060 -27497 150084 -27441
rect 150140 -27497 150164 -27441
rect 150220 -27497 150244 -27441
rect 150300 -27497 150324 -27441
rect 150380 -27497 150404 -27441
rect 150460 -27497 150484 -27441
rect 150540 -27497 150564 -27441
rect 150620 -27497 150644 -27441
rect 150700 -27497 150724 -27441
rect 150780 -27497 150804 -27441
rect 150860 -27497 150884 -27441
rect 150940 -27497 150964 -27441
rect 151020 -27497 151044 -27441
rect 151100 -27497 151124 -27441
rect 151180 -27497 151204 -27441
rect 151260 -27497 151284 -27441
rect 151340 -27497 151364 -27441
rect 151420 -27497 151444 -27441
rect 151500 -27497 151524 -27441
rect 151580 -27497 151604 -27441
rect 151660 -27497 151684 -27441
rect 151740 -27497 151764 -27441
rect 151820 -27497 151844 -27441
rect 151900 -27497 151924 -27441
rect 151980 -27497 152004 -27441
rect 152060 -27497 152084 -27441
rect 152140 -27497 152164 -27441
rect 152220 -27497 152244 -27441
rect 152300 -27497 152324 -27441
rect 152380 -27497 152404 -27441
rect 152460 -27497 152484 -27441
rect 152540 -27497 152564 -27441
rect 152620 -27497 152644 -27441
rect 152700 -27497 152724 -27441
rect 152780 -27497 152804 -27441
rect 152860 -27497 152884 -27441
rect 152940 -27497 152964 -27441
rect 153020 -27497 153044 -27441
rect 153100 -27497 153124 -27441
rect 153180 -27497 153204 -27441
rect 153260 -27497 153284 -27441
rect 153340 -27497 153364 -27441
rect 153420 -27497 153444 -27441
rect 153500 -27497 153524 -27441
rect 153580 -27497 153604 -27441
rect 153660 -27497 153684 -27441
rect 153740 -27497 153764 -27441
rect 153820 -27497 153844 -27441
rect 153900 -27497 153924 -27441
rect 153980 -27497 154004 -27441
rect 154060 -27497 154084 -27441
rect 154140 -27497 154164 -27441
rect 154220 -27497 154244 -27441
rect 154300 -27497 154324 -27441
rect 154380 -27497 154404 -27441
rect 154460 -27497 154484 -27441
rect 154540 -27497 154564 -27441
rect 154620 -27497 154644 -27441
rect 154700 -27497 154724 -27441
rect 154780 -27497 154804 -27441
rect 154860 -27497 154884 -27441
rect 154940 -27497 154964 -27441
rect 155020 -27497 155044 -27441
rect 155100 -27497 155124 -27441
rect 155180 -27497 155204 -27441
rect 155260 -27497 155284 -27441
rect 155340 -27497 155364 -27441
rect 155420 -27497 155444 -27441
rect 155500 -27497 155524 -27441
rect 155580 -27497 155604 -27441
rect 155660 -27497 155684 -27441
rect 155740 -27497 155764 -27441
rect 155820 -27497 155844 -27441
rect 155900 -27497 155924 -27441
rect 155980 -27497 156004 -27441
rect 156060 -27497 156084 -27441
rect 156140 -27497 156164 -27441
rect 156220 -27497 156244 -27441
rect 156300 -27497 156324 -27441
rect 156380 -27497 156428 -27441
rect 146912 -28138 156428 -27497
rect 169409 -27961 170803 -27925
rect 166710 -28096 167694 -28012
rect 166710 -28152 166967 -28096
rect 167023 -28152 167047 -28096
rect 167103 -28152 167127 -28096
rect 167183 -28152 167207 -28096
rect 167263 -28152 167287 -28096
rect 167343 -28152 167367 -28096
rect 167423 -28152 167447 -28096
rect 167503 -28152 167527 -28096
rect 167583 -28152 167694 -28096
rect 166710 -28165 167694 -28152
rect 166772 -28168 167694 -28165
rect 166804 -28208 167656 -28168
rect 169409 -28177 169494 -27961
rect 169710 -27962 170803 -27961
rect 169710 -28177 170460 -27962
rect 169409 -28186 170460 -28177
rect 170764 -28186 170803 -27962
rect 169409 -28213 170803 -28186
rect 146772 -31334 168651 -31277
rect 146772 -31380 168184 -31334
rect 146772 -31516 146865 -31380
rect 167401 -31516 168184 -31380
rect 146772 -31558 168184 -31516
rect 168568 -31558 168651 -31334
rect 146772 -31615 168651 -31558
<< via3 >>
rect 148571 1932 154635 14156
rect 160198 -21572 160742 -20628
rect 160467 -23323 164211 -23179
rect 170460 -28186 170764 -27962
rect 168184 -31558 168568 -31334
<< metal4 >>
rect 146874 14823 156352 16000
rect 146874 1147 147936 14823
rect 155212 1147 156352 14823
rect 146874 0 156352 1147
rect 160074 -20628 164284 -20476
rect 160074 -21572 160198 -20628
rect 160742 -20659 164284 -20628
rect 160742 -21535 163188 -20659
rect 163744 -21535 164284 -20659
rect 160742 -21572 164284 -21535
rect 160074 -21689 164284 -21572
rect 160343 -22665 165003 -22504
rect 160343 -22901 164648 -22665
rect 164884 -22901 165003 -22665
rect 160343 -22985 165003 -22901
rect 160343 -23179 164648 -22985
rect 160343 -23323 160467 -23179
rect 164211 -23221 164648 -23179
rect 164884 -23221 165003 -22985
rect 164211 -23323 165003 -23221
rect 160343 -23370 165003 -23323
rect 170438 -27962 171909 -27925
rect 170438 -28186 170460 -27962
rect 170764 -27964 171909 -27962
rect 170764 -28186 171582 -27964
rect 170438 -28200 171582 -28186
rect 171818 -28200 171909 -27964
rect 170438 -28213 171909 -28200
rect 168109 -30883 170325 -30630
rect 168109 -31119 169861 -30883
rect 170097 -31119 170325 -30883
rect 168109 -31203 170325 -31119
rect 168109 -31334 169861 -31203
rect 168109 -31558 168184 -31334
rect 168568 -31439 169861 -31334
rect 170097 -31439 170325 -31203
rect 168568 -31558 170325 -31439
rect 168109 -31651 170325 -31558
<< via4 >>
rect 147936 14156 155212 14823
rect 147936 1932 148571 14156
rect 148571 1932 154635 14156
rect 154635 1932 155212 14156
rect 147936 1147 155212 1932
rect 163188 -21535 163744 -20659
rect 164648 -22901 164884 -22665
rect 164648 -23221 164884 -22985
rect 171582 -28200 171818 -27964
rect 169861 -31119 170097 -30883
rect 169861 -31439 170097 -31203
<< metal5 >>
rect 146874 14823 156352 16000
rect 146874 1147 147936 14823
rect 155212 1147 156352 14823
rect 146874 0 156352 1147
rect 163107 -20659 167317 -20476
rect 163107 -21535 163188 -20659
rect 163744 -21535 167317 -20659
rect 163107 -21689 167317 -21535
rect 164597 -22665 169257 -22504
rect 164597 -22901 164648 -22665
rect 164884 -22901 169257 -22665
rect 164597 -22985 169257 -22901
rect 164597 -23221 164648 -22985
rect 164884 -23221 169257 -22985
rect 164597 -23370 169257 -23221
rect 171445 -27964 172056 -27810
rect 171445 -28200 171582 -27964
rect 171818 -28200 172056 -27964
rect 171445 -28303 172056 -28200
rect 169750 -30883 171581 -30396
rect 169750 -31119 169861 -30883
rect 170097 -31119 171581 -30883
rect 169750 -31203 171581 -31119
rect 169750 -31439 169861 -31203
rect 170097 -31439 171581 -31203
rect 169750 -31847 171581 -31439
use sky130_fd_pr__res_generic_po_u1tz6h  sky130_fd_pr__res_generic_po_u1tz6h_0
timestamp 1611881054
transform 1 0 162342 0 1 -26306
box -2166 -404 2166 404
use sky130_fd_pr__res_high_po_0p35_i8je6j  sky130_fd_pr__res_high_po_0p35_i8je6j_0
timestamp 1611881054
transform 1 0 167251 0 1 -26054
box -1596 -1562 1596 1562
use transistor_1m  transistor_1m_0
timestamp 1611881054
transform 1 0 128835 0 1 -31687
box 28923 745 38986 3606
use transistor_1m  transistor_1m_1
timestamp 1611881054
transform 1 0 117795 0 1 -31685
box 28923 745 38986 3606
use transistor_1m  transistor_1m_2
timestamp 1611881054
transform 1 0 117759 0 1 -28251
box 28923 745 38986 3606
use INDUCTOR_L  INDUCTOR_L_0
timestamp 1611881054
transform 1 0 432600 0 1 171000
box -432600 -171000 -79800 178200
<< labels >>
rlabel metal3 s 147547 -13778 155259 -3811 4 out
rlabel metal5 s 166668 -21526 167008 -20656 4 Vgate
port 1 nsew
rlabel metal5 s 171926 -28261 172027 -27853 4 Isource
port 2 nsew
rlabel metal5 s 168834 -23282 169169 -22611 4 Rnode
port 3 nsew
rlabel metal5 s 171123 -31584 171405 -30698 4 vss
port 4 nsew
<< end >>
