magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -227 194 227 228
rect -227 -194 -193 194
rect 193 -194 227 194
rect -227 -228 227 -194
<< nmos >>
rect -63 -54 -33 54
rect 33 -54 63 54
<< ndiff >>
rect -125 17 -63 54
rect -125 -17 -113 17
rect -79 -17 -63 17
rect -125 -54 -63 -17
rect -33 17 33 54
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -54 33 -17
rect 63 17 125 54
rect 63 -17 79 17
rect 113 -17 125 17
rect 63 -54 125 -17
<< ndiffc >>
rect -113 -17 -79 17
rect -17 -17 17 17
rect 79 -17 113 17
<< psubdiff >>
rect -227 194 -119 228
rect -85 194 -51 228
rect -17 194 17 228
rect 51 194 85 228
rect 119 194 227 228
rect -227 119 -193 194
rect -227 51 -193 85
rect 193 119 227 194
rect -227 -17 -193 17
rect -227 -85 -193 -51
rect 193 51 227 85
rect 193 -17 227 17
rect -227 -194 -193 -119
rect 193 -85 227 -51
rect 193 -194 227 -119
rect -227 -228 -119 -194
rect -85 -228 -51 -194
rect -17 -228 17 -194
rect 51 -228 85 -194
rect 119 -228 227 -194
<< psubdiffcont >>
rect -119 194 -85 228
rect -51 194 -17 228
rect 17 194 51 228
rect 85 194 119 228
rect -227 85 -193 119
rect 193 85 227 119
rect -227 17 -193 51
rect -227 -51 -193 -17
rect 193 17 227 51
rect 193 -51 227 -17
rect -227 -119 -193 -85
rect 193 -119 227 -85
rect -119 -228 -85 -194
rect -51 -228 -17 -194
rect 17 -228 51 -194
rect 85 -228 119 -194
<< poly >>
rect 15 126 81 142
rect 15 92 31 126
rect 65 92 81 126
rect -63 54 -33 80
rect 15 76 81 92
rect 33 54 63 76
rect -63 -76 -33 -54
rect -81 -92 -15 -76
rect 33 -80 63 -54
rect -81 -126 -65 -92
rect -31 -126 -15 -92
rect -81 -142 -15 -126
<< polycont >>
rect 31 92 65 126
rect -65 -126 -31 -92
<< locali >>
rect -227 194 -119 228
rect -85 194 -51 228
rect -17 194 17 228
rect 51 194 85 228
rect 119 194 227 228
rect -227 119 -193 194
rect 15 92 31 126
rect 65 92 81 126
rect 193 119 227 194
rect -227 51 -193 85
rect -227 -17 -193 17
rect -227 -85 -193 -51
rect -113 17 -79 58
rect -113 -58 -79 -17
rect -17 17 17 58
rect -17 -58 17 -17
rect 79 17 113 58
rect 79 -58 113 -17
rect 193 51 227 85
rect 193 -17 227 17
rect 193 -85 227 -51
rect -227 -194 -193 -119
rect -81 -126 -65 -92
rect -31 -126 -15 -92
rect 193 -194 227 -119
rect -227 -228 -119 -194
rect -85 -228 -51 -194
rect -17 -228 17 -194
rect 51 -228 85 -194
rect 119 -228 227 -194
<< viali >>
rect -113 -17 -79 17
rect -17 -17 17 17
rect 79 -17 113 17
<< metal1 >>
rect -119 17 -73 54
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -54 -73 -17
rect -23 17 23 54
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -54 23 -17
rect 73 17 119 54
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -54 119 -17
<< properties >>
string FIXED_BBOX -210 -211 210 211
<< end >>
