magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< error_p >>
rect -29 1072 29 1078
rect -29 1038 -17 1072
rect -29 1032 29 1038
rect -29 -1038 29 -1032
rect -29 -1072 -17 -1038
rect -29 -1078 29 -1072
<< pwell >>
rect -175 1140 175 1174
rect -175 -1140 -141 1140
rect 141 -1140 175 1140
rect -175 -1174 175 -1140
<< nmos >>
rect -15 -1000 15 1000
<< ndiff >>
rect -73 969 -15 1000
rect -73 935 -61 969
rect -27 935 -15 969
rect -73 901 -15 935
rect -73 867 -61 901
rect -27 867 -15 901
rect -73 833 -15 867
rect -73 799 -61 833
rect -27 799 -15 833
rect -73 765 -15 799
rect -73 731 -61 765
rect -27 731 -15 765
rect -73 697 -15 731
rect -73 663 -61 697
rect -27 663 -15 697
rect -73 629 -15 663
rect -73 595 -61 629
rect -27 595 -15 629
rect -73 561 -15 595
rect -73 527 -61 561
rect -27 527 -15 561
rect -73 493 -15 527
rect -73 459 -61 493
rect -27 459 -15 493
rect -73 425 -15 459
rect -73 391 -61 425
rect -27 391 -15 425
rect -73 357 -15 391
rect -73 323 -61 357
rect -27 323 -15 357
rect -73 289 -15 323
rect -73 255 -61 289
rect -27 255 -15 289
rect -73 221 -15 255
rect -73 187 -61 221
rect -27 187 -15 221
rect -73 153 -15 187
rect -73 119 -61 153
rect -27 119 -15 153
rect -73 85 -15 119
rect -73 51 -61 85
rect -27 51 -15 85
rect -73 17 -15 51
rect -73 -17 -61 17
rect -27 -17 -15 17
rect -73 -51 -15 -17
rect -73 -85 -61 -51
rect -27 -85 -15 -51
rect -73 -119 -15 -85
rect -73 -153 -61 -119
rect -27 -153 -15 -119
rect -73 -187 -15 -153
rect -73 -221 -61 -187
rect -27 -221 -15 -187
rect -73 -255 -15 -221
rect -73 -289 -61 -255
rect -27 -289 -15 -255
rect -73 -323 -15 -289
rect -73 -357 -61 -323
rect -27 -357 -15 -323
rect -73 -391 -15 -357
rect -73 -425 -61 -391
rect -27 -425 -15 -391
rect -73 -459 -15 -425
rect -73 -493 -61 -459
rect -27 -493 -15 -459
rect -73 -527 -15 -493
rect -73 -561 -61 -527
rect -27 -561 -15 -527
rect -73 -595 -15 -561
rect -73 -629 -61 -595
rect -27 -629 -15 -595
rect -73 -663 -15 -629
rect -73 -697 -61 -663
rect -27 -697 -15 -663
rect -73 -731 -15 -697
rect -73 -765 -61 -731
rect -27 -765 -15 -731
rect -73 -799 -15 -765
rect -73 -833 -61 -799
rect -27 -833 -15 -799
rect -73 -867 -15 -833
rect -73 -901 -61 -867
rect -27 -901 -15 -867
rect -73 -935 -15 -901
rect -73 -969 -61 -935
rect -27 -969 -15 -935
rect -73 -1000 -15 -969
rect 15 969 73 1000
rect 15 935 27 969
rect 61 935 73 969
rect 15 901 73 935
rect 15 867 27 901
rect 61 867 73 901
rect 15 833 73 867
rect 15 799 27 833
rect 61 799 73 833
rect 15 765 73 799
rect 15 731 27 765
rect 61 731 73 765
rect 15 697 73 731
rect 15 663 27 697
rect 61 663 73 697
rect 15 629 73 663
rect 15 595 27 629
rect 61 595 73 629
rect 15 561 73 595
rect 15 527 27 561
rect 61 527 73 561
rect 15 493 73 527
rect 15 459 27 493
rect 61 459 73 493
rect 15 425 73 459
rect 15 391 27 425
rect 61 391 73 425
rect 15 357 73 391
rect 15 323 27 357
rect 61 323 73 357
rect 15 289 73 323
rect 15 255 27 289
rect 61 255 73 289
rect 15 221 73 255
rect 15 187 27 221
rect 61 187 73 221
rect 15 153 73 187
rect 15 119 27 153
rect 61 119 73 153
rect 15 85 73 119
rect 15 51 27 85
rect 61 51 73 85
rect 15 17 73 51
rect 15 -17 27 17
rect 61 -17 73 17
rect 15 -51 73 -17
rect 15 -85 27 -51
rect 61 -85 73 -51
rect 15 -119 73 -85
rect 15 -153 27 -119
rect 61 -153 73 -119
rect 15 -187 73 -153
rect 15 -221 27 -187
rect 61 -221 73 -187
rect 15 -255 73 -221
rect 15 -289 27 -255
rect 61 -289 73 -255
rect 15 -323 73 -289
rect 15 -357 27 -323
rect 61 -357 73 -323
rect 15 -391 73 -357
rect 15 -425 27 -391
rect 61 -425 73 -391
rect 15 -459 73 -425
rect 15 -493 27 -459
rect 61 -493 73 -459
rect 15 -527 73 -493
rect 15 -561 27 -527
rect 61 -561 73 -527
rect 15 -595 73 -561
rect 15 -629 27 -595
rect 61 -629 73 -595
rect 15 -663 73 -629
rect 15 -697 27 -663
rect 61 -697 73 -663
rect 15 -731 73 -697
rect 15 -765 27 -731
rect 61 -765 73 -731
rect 15 -799 73 -765
rect 15 -833 27 -799
rect 61 -833 73 -799
rect 15 -867 73 -833
rect 15 -901 27 -867
rect 61 -901 73 -867
rect 15 -935 73 -901
rect 15 -969 27 -935
rect 61 -969 73 -935
rect 15 -1000 73 -969
<< ndiffc >>
rect -61 935 -27 969
rect -61 867 -27 901
rect -61 799 -27 833
rect -61 731 -27 765
rect -61 663 -27 697
rect -61 595 -27 629
rect -61 527 -27 561
rect -61 459 -27 493
rect -61 391 -27 425
rect -61 323 -27 357
rect -61 255 -27 289
rect -61 187 -27 221
rect -61 119 -27 153
rect -61 51 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -51
rect -61 -153 -27 -119
rect -61 -221 -27 -187
rect -61 -289 -27 -255
rect -61 -357 -27 -323
rect -61 -425 -27 -391
rect -61 -493 -27 -459
rect -61 -561 -27 -527
rect -61 -629 -27 -595
rect -61 -697 -27 -663
rect -61 -765 -27 -731
rect -61 -833 -27 -799
rect -61 -901 -27 -867
rect -61 -969 -27 -935
rect 27 935 61 969
rect 27 867 61 901
rect 27 799 61 833
rect 27 731 61 765
rect 27 663 61 697
rect 27 595 61 629
rect 27 527 61 561
rect 27 459 61 493
rect 27 391 61 425
rect 27 323 61 357
rect 27 255 61 289
rect 27 187 61 221
rect 27 119 61 153
rect 27 51 61 85
rect 27 -17 61 17
rect 27 -85 61 -51
rect 27 -153 61 -119
rect 27 -221 61 -187
rect 27 -289 61 -255
rect 27 -357 61 -323
rect 27 -425 61 -391
rect 27 -493 61 -459
rect 27 -561 61 -527
rect 27 -629 61 -595
rect 27 -697 61 -663
rect 27 -765 61 -731
rect 27 -833 61 -799
rect 27 -901 61 -867
rect 27 -969 61 -935
<< psubdiff >>
rect -175 1140 -51 1174
rect -17 1140 17 1174
rect 51 1140 175 1174
rect -175 1071 -141 1140
rect -175 1003 -141 1037
rect 141 1071 175 1140
rect 141 1003 175 1037
rect -175 935 -141 969
rect -175 867 -141 901
rect -175 799 -141 833
rect -175 731 -141 765
rect -175 663 -141 697
rect -175 595 -141 629
rect -175 527 -141 561
rect -175 459 -141 493
rect -175 391 -141 425
rect -175 323 -141 357
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -175 -357 -141 -323
rect -175 -425 -141 -391
rect -175 -493 -141 -459
rect -175 -561 -141 -527
rect -175 -629 -141 -595
rect -175 -697 -141 -663
rect -175 -765 -141 -731
rect -175 -833 -141 -799
rect -175 -901 -141 -867
rect -175 -969 -141 -935
rect 141 935 175 969
rect 141 867 175 901
rect 141 799 175 833
rect 141 731 175 765
rect 141 663 175 697
rect 141 595 175 629
rect 141 527 175 561
rect 141 459 175 493
rect 141 391 175 425
rect 141 323 175 357
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect 141 -357 175 -323
rect 141 -425 175 -391
rect 141 -493 175 -459
rect 141 -561 175 -527
rect 141 -629 175 -595
rect 141 -697 175 -663
rect 141 -765 175 -731
rect 141 -833 175 -799
rect 141 -901 175 -867
rect 141 -969 175 -935
rect -175 -1037 -141 -1003
rect -175 -1140 -141 -1071
rect 141 -1037 175 -1003
rect 141 -1140 175 -1071
rect -175 -1174 -51 -1140
rect -17 -1174 17 -1140
rect 51 -1174 175 -1140
<< psubdiffcont >>
rect -51 1140 -17 1174
rect 17 1140 51 1174
rect -175 1037 -141 1071
rect 141 1037 175 1071
rect -175 969 -141 1003
rect -175 901 -141 935
rect -175 833 -141 867
rect -175 765 -141 799
rect -175 697 -141 731
rect -175 629 -141 663
rect -175 561 -141 595
rect -175 493 -141 527
rect -175 425 -141 459
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -459 -141 -425
rect -175 -527 -141 -493
rect -175 -595 -141 -561
rect -175 -663 -141 -629
rect -175 -731 -141 -697
rect -175 -799 -141 -765
rect -175 -867 -141 -833
rect -175 -935 -141 -901
rect -175 -1003 -141 -969
rect 141 969 175 1003
rect 141 901 175 935
rect 141 833 175 867
rect 141 765 175 799
rect 141 697 175 731
rect 141 629 175 663
rect 141 561 175 595
rect 141 493 175 527
rect 141 425 175 459
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -459 175 -425
rect 141 -527 175 -493
rect 141 -595 175 -561
rect 141 -663 175 -629
rect 141 -731 175 -697
rect 141 -799 175 -765
rect 141 -867 175 -833
rect 141 -935 175 -901
rect 141 -1003 175 -969
rect -175 -1071 -141 -1037
rect 141 -1071 175 -1037
rect -51 -1174 -17 -1140
rect 17 -1174 51 -1140
<< poly >>
rect -33 1072 33 1088
rect -33 1038 -17 1072
rect 17 1038 33 1072
rect -33 1022 33 1038
rect -15 1000 15 1022
rect -15 -1022 15 -1000
rect -33 -1038 33 -1022
rect -33 -1072 -17 -1038
rect 17 -1072 33 -1038
rect -33 -1088 33 -1072
<< polycont >>
rect -17 1038 17 1072
rect -17 -1072 17 -1038
<< locali >>
rect -175 1140 -51 1174
rect -17 1140 17 1174
rect 51 1140 175 1174
rect -175 1071 -141 1140
rect -33 1038 -17 1072
rect 17 1038 33 1072
rect 141 1071 175 1140
rect -175 1003 -141 1037
rect -175 935 -141 969
rect -175 867 -141 901
rect -175 799 -141 833
rect -175 731 -141 765
rect -175 663 -141 697
rect -175 595 -141 629
rect -175 527 -141 561
rect -175 459 -141 493
rect -175 391 -141 425
rect -175 323 -141 357
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -175 -357 -141 -323
rect -175 -425 -141 -391
rect -175 -493 -141 -459
rect -175 -561 -141 -527
rect -175 -629 -141 -595
rect -175 -697 -141 -663
rect -175 -765 -141 -731
rect -175 -833 -141 -799
rect -175 -901 -141 -867
rect -175 -969 -141 -935
rect -175 -1037 -141 -1003
rect -61 969 -27 1004
rect -61 901 -27 919
rect -61 833 -27 847
rect -61 765 -27 775
rect -61 697 -27 703
rect -61 629 -27 631
rect -61 593 -27 595
rect -61 521 -27 527
rect -61 449 -27 459
rect -61 377 -27 391
rect -61 305 -27 323
rect -61 233 -27 255
rect -61 161 -27 187
rect -61 89 -27 119
rect -61 17 -27 51
rect -61 -51 -27 -17
rect -61 -119 -27 -89
rect -61 -187 -27 -161
rect -61 -255 -27 -233
rect -61 -323 -27 -305
rect -61 -391 -27 -377
rect -61 -459 -27 -449
rect -61 -527 -27 -521
rect -61 -595 -27 -593
rect -61 -631 -27 -629
rect -61 -703 -27 -697
rect -61 -775 -27 -765
rect -61 -847 -27 -833
rect -61 -919 -27 -901
rect -61 -1004 -27 -969
rect 27 969 61 1004
rect 27 901 61 919
rect 27 833 61 847
rect 27 765 61 775
rect 27 697 61 703
rect 27 629 61 631
rect 27 593 61 595
rect 27 521 61 527
rect 27 449 61 459
rect 27 377 61 391
rect 27 305 61 323
rect 27 233 61 255
rect 27 161 61 187
rect 27 89 61 119
rect 27 17 61 51
rect 27 -51 61 -17
rect 27 -119 61 -89
rect 27 -187 61 -161
rect 27 -255 61 -233
rect 27 -323 61 -305
rect 27 -391 61 -377
rect 27 -459 61 -449
rect 27 -527 61 -521
rect 27 -595 61 -593
rect 27 -631 61 -629
rect 27 -703 61 -697
rect 27 -775 61 -765
rect 27 -847 61 -833
rect 27 -919 61 -901
rect 27 -1004 61 -969
rect 141 1003 175 1037
rect 141 935 175 969
rect 141 867 175 901
rect 141 799 175 833
rect 141 731 175 765
rect 141 663 175 697
rect 141 595 175 629
rect 141 527 175 561
rect 141 459 175 493
rect 141 391 175 425
rect 141 323 175 357
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect 141 -357 175 -323
rect 141 -425 175 -391
rect 141 -493 175 -459
rect 141 -561 175 -527
rect 141 -629 175 -595
rect 141 -697 175 -663
rect 141 -765 175 -731
rect 141 -833 175 -799
rect 141 -901 175 -867
rect 141 -969 175 -935
rect 141 -1037 175 -1003
rect -175 -1140 -141 -1071
rect -33 -1072 -17 -1038
rect 17 -1072 33 -1038
rect 141 -1140 175 -1071
rect -175 -1174 -51 -1140
rect -17 -1174 17 -1140
rect 51 -1174 175 -1140
<< viali >>
rect -17 1038 17 1072
rect -61 935 -27 953
rect -61 919 -27 935
rect -61 867 -27 881
rect -61 847 -27 867
rect -61 799 -27 809
rect -61 775 -27 799
rect -61 731 -27 737
rect -61 703 -27 731
rect -61 663 -27 665
rect -61 631 -27 663
rect -61 561 -27 593
rect -61 559 -27 561
rect -61 493 -27 521
rect -61 487 -27 493
rect -61 425 -27 449
rect -61 415 -27 425
rect -61 357 -27 377
rect -61 343 -27 357
rect -61 289 -27 305
rect -61 271 -27 289
rect -61 221 -27 233
rect -61 199 -27 221
rect -61 153 -27 161
rect -61 127 -27 153
rect -61 85 -27 89
rect -61 55 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -55
rect -61 -89 -27 -85
rect -61 -153 -27 -127
rect -61 -161 -27 -153
rect -61 -221 -27 -199
rect -61 -233 -27 -221
rect -61 -289 -27 -271
rect -61 -305 -27 -289
rect -61 -357 -27 -343
rect -61 -377 -27 -357
rect -61 -425 -27 -415
rect -61 -449 -27 -425
rect -61 -493 -27 -487
rect -61 -521 -27 -493
rect -61 -561 -27 -559
rect -61 -593 -27 -561
rect -61 -663 -27 -631
rect -61 -665 -27 -663
rect -61 -731 -27 -703
rect -61 -737 -27 -731
rect -61 -799 -27 -775
rect -61 -809 -27 -799
rect -61 -867 -27 -847
rect -61 -881 -27 -867
rect -61 -935 -27 -919
rect -61 -953 -27 -935
rect 27 935 61 953
rect 27 919 61 935
rect 27 867 61 881
rect 27 847 61 867
rect 27 799 61 809
rect 27 775 61 799
rect 27 731 61 737
rect 27 703 61 731
rect 27 663 61 665
rect 27 631 61 663
rect 27 561 61 593
rect 27 559 61 561
rect 27 493 61 521
rect 27 487 61 493
rect 27 425 61 449
rect 27 415 61 425
rect 27 357 61 377
rect 27 343 61 357
rect 27 289 61 305
rect 27 271 61 289
rect 27 221 61 233
rect 27 199 61 221
rect 27 153 61 161
rect 27 127 61 153
rect 27 85 61 89
rect 27 55 61 85
rect 27 -17 61 17
rect 27 -85 61 -55
rect 27 -89 61 -85
rect 27 -153 61 -127
rect 27 -161 61 -153
rect 27 -221 61 -199
rect 27 -233 61 -221
rect 27 -289 61 -271
rect 27 -305 61 -289
rect 27 -357 61 -343
rect 27 -377 61 -357
rect 27 -425 61 -415
rect 27 -449 61 -425
rect 27 -493 61 -487
rect 27 -521 61 -493
rect 27 -561 61 -559
rect 27 -593 61 -561
rect 27 -663 61 -631
rect 27 -665 61 -663
rect 27 -731 61 -703
rect 27 -737 61 -731
rect 27 -799 61 -775
rect 27 -809 61 -799
rect 27 -867 61 -847
rect 27 -881 61 -867
rect 27 -935 61 -919
rect 27 -953 61 -935
rect -17 -1072 17 -1038
<< metal1 >>
rect -29 1072 29 1078
rect -29 1038 -17 1072
rect 17 1038 29 1072
rect -29 1032 29 1038
rect -67 953 -21 1000
rect -67 919 -61 953
rect -27 919 -21 953
rect -67 881 -21 919
rect -67 847 -61 881
rect -27 847 -21 881
rect -67 809 -21 847
rect -67 775 -61 809
rect -27 775 -21 809
rect -67 737 -21 775
rect -67 703 -61 737
rect -27 703 -21 737
rect -67 665 -21 703
rect -67 631 -61 665
rect -27 631 -21 665
rect -67 593 -21 631
rect -67 559 -61 593
rect -27 559 -21 593
rect -67 521 -21 559
rect -67 487 -61 521
rect -27 487 -21 521
rect -67 449 -21 487
rect -67 415 -61 449
rect -27 415 -21 449
rect -67 377 -21 415
rect -67 343 -61 377
rect -27 343 -21 377
rect -67 305 -21 343
rect -67 271 -61 305
rect -27 271 -21 305
rect -67 233 -21 271
rect -67 199 -61 233
rect -27 199 -21 233
rect -67 161 -21 199
rect -67 127 -61 161
rect -27 127 -21 161
rect -67 89 -21 127
rect -67 55 -61 89
rect -27 55 -21 89
rect -67 17 -21 55
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -55 -21 -17
rect -67 -89 -61 -55
rect -27 -89 -21 -55
rect -67 -127 -21 -89
rect -67 -161 -61 -127
rect -27 -161 -21 -127
rect -67 -199 -21 -161
rect -67 -233 -61 -199
rect -27 -233 -21 -199
rect -67 -271 -21 -233
rect -67 -305 -61 -271
rect -27 -305 -21 -271
rect -67 -343 -21 -305
rect -67 -377 -61 -343
rect -27 -377 -21 -343
rect -67 -415 -21 -377
rect -67 -449 -61 -415
rect -27 -449 -21 -415
rect -67 -487 -21 -449
rect -67 -521 -61 -487
rect -27 -521 -21 -487
rect -67 -559 -21 -521
rect -67 -593 -61 -559
rect -27 -593 -21 -559
rect -67 -631 -21 -593
rect -67 -665 -61 -631
rect -27 -665 -21 -631
rect -67 -703 -21 -665
rect -67 -737 -61 -703
rect -27 -737 -21 -703
rect -67 -775 -21 -737
rect -67 -809 -61 -775
rect -27 -809 -21 -775
rect -67 -847 -21 -809
rect -67 -881 -61 -847
rect -27 -881 -21 -847
rect -67 -919 -21 -881
rect -67 -953 -61 -919
rect -27 -953 -21 -919
rect -67 -1000 -21 -953
rect 21 953 67 1000
rect 21 919 27 953
rect 61 919 67 953
rect 21 881 67 919
rect 21 847 27 881
rect 61 847 67 881
rect 21 809 67 847
rect 21 775 27 809
rect 61 775 67 809
rect 21 737 67 775
rect 21 703 27 737
rect 61 703 67 737
rect 21 665 67 703
rect 21 631 27 665
rect 61 631 67 665
rect 21 593 67 631
rect 21 559 27 593
rect 61 559 67 593
rect 21 521 67 559
rect 21 487 27 521
rect 61 487 67 521
rect 21 449 67 487
rect 21 415 27 449
rect 61 415 67 449
rect 21 377 67 415
rect 21 343 27 377
rect 61 343 67 377
rect 21 305 67 343
rect 21 271 27 305
rect 61 271 67 305
rect 21 233 67 271
rect 21 199 27 233
rect 61 199 67 233
rect 21 161 67 199
rect 21 127 27 161
rect 61 127 67 161
rect 21 89 67 127
rect 21 55 27 89
rect 61 55 67 89
rect 21 17 67 55
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -55 67 -17
rect 21 -89 27 -55
rect 61 -89 67 -55
rect 21 -127 67 -89
rect 21 -161 27 -127
rect 61 -161 67 -127
rect 21 -199 67 -161
rect 21 -233 27 -199
rect 61 -233 67 -199
rect 21 -271 67 -233
rect 21 -305 27 -271
rect 61 -305 67 -271
rect 21 -343 67 -305
rect 21 -377 27 -343
rect 61 -377 67 -343
rect 21 -415 67 -377
rect 21 -449 27 -415
rect 61 -449 67 -415
rect 21 -487 67 -449
rect 21 -521 27 -487
rect 61 -521 67 -487
rect 21 -559 67 -521
rect 21 -593 27 -559
rect 61 -593 67 -559
rect 21 -631 67 -593
rect 21 -665 27 -631
rect 61 -665 67 -631
rect 21 -703 67 -665
rect 21 -737 27 -703
rect 61 -737 67 -703
rect 21 -775 67 -737
rect 21 -809 27 -775
rect 61 -809 67 -775
rect 21 -847 67 -809
rect 21 -881 27 -847
rect 61 -881 67 -847
rect 21 -919 67 -881
rect 21 -953 27 -919
rect 61 -953 67 -919
rect 21 -1000 67 -953
rect -29 -1038 29 -1032
rect -29 -1072 -17 -1038
rect 17 -1072 29 -1038
rect -29 -1078 29 -1072
<< properties >>
string FIXED_BBOX -158 -1157 158 1157
<< end >>
