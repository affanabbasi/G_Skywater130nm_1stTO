magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -801 728 801 762
rect -801 -728 -767 728
rect 767 -728 801 728
rect -801 -762 801 -728
<< psubdiff >>
rect -801 728 -697 762
rect -663 728 -629 762
rect -595 728 -561 762
rect -527 728 -493 762
rect -459 728 -425 762
rect -391 728 -357 762
rect -323 728 -289 762
rect -255 728 -221 762
rect -187 728 -153 762
rect -119 728 -85 762
rect -51 728 -17 762
rect 17 728 51 762
rect 85 728 119 762
rect 153 728 187 762
rect 221 728 255 762
rect 289 728 323 762
rect 357 728 391 762
rect 425 728 459 762
rect 493 728 527 762
rect 561 728 595 762
rect 629 728 663 762
rect 697 728 801 762
rect -801 663 -767 728
rect 767 663 801 728
rect -801 595 -767 629
rect -801 527 -767 561
rect -801 459 -767 493
rect -801 391 -767 425
rect -801 323 -767 357
rect -801 255 -767 289
rect -801 187 -767 221
rect -801 119 -767 153
rect -801 51 -767 85
rect -801 -17 -767 17
rect -801 -85 -767 -51
rect -801 -153 -767 -119
rect -801 -221 -767 -187
rect -801 -289 -767 -255
rect -801 -357 -767 -323
rect -801 -425 -767 -391
rect -801 -493 -767 -459
rect -801 -561 -767 -527
rect -801 -629 -767 -595
rect 767 595 801 629
rect 767 527 801 561
rect 767 459 801 493
rect 767 391 801 425
rect 767 323 801 357
rect 767 255 801 289
rect 767 187 801 221
rect 767 119 801 153
rect 767 51 801 85
rect 767 -17 801 17
rect 767 -85 801 -51
rect 767 -153 801 -119
rect 767 -221 801 -187
rect 767 -289 801 -255
rect 767 -357 801 -323
rect 767 -425 801 -391
rect 767 -493 801 -459
rect 767 -561 801 -527
rect 767 -629 801 -595
rect -801 -728 -767 -663
rect 767 -728 801 -663
rect -801 -762 -697 -728
rect -663 -762 -629 -728
rect -595 -762 -561 -728
rect -527 -762 -493 -728
rect -459 -762 -425 -728
rect -391 -762 -357 -728
rect -323 -762 -289 -728
rect -255 -762 -221 -728
rect -187 -762 -153 -728
rect -119 -762 -85 -728
rect -51 -762 -17 -728
rect 17 -762 51 -728
rect 85 -762 119 -728
rect 153 -762 187 -728
rect 221 -762 255 -728
rect 289 -762 323 -728
rect 357 -762 391 -728
rect 425 -762 459 -728
rect 493 -762 527 -728
rect 561 -762 595 -728
rect 629 -762 663 -728
rect 697 -762 801 -728
<< psubdiffcont >>
rect -697 728 -663 762
rect -629 728 -595 762
rect -561 728 -527 762
rect -493 728 -459 762
rect -425 728 -391 762
rect -357 728 -323 762
rect -289 728 -255 762
rect -221 728 -187 762
rect -153 728 -119 762
rect -85 728 -51 762
rect -17 728 17 762
rect 51 728 85 762
rect 119 728 153 762
rect 187 728 221 762
rect 255 728 289 762
rect 323 728 357 762
rect 391 728 425 762
rect 459 728 493 762
rect 527 728 561 762
rect 595 728 629 762
rect 663 728 697 762
rect -801 629 -767 663
rect -801 561 -767 595
rect -801 493 -767 527
rect -801 425 -767 459
rect -801 357 -767 391
rect -801 289 -767 323
rect -801 221 -767 255
rect -801 153 -767 187
rect -801 85 -767 119
rect -801 17 -767 51
rect -801 -51 -767 -17
rect -801 -119 -767 -85
rect -801 -187 -767 -153
rect -801 -255 -767 -221
rect -801 -323 -767 -289
rect -801 -391 -767 -357
rect -801 -459 -767 -425
rect -801 -527 -767 -493
rect -801 -595 -767 -561
rect -801 -663 -767 -629
rect 767 629 801 663
rect 767 561 801 595
rect 767 493 801 527
rect 767 425 801 459
rect 767 357 801 391
rect 767 289 801 323
rect 767 221 801 255
rect 767 153 801 187
rect 767 85 801 119
rect 767 17 801 51
rect 767 -51 801 -17
rect 767 -119 801 -85
rect 767 -187 801 -153
rect 767 -255 801 -221
rect 767 -323 801 -289
rect 767 -391 801 -357
rect 767 -459 801 -425
rect 767 -527 801 -493
rect 767 -595 801 -561
rect 767 -663 801 -629
rect -697 -762 -663 -728
rect -629 -762 -595 -728
rect -561 -762 -527 -728
rect -493 -762 -459 -728
rect -425 -762 -391 -728
rect -357 -762 -323 -728
rect -289 -762 -255 -728
rect -221 -762 -187 -728
rect -153 -762 -119 -728
rect -85 -762 -51 -728
rect -17 -762 17 -728
rect 51 -762 85 -728
rect 119 -762 153 -728
rect 187 -762 221 -728
rect 255 -762 289 -728
rect 323 -762 357 -728
rect 391 -762 425 -728
rect 459 -762 493 -728
rect 527 -762 561 -728
rect 595 -762 629 -728
rect 663 -762 697 -728
<< xpolycontact >>
rect -671 200 -601 632
rect -671 -632 -601 -200
rect -353 200 -283 632
rect -353 -632 -283 -200
rect -35 200 35 632
rect -35 -632 35 -200
rect 283 200 353 632
rect 283 -632 353 -200
rect 601 200 671 632
rect 601 -632 671 -200
<< xpolyres >>
rect -671 -200 -601 200
rect -353 -200 -283 200
rect -35 -200 35 200
rect 283 -200 353 200
rect 601 -200 671 200
<< locali >>
rect -801 728 -697 762
rect -663 728 -629 762
rect -595 728 -561 762
rect -527 728 -493 762
rect -459 728 -425 762
rect -391 728 -357 762
rect -323 728 -289 762
rect -255 728 -221 762
rect -187 728 -153 762
rect -119 728 -85 762
rect -51 728 -17 762
rect 17 728 51 762
rect 85 728 119 762
rect 153 728 187 762
rect 221 728 255 762
rect 289 728 323 762
rect 357 728 391 762
rect 425 728 459 762
rect 493 728 527 762
rect 561 728 595 762
rect 629 728 663 762
rect 697 728 801 762
rect -801 663 -767 728
rect 767 663 801 728
rect -801 595 -767 629
rect -801 527 -767 561
rect -801 459 -767 493
rect -801 391 -767 425
rect -801 323 -767 357
rect -801 255 -767 289
rect -801 187 -767 221
rect 767 595 801 629
rect 767 527 801 561
rect 767 459 801 493
rect 767 391 801 425
rect 767 323 801 357
rect 767 255 801 289
rect -801 119 -767 153
rect -801 51 -767 85
rect -801 -17 -767 17
rect -801 -85 -767 -51
rect -801 -153 -767 -119
rect -801 -221 -767 -187
rect 767 187 801 221
rect 767 119 801 153
rect 767 51 801 85
rect 767 -17 801 17
rect 767 -85 801 -51
rect 767 -153 801 -119
rect -801 -289 -767 -255
rect -801 -357 -767 -323
rect -801 -425 -767 -391
rect -801 -493 -767 -459
rect -801 -561 -767 -527
rect -801 -629 -767 -595
rect 767 -221 801 -187
rect 767 -289 801 -255
rect 767 -357 801 -323
rect 767 -425 801 -391
rect 767 -493 801 -459
rect 767 -561 801 -527
rect 767 -629 801 -595
rect -801 -728 -767 -663
rect 767 -728 801 -663
rect -801 -762 -697 -728
rect -663 -762 -629 -728
rect -595 -762 -561 -728
rect -527 -762 -493 -728
rect -459 -762 -425 -728
rect -391 -762 -357 -728
rect -323 -762 -289 -728
rect -255 -762 -221 -728
rect -187 -762 -153 -728
rect -119 -762 -85 -728
rect -51 -762 -17 -728
rect 17 -762 51 -728
rect 85 -762 119 -728
rect 153 -762 187 -728
rect 221 -762 255 -728
rect 289 -762 323 -728
rect 357 -762 391 -728
rect 425 -762 459 -728
rect 493 -762 527 -728
rect 561 -762 595 -728
rect 629 -762 663 -728
rect 697 -762 801 -728
<< properties >>
string FIXED_BBOX -784 -745 784 745
<< end >>
