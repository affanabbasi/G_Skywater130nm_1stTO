magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -2879 840 2879 874
rect -2879 -840 -2845 840
rect 2845 -840 2879 840
rect -2879 -874 2879 -840
<< nmoslvt >>
rect -2719 -700 -2319 700
rect -2261 -700 -1861 700
rect -1803 -700 -1403 700
rect -1345 -700 -945 700
rect -887 -700 -487 700
rect -429 -700 -29 700
rect 29 -700 429 700
rect 487 -700 887 700
rect 945 -700 1345 700
rect 1403 -700 1803 700
rect 1861 -700 2261 700
rect 2319 -700 2719 700
<< ndiff >>
rect -2777 663 -2719 700
rect -2777 629 -2765 663
rect -2731 629 -2719 663
rect -2777 595 -2719 629
rect -2777 561 -2765 595
rect -2731 561 -2719 595
rect -2777 527 -2719 561
rect -2777 493 -2765 527
rect -2731 493 -2719 527
rect -2777 459 -2719 493
rect -2777 425 -2765 459
rect -2731 425 -2719 459
rect -2777 391 -2719 425
rect -2777 357 -2765 391
rect -2731 357 -2719 391
rect -2777 323 -2719 357
rect -2777 289 -2765 323
rect -2731 289 -2719 323
rect -2777 255 -2719 289
rect -2777 221 -2765 255
rect -2731 221 -2719 255
rect -2777 187 -2719 221
rect -2777 153 -2765 187
rect -2731 153 -2719 187
rect -2777 119 -2719 153
rect -2777 85 -2765 119
rect -2731 85 -2719 119
rect -2777 51 -2719 85
rect -2777 17 -2765 51
rect -2731 17 -2719 51
rect -2777 -17 -2719 17
rect -2777 -51 -2765 -17
rect -2731 -51 -2719 -17
rect -2777 -85 -2719 -51
rect -2777 -119 -2765 -85
rect -2731 -119 -2719 -85
rect -2777 -153 -2719 -119
rect -2777 -187 -2765 -153
rect -2731 -187 -2719 -153
rect -2777 -221 -2719 -187
rect -2777 -255 -2765 -221
rect -2731 -255 -2719 -221
rect -2777 -289 -2719 -255
rect -2777 -323 -2765 -289
rect -2731 -323 -2719 -289
rect -2777 -357 -2719 -323
rect -2777 -391 -2765 -357
rect -2731 -391 -2719 -357
rect -2777 -425 -2719 -391
rect -2777 -459 -2765 -425
rect -2731 -459 -2719 -425
rect -2777 -493 -2719 -459
rect -2777 -527 -2765 -493
rect -2731 -527 -2719 -493
rect -2777 -561 -2719 -527
rect -2777 -595 -2765 -561
rect -2731 -595 -2719 -561
rect -2777 -629 -2719 -595
rect -2777 -663 -2765 -629
rect -2731 -663 -2719 -629
rect -2777 -700 -2719 -663
rect -2319 663 -2261 700
rect -2319 629 -2307 663
rect -2273 629 -2261 663
rect -2319 595 -2261 629
rect -2319 561 -2307 595
rect -2273 561 -2261 595
rect -2319 527 -2261 561
rect -2319 493 -2307 527
rect -2273 493 -2261 527
rect -2319 459 -2261 493
rect -2319 425 -2307 459
rect -2273 425 -2261 459
rect -2319 391 -2261 425
rect -2319 357 -2307 391
rect -2273 357 -2261 391
rect -2319 323 -2261 357
rect -2319 289 -2307 323
rect -2273 289 -2261 323
rect -2319 255 -2261 289
rect -2319 221 -2307 255
rect -2273 221 -2261 255
rect -2319 187 -2261 221
rect -2319 153 -2307 187
rect -2273 153 -2261 187
rect -2319 119 -2261 153
rect -2319 85 -2307 119
rect -2273 85 -2261 119
rect -2319 51 -2261 85
rect -2319 17 -2307 51
rect -2273 17 -2261 51
rect -2319 -17 -2261 17
rect -2319 -51 -2307 -17
rect -2273 -51 -2261 -17
rect -2319 -85 -2261 -51
rect -2319 -119 -2307 -85
rect -2273 -119 -2261 -85
rect -2319 -153 -2261 -119
rect -2319 -187 -2307 -153
rect -2273 -187 -2261 -153
rect -2319 -221 -2261 -187
rect -2319 -255 -2307 -221
rect -2273 -255 -2261 -221
rect -2319 -289 -2261 -255
rect -2319 -323 -2307 -289
rect -2273 -323 -2261 -289
rect -2319 -357 -2261 -323
rect -2319 -391 -2307 -357
rect -2273 -391 -2261 -357
rect -2319 -425 -2261 -391
rect -2319 -459 -2307 -425
rect -2273 -459 -2261 -425
rect -2319 -493 -2261 -459
rect -2319 -527 -2307 -493
rect -2273 -527 -2261 -493
rect -2319 -561 -2261 -527
rect -2319 -595 -2307 -561
rect -2273 -595 -2261 -561
rect -2319 -629 -2261 -595
rect -2319 -663 -2307 -629
rect -2273 -663 -2261 -629
rect -2319 -700 -2261 -663
rect -1861 663 -1803 700
rect -1861 629 -1849 663
rect -1815 629 -1803 663
rect -1861 595 -1803 629
rect -1861 561 -1849 595
rect -1815 561 -1803 595
rect -1861 527 -1803 561
rect -1861 493 -1849 527
rect -1815 493 -1803 527
rect -1861 459 -1803 493
rect -1861 425 -1849 459
rect -1815 425 -1803 459
rect -1861 391 -1803 425
rect -1861 357 -1849 391
rect -1815 357 -1803 391
rect -1861 323 -1803 357
rect -1861 289 -1849 323
rect -1815 289 -1803 323
rect -1861 255 -1803 289
rect -1861 221 -1849 255
rect -1815 221 -1803 255
rect -1861 187 -1803 221
rect -1861 153 -1849 187
rect -1815 153 -1803 187
rect -1861 119 -1803 153
rect -1861 85 -1849 119
rect -1815 85 -1803 119
rect -1861 51 -1803 85
rect -1861 17 -1849 51
rect -1815 17 -1803 51
rect -1861 -17 -1803 17
rect -1861 -51 -1849 -17
rect -1815 -51 -1803 -17
rect -1861 -85 -1803 -51
rect -1861 -119 -1849 -85
rect -1815 -119 -1803 -85
rect -1861 -153 -1803 -119
rect -1861 -187 -1849 -153
rect -1815 -187 -1803 -153
rect -1861 -221 -1803 -187
rect -1861 -255 -1849 -221
rect -1815 -255 -1803 -221
rect -1861 -289 -1803 -255
rect -1861 -323 -1849 -289
rect -1815 -323 -1803 -289
rect -1861 -357 -1803 -323
rect -1861 -391 -1849 -357
rect -1815 -391 -1803 -357
rect -1861 -425 -1803 -391
rect -1861 -459 -1849 -425
rect -1815 -459 -1803 -425
rect -1861 -493 -1803 -459
rect -1861 -527 -1849 -493
rect -1815 -527 -1803 -493
rect -1861 -561 -1803 -527
rect -1861 -595 -1849 -561
rect -1815 -595 -1803 -561
rect -1861 -629 -1803 -595
rect -1861 -663 -1849 -629
rect -1815 -663 -1803 -629
rect -1861 -700 -1803 -663
rect -1403 663 -1345 700
rect -1403 629 -1391 663
rect -1357 629 -1345 663
rect -1403 595 -1345 629
rect -1403 561 -1391 595
rect -1357 561 -1345 595
rect -1403 527 -1345 561
rect -1403 493 -1391 527
rect -1357 493 -1345 527
rect -1403 459 -1345 493
rect -1403 425 -1391 459
rect -1357 425 -1345 459
rect -1403 391 -1345 425
rect -1403 357 -1391 391
rect -1357 357 -1345 391
rect -1403 323 -1345 357
rect -1403 289 -1391 323
rect -1357 289 -1345 323
rect -1403 255 -1345 289
rect -1403 221 -1391 255
rect -1357 221 -1345 255
rect -1403 187 -1345 221
rect -1403 153 -1391 187
rect -1357 153 -1345 187
rect -1403 119 -1345 153
rect -1403 85 -1391 119
rect -1357 85 -1345 119
rect -1403 51 -1345 85
rect -1403 17 -1391 51
rect -1357 17 -1345 51
rect -1403 -17 -1345 17
rect -1403 -51 -1391 -17
rect -1357 -51 -1345 -17
rect -1403 -85 -1345 -51
rect -1403 -119 -1391 -85
rect -1357 -119 -1345 -85
rect -1403 -153 -1345 -119
rect -1403 -187 -1391 -153
rect -1357 -187 -1345 -153
rect -1403 -221 -1345 -187
rect -1403 -255 -1391 -221
rect -1357 -255 -1345 -221
rect -1403 -289 -1345 -255
rect -1403 -323 -1391 -289
rect -1357 -323 -1345 -289
rect -1403 -357 -1345 -323
rect -1403 -391 -1391 -357
rect -1357 -391 -1345 -357
rect -1403 -425 -1345 -391
rect -1403 -459 -1391 -425
rect -1357 -459 -1345 -425
rect -1403 -493 -1345 -459
rect -1403 -527 -1391 -493
rect -1357 -527 -1345 -493
rect -1403 -561 -1345 -527
rect -1403 -595 -1391 -561
rect -1357 -595 -1345 -561
rect -1403 -629 -1345 -595
rect -1403 -663 -1391 -629
rect -1357 -663 -1345 -629
rect -1403 -700 -1345 -663
rect -945 663 -887 700
rect -945 629 -933 663
rect -899 629 -887 663
rect -945 595 -887 629
rect -945 561 -933 595
rect -899 561 -887 595
rect -945 527 -887 561
rect -945 493 -933 527
rect -899 493 -887 527
rect -945 459 -887 493
rect -945 425 -933 459
rect -899 425 -887 459
rect -945 391 -887 425
rect -945 357 -933 391
rect -899 357 -887 391
rect -945 323 -887 357
rect -945 289 -933 323
rect -899 289 -887 323
rect -945 255 -887 289
rect -945 221 -933 255
rect -899 221 -887 255
rect -945 187 -887 221
rect -945 153 -933 187
rect -899 153 -887 187
rect -945 119 -887 153
rect -945 85 -933 119
rect -899 85 -887 119
rect -945 51 -887 85
rect -945 17 -933 51
rect -899 17 -887 51
rect -945 -17 -887 17
rect -945 -51 -933 -17
rect -899 -51 -887 -17
rect -945 -85 -887 -51
rect -945 -119 -933 -85
rect -899 -119 -887 -85
rect -945 -153 -887 -119
rect -945 -187 -933 -153
rect -899 -187 -887 -153
rect -945 -221 -887 -187
rect -945 -255 -933 -221
rect -899 -255 -887 -221
rect -945 -289 -887 -255
rect -945 -323 -933 -289
rect -899 -323 -887 -289
rect -945 -357 -887 -323
rect -945 -391 -933 -357
rect -899 -391 -887 -357
rect -945 -425 -887 -391
rect -945 -459 -933 -425
rect -899 -459 -887 -425
rect -945 -493 -887 -459
rect -945 -527 -933 -493
rect -899 -527 -887 -493
rect -945 -561 -887 -527
rect -945 -595 -933 -561
rect -899 -595 -887 -561
rect -945 -629 -887 -595
rect -945 -663 -933 -629
rect -899 -663 -887 -629
rect -945 -700 -887 -663
rect -487 663 -429 700
rect -487 629 -475 663
rect -441 629 -429 663
rect -487 595 -429 629
rect -487 561 -475 595
rect -441 561 -429 595
rect -487 527 -429 561
rect -487 493 -475 527
rect -441 493 -429 527
rect -487 459 -429 493
rect -487 425 -475 459
rect -441 425 -429 459
rect -487 391 -429 425
rect -487 357 -475 391
rect -441 357 -429 391
rect -487 323 -429 357
rect -487 289 -475 323
rect -441 289 -429 323
rect -487 255 -429 289
rect -487 221 -475 255
rect -441 221 -429 255
rect -487 187 -429 221
rect -487 153 -475 187
rect -441 153 -429 187
rect -487 119 -429 153
rect -487 85 -475 119
rect -441 85 -429 119
rect -487 51 -429 85
rect -487 17 -475 51
rect -441 17 -429 51
rect -487 -17 -429 17
rect -487 -51 -475 -17
rect -441 -51 -429 -17
rect -487 -85 -429 -51
rect -487 -119 -475 -85
rect -441 -119 -429 -85
rect -487 -153 -429 -119
rect -487 -187 -475 -153
rect -441 -187 -429 -153
rect -487 -221 -429 -187
rect -487 -255 -475 -221
rect -441 -255 -429 -221
rect -487 -289 -429 -255
rect -487 -323 -475 -289
rect -441 -323 -429 -289
rect -487 -357 -429 -323
rect -487 -391 -475 -357
rect -441 -391 -429 -357
rect -487 -425 -429 -391
rect -487 -459 -475 -425
rect -441 -459 -429 -425
rect -487 -493 -429 -459
rect -487 -527 -475 -493
rect -441 -527 -429 -493
rect -487 -561 -429 -527
rect -487 -595 -475 -561
rect -441 -595 -429 -561
rect -487 -629 -429 -595
rect -487 -663 -475 -629
rect -441 -663 -429 -629
rect -487 -700 -429 -663
rect -29 663 29 700
rect -29 629 -17 663
rect 17 629 29 663
rect -29 595 29 629
rect -29 561 -17 595
rect 17 561 29 595
rect -29 527 29 561
rect -29 493 -17 527
rect 17 493 29 527
rect -29 459 29 493
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -493 29 -459
rect -29 -527 -17 -493
rect 17 -527 29 -493
rect -29 -561 29 -527
rect -29 -595 -17 -561
rect 17 -595 29 -561
rect -29 -629 29 -595
rect -29 -663 -17 -629
rect 17 -663 29 -629
rect -29 -700 29 -663
rect 429 663 487 700
rect 429 629 441 663
rect 475 629 487 663
rect 429 595 487 629
rect 429 561 441 595
rect 475 561 487 595
rect 429 527 487 561
rect 429 493 441 527
rect 475 493 487 527
rect 429 459 487 493
rect 429 425 441 459
rect 475 425 487 459
rect 429 391 487 425
rect 429 357 441 391
rect 475 357 487 391
rect 429 323 487 357
rect 429 289 441 323
rect 475 289 487 323
rect 429 255 487 289
rect 429 221 441 255
rect 475 221 487 255
rect 429 187 487 221
rect 429 153 441 187
rect 475 153 487 187
rect 429 119 487 153
rect 429 85 441 119
rect 475 85 487 119
rect 429 51 487 85
rect 429 17 441 51
rect 475 17 487 51
rect 429 -17 487 17
rect 429 -51 441 -17
rect 475 -51 487 -17
rect 429 -85 487 -51
rect 429 -119 441 -85
rect 475 -119 487 -85
rect 429 -153 487 -119
rect 429 -187 441 -153
rect 475 -187 487 -153
rect 429 -221 487 -187
rect 429 -255 441 -221
rect 475 -255 487 -221
rect 429 -289 487 -255
rect 429 -323 441 -289
rect 475 -323 487 -289
rect 429 -357 487 -323
rect 429 -391 441 -357
rect 475 -391 487 -357
rect 429 -425 487 -391
rect 429 -459 441 -425
rect 475 -459 487 -425
rect 429 -493 487 -459
rect 429 -527 441 -493
rect 475 -527 487 -493
rect 429 -561 487 -527
rect 429 -595 441 -561
rect 475 -595 487 -561
rect 429 -629 487 -595
rect 429 -663 441 -629
rect 475 -663 487 -629
rect 429 -700 487 -663
rect 887 663 945 700
rect 887 629 899 663
rect 933 629 945 663
rect 887 595 945 629
rect 887 561 899 595
rect 933 561 945 595
rect 887 527 945 561
rect 887 493 899 527
rect 933 493 945 527
rect 887 459 945 493
rect 887 425 899 459
rect 933 425 945 459
rect 887 391 945 425
rect 887 357 899 391
rect 933 357 945 391
rect 887 323 945 357
rect 887 289 899 323
rect 933 289 945 323
rect 887 255 945 289
rect 887 221 899 255
rect 933 221 945 255
rect 887 187 945 221
rect 887 153 899 187
rect 933 153 945 187
rect 887 119 945 153
rect 887 85 899 119
rect 933 85 945 119
rect 887 51 945 85
rect 887 17 899 51
rect 933 17 945 51
rect 887 -17 945 17
rect 887 -51 899 -17
rect 933 -51 945 -17
rect 887 -85 945 -51
rect 887 -119 899 -85
rect 933 -119 945 -85
rect 887 -153 945 -119
rect 887 -187 899 -153
rect 933 -187 945 -153
rect 887 -221 945 -187
rect 887 -255 899 -221
rect 933 -255 945 -221
rect 887 -289 945 -255
rect 887 -323 899 -289
rect 933 -323 945 -289
rect 887 -357 945 -323
rect 887 -391 899 -357
rect 933 -391 945 -357
rect 887 -425 945 -391
rect 887 -459 899 -425
rect 933 -459 945 -425
rect 887 -493 945 -459
rect 887 -527 899 -493
rect 933 -527 945 -493
rect 887 -561 945 -527
rect 887 -595 899 -561
rect 933 -595 945 -561
rect 887 -629 945 -595
rect 887 -663 899 -629
rect 933 -663 945 -629
rect 887 -700 945 -663
rect 1345 663 1403 700
rect 1345 629 1357 663
rect 1391 629 1403 663
rect 1345 595 1403 629
rect 1345 561 1357 595
rect 1391 561 1403 595
rect 1345 527 1403 561
rect 1345 493 1357 527
rect 1391 493 1403 527
rect 1345 459 1403 493
rect 1345 425 1357 459
rect 1391 425 1403 459
rect 1345 391 1403 425
rect 1345 357 1357 391
rect 1391 357 1403 391
rect 1345 323 1403 357
rect 1345 289 1357 323
rect 1391 289 1403 323
rect 1345 255 1403 289
rect 1345 221 1357 255
rect 1391 221 1403 255
rect 1345 187 1403 221
rect 1345 153 1357 187
rect 1391 153 1403 187
rect 1345 119 1403 153
rect 1345 85 1357 119
rect 1391 85 1403 119
rect 1345 51 1403 85
rect 1345 17 1357 51
rect 1391 17 1403 51
rect 1345 -17 1403 17
rect 1345 -51 1357 -17
rect 1391 -51 1403 -17
rect 1345 -85 1403 -51
rect 1345 -119 1357 -85
rect 1391 -119 1403 -85
rect 1345 -153 1403 -119
rect 1345 -187 1357 -153
rect 1391 -187 1403 -153
rect 1345 -221 1403 -187
rect 1345 -255 1357 -221
rect 1391 -255 1403 -221
rect 1345 -289 1403 -255
rect 1345 -323 1357 -289
rect 1391 -323 1403 -289
rect 1345 -357 1403 -323
rect 1345 -391 1357 -357
rect 1391 -391 1403 -357
rect 1345 -425 1403 -391
rect 1345 -459 1357 -425
rect 1391 -459 1403 -425
rect 1345 -493 1403 -459
rect 1345 -527 1357 -493
rect 1391 -527 1403 -493
rect 1345 -561 1403 -527
rect 1345 -595 1357 -561
rect 1391 -595 1403 -561
rect 1345 -629 1403 -595
rect 1345 -663 1357 -629
rect 1391 -663 1403 -629
rect 1345 -700 1403 -663
rect 1803 663 1861 700
rect 1803 629 1815 663
rect 1849 629 1861 663
rect 1803 595 1861 629
rect 1803 561 1815 595
rect 1849 561 1861 595
rect 1803 527 1861 561
rect 1803 493 1815 527
rect 1849 493 1861 527
rect 1803 459 1861 493
rect 1803 425 1815 459
rect 1849 425 1861 459
rect 1803 391 1861 425
rect 1803 357 1815 391
rect 1849 357 1861 391
rect 1803 323 1861 357
rect 1803 289 1815 323
rect 1849 289 1861 323
rect 1803 255 1861 289
rect 1803 221 1815 255
rect 1849 221 1861 255
rect 1803 187 1861 221
rect 1803 153 1815 187
rect 1849 153 1861 187
rect 1803 119 1861 153
rect 1803 85 1815 119
rect 1849 85 1861 119
rect 1803 51 1861 85
rect 1803 17 1815 51
rect 1849 17 1861 51
rect 1803 -17 1861 17
rect 1803 -51 1815 -17
rect 1849 -51 1861 -17
rect 1803 -85 1861 -51
rect 1803 -119 1815 -85
rect 1849 -119 1861 -85
rect 1803 -153 1861 -119
rect 1803 -187 1815 -153
rect 1849 -187 1861 -153
rect 1803 -221 1861 -187
rect 1803 -255 1815 -221
rect 1849 -255 1861 -221
rect 1803 -289 1861 -255
rect 1803 -323 1815 -289
rect 1849 -323 1861 -289
rect 1803 -357 1861 -323
rect 1803 -391 1815 -357
rect 1849 -391 1861 -357
rect 1803 -425 1861 -391
rect 1803 -459 1815 -425
rect 1849 -459 1861 -425
rect 1803 -493 1861 -459
rect 1803 -527 1815 -493
rect 1849 -527 1861 -493
rect 1803 -561 1861 -527
rect 1803 -595 1815 -561
rect 1849 -595 1861 -561
rect 1803 -629 1861 -595
rect 1803 -663 1815 -629
rect 1849 -663 1861 -629
rect 1803 -700 1861 -663
rect 2261 663 2319 700
rect 2261 629 2273 663
rect 2307 629 2319 663
rect 2261 595 2319 629
rect 2261 561 2273 595
rect 2307 561 2319 595
rect 2261 527 2319 561
rect 2261 493 2273 527
rect 2307 493 2319 527
rect 2261 459 2319 493
rect 2261 425 2273 459
rect 2307 425 2319 459
rect 2261 391 2319 425
rect 2261 357 2273 391
rect 2307 357 2319 391
rect 2261 323 2319 357
rect 2261 289 2273 323
rect 2307 289 2319 323
rect 2261 255 2319 289
rect 2261 221 2273 255
rect 2307 221 2319 255
rect 2261 187 2319 221
rect 2261 153 2273 187
rect 2307 153 2319 187
rect 2261 119 2319 153
rect 2261 85 2273 119
rect 2307 85 2319 119
rect 2261 51 2319 85
rect 2261 17 2273 51
rect 2307 17 2319 51
rect 2261 -17 2319 17
rect 2261 -51 2273 -17
rect 2307 -51 2319 -17
rect 2261 -85 2319 -51
rect 2261 -119 2273 -85
rect 2307 -119 2319 -85
rect 2261 -153 2319 -119
rect 2261 -187 2273 -153
rect 2307 -187 2319 -153
rect 2261 -221 2319 -187
rect 2261 -255 2273 -221
rect 2307 -255 2319 -221
rect 2261 -289 2319 -255
rect 2261 -323 2273 -289
rect 2307 -323 2319 -289
rect 2261 -357 2319 -323
rect 2261 -391 2273 -357
rect 2307 -391 2319 -357
rect 2261 -425 2319 -391
rect 2261 -459 2273 -425
rect 2307 -459 2319 -425
rect 2261 -493 2319 -459
rect 2261 -527 2273 -493
rect 2307 -527 2319 -493
rect 2261 -561 2319 -527
rect 2261 -595 2273 -561
rect 2307 -595 2319 -561
rect 2261 -629 2319 -595
rect 2261 -663 2273 -629
rect 2307 -663 2319 -629
rect 2261 -700 2319 -663
rect 2719 663 2777 700
rect 2719 629 2731 663
rect 2765 629 2777 663
rect 2719 595 2777 629
rect 2719 561 2731 595
rect 2765 561 2777 595
rect 2719 527 2777 561
rect 2719 493 2731 527
rect 2765 493 2777 527
rect 2719 459 2777 493
rect 2719 425 2731 459
rect 2765 425 2777 459
rect 2719 391 2777 425
rect 2719 357 2731 391
rect 2765 357 2777 391
rect 2719 323 2777 357
rect 2719 289 2731 323
rect 2765 289 2777 323
rect 2719 255 2777 289
rect 2719 221 2731 255
rect 2765 221 2777 255
rect 2719 187 2777 221
rect 2719 153 2731 187
rect 2765 153 2777 187
rect 2719 119 2777 153
rect 2719 85 2731 119
rect 2765 85 2777 119
rect 2719 51 2777 85
rect 2719 17 2731 51
rect 2765 17 2777 51
rect 2719 -17 2777 17
rect 2719 -51 2731 -17
rect 2765 -51 2777 -17
rect 2719 -85 2777 -51
rect 2719 -119 2731 -85
rect 2765 -119 2777 -85
rect 2719 -153 2777 -119
rect 2719 -187 2731 -153
rect 2765 -187 2777 -153
rect 2719 -221 2777 -187
rect 2719 -255 2731 -221
rect 2765 -255 2777 -221
rect 2719 -289 2777 -255
rect 2719 -323 2731 -289
rect 2765 -323 2777 -289
rect 2719 -357 2777 -323
rect 2719 -391 2731 -357
rect 2765 -391 2777 -357
rect 2719 -425 2777 -391
rect 2719 -459 2731 -425
rect 2765 -459 2777 -425
rect 2719 -493 2777 -459
rect 2719 -527 2731 -493
rect 2765 -527 2777 -493
rect 2719 -561 2777 -527
rect 2719 -595 2731 -561
rect 2765 -595 2777 -561
rect 2719 -629 2777 -595
rect 2719 -663 2731 -629
rect 2765 -663 2777 -629
rect 2719 -700 2777 -663
<< ndiffc >>
rect -2765 629 -2731 663
rect -2765 561 -2731 595
rect -2765 493 -2731 527
rect -2765 425 -2731 459
rect -2765 357 -2731 391
rect -2765 289 -2731 323
rect -2765 221 -2731 255
rect -2765 153 -2731 187
rect -2765 85 -2731 119
rect -2765 17 -2731 51
rect -2765 -51 -2731 -17
rect -2765 -119 -2731 -85
rect -2765 -187 -2731 -153
rect -2765 -255 -2731 -221
rect -2765 -323 -2731 -289
rect -2765 -391 -2731 -357
rect -2765 -459 -2731 -425
rect -2765 -527 -2731 -493
rect -2765 -595 -2731 -561
rect -2765 -663 -2731 -629
rect -2307 629 -2273 663
rect -2307 561 -2273 595
rect -2307 493 -2273 527
rect -2307 425 -2273 459
rect -2307 357 -2273 391
rect -2307 289 -2273 323
rect -2307 221 -2273 255
rect -2307 153 -2273 187
rect -2307 85 -2273 119
rect -2307 17 -2273 51
rect -2307 -51 -2273 -17
rect -2307 -119 -2273 -85
rect -2307 -187 -2273 -153
rect -2307 -255 -2273 -221
rect -2307 -323 -2273 -289
rect -2307 -391 -2273 -357
rect -2307 -459 -2273 -425
rect -2307 -527 -2273 -493
rect -2307 -595 -2273 -561
rect -2307 -663 -2273 -629
rect -1849 629 -1815 663
rect -1849 561 -1815 595
rect -1849 493 -1815 527
rect -1849 425 -1815 459
rect -1849 357 -1815 391
rect -1849 289 -1815 323
rect -1849 221 -1815 255
rect -1849 153 -1815 187
rect -1849 85 -1815 119
rect -1849 17 -1815 51
rect -1849 -51 -1815 -17
rect -1849 -119 -1815 -85
rect -1849 -187 -1815 -153
rect -1849 -255 -1815 -221
rect -1849 -323 -1815 -289
rect -1849 -391 -1815 -357
rect -1849 -459 -1815 -425
rect -1849 -527 -1815 -493
rect -1849 -595 -1815 -561
rect -1849 -663 -1815 -629
rect -1391 629 -1357 663
rect -1391 561 -1357 595
rect -1391 493 -1357 527
rect -1391 425 -1357 459
rect -1391 357 -1357 391
rect -1391 289 -1357 323
rect -1391 221 -1357 255
rect -1391 153 -1357 187
rect -1391 85 -1357 119
rect -1391 17 -1357 51
rect -1391 -51 -1357 -17
rect -1391 -119 -1357 -85
rect -1391 -187 -1357 -153
rect -1391 -255 -1357 -221
rect -1391 -323 -1357 -289
rect -1391 -391 -1357 -357
rect -1391 -459 -1357 -425
rect -1391 -527 -1357 -493
rect -1391 -595 -1357 -561
rect -1391 -663 -1357 -629
rect -933 629 -899 663
rect -933 561 -899 595
rect -933 493 -899 527
rect -933 425 -899 459
rect -933 357 -899 391
rect -933 289 -899 323
rect -933 221 -899 255
rect -933 153 -899 187
rect -933 85 -899 119
rect -933 17 -899 51
rect -933 -51 -899 -17
rect -933 -119 -899 -85
rect -933 -187 -899 -153
rect -933 -255 -899 -221
rect -933 -323 -899 -289
rect -933 -391 -899 -357
rect -933 -459 -899 -425
rect -933 -527 -899 -493
rect -933 -595 -899 -561
rect -933 -663 -899 -629
rect -475 629 -441 663
rect -475 561 -441 595
rect -475 493 -441 527
rect -475 425 -441 459
rect -475 357 -441 391
rect -475 289 -441 323
rect -475 221 -441 255
rect -475 153 -441 187
rect -475 85 -441 119
rect -475 17 -441 51
rect -475 -51 -441 -17
rect -475 -119 -441 -85
rect -475 -187 -441 -153
rect -475 -255 -441 -221
rect -475 -323 -441 -289
rect -475 -391 -441 -357
rect -475 -459 -441 -425
rect -475 -527 -441 -493
rect -475 -595 -441 -561
rect -475 -663 -441 -629
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect 441 629 475 663
rect 441 561 475 595
rect 441 493 475 527
rect 441 425 475 459
rect 441 357 475 391
rect 441 289 475 323
rect 441 221 475 255
rect 441 153 475 187
rect 441 85 475 119
rect 441 17 475 51
rect 441 -51 475 -17
rect 441 -119 475 -85
rect 441 -187 475 -153
rect 441 -255 475 -221
rect 441 -323 475 -289
rect 441 -391 475 -357
rect 441 -459 475 -425
rect 441 -527 475 -493
rect 441 -595 475 -561
rect 441 -663 475 -629
rect 899 629 933 663
rect 899 561 933 595
rect 899 493 933 527
rect 899 425 933 459
rect 899 357 933 391
rect 899 289 933 323
rect 899 221 933 255
rect 899 153 933 187
rect 899 85 933 119
rect 899 17 933 51
rect 899 -51 933 -17
rect 899 -119 933 -85
rect 899 -187 933 -153
rect 899 -255 933 -221
rect 899 -323 933 -289
rect 899 -391 933 -357
rect 899 -459 933 -425
rect 899 -527 933 -493
rect 899 -595 933 -561
rect 899 -663 933 -629
rect 1357 629 1391 663
rect 1357 561 1391 595
rect 1357 493 1391 527
rect 1357 425 1391 459
rect 1357 357 1391 391
rect 1357 289 1391 323
rect 1357 221 1391 255
rect 1357 153 1391 187
rect 1357 85 1391 119
rect 1357 17 1391 51
rect 1357 -51 1391 -17
rect 1357 -119 1391 -85
rect 1357 -187 1391 -153
rect 1357 -255 1391 -221
rect 1357 -323 1391 -289
rect 1357 -391 1391 -357
rect 1357 -459 1391 -425
rect 1357 -527 1391 -493
rect 1357 -595 1391 -561
rect 1357 -663 1391 -629
rect 1815 629 1849 663
rect 1815 561 1849 595
rect 1815 493 1849 527
rect 1815 425 1849 459
rect 1815 357 1849 391
rect 1815 289 1849 323
rect 1815 221 1849 255
rect 1815 153 1849 187
rect 1815 85 1849 119
rect 1815 17 1849 51
rect 1815 -51 1849 -17
rect 1815 -119 1849 -85
rect 1815 -187 1849 -153
rect 1815 -255 1849 -221
rect 1815 -323 1849 -289
rect 1815 -391 1849 -357
rect 1815 -459 1849 -425
rect 1815 -527 1849 -493
rect 1815 -595 1849 -561
rect 1815 -663 1849 -629
rect 2273 629 2307 663
rect 2273 561 2307 595
rect 2273 493 2307 527
rect 2273 425 2307 459
rect 2273 357 2307 391
rect 2273 289 2307 323
rect 2273 221 2307 255
rect 2273 153 2307 187
rect 2273 85 2307 119
rect 2273 17 2307 51
rect 2273 -51 2307 -17
rect 2273 -119 2307 -85
rect 2273 -187 2307 -153
rect 2273 -255 2307 -221
rect 2273 -323 2307 -289
rect 2273 -391 2307 -357
rect 2273 -459 2307 -425
rect 2273 -527 2307 -493
rect 2273 -595 2307 -561
rect 2273 -663 2307 -629
rect 2731 629 2765 663
rect 2731 561 2765 595
rect 2731 493 2765 527
rect 2731 425 2765 459
rect 2731 357 2765 391
rect 2731 289 2765 323
rect 2731 221 2765 255
rect 2731 153 2765 187
rect 2731 85 2765 119
rect 2731 17 2765 51
rect 2731 -51 2765 -17
rect 2731 -119 2765 -85
rect 2731 -187 2765 -153
rect 2731 -255 2765 -221
rect 2731 -323 2765 -289
rect 2731 -391 2765 -357
rect 2731 -459 2765 -425
rect 2731 -527 2765 -493
rect 2731 -595 2765 -561
rect 2731 -663 2765 -629
<< psubdiff >>
rect -2879 840 -2771 874
rect -2737 840 -2703 874
rect -2669 840 -2635 874
rect -2601 840 -2567 874
rect -2533 840 -2499 874
rect -2465 840 -2431 874
rect -2397 840 -2363 874
rect -2329 840 -2295 874
rect -2261 840 -2227 874
rect -2193 840 -2159 874
rect -2125 840 -2091 874
rect -2057 840 -2023 874
rect -1989 840 -1955 874
rect -1921 840 -1887 874
rect -1853 840 -1819 874
rect -1785 840 -1751 874
rect -1717 840 -1683 874
rect -1649 840 -1615 874
rect -1581 840 -1547 874
rect -1513 840 -1479 874
rect -1445 840 -1411 874
rect -1377 840 -1343 874
rect -1309 840 -1275 874
rect -1241 840 -1207 874
rect -1173 840 -1139 874
rect -1105 840 -1071 874
rect -1037 840 -1003 874
rect -969 840 -935 874
rect -901 840 -867 874
rect -833 840 -799 874
rect -765 840 -731 874
rect -697 840 -663 874
rect -629 840 -595 874
rect -561 840 -527 874
rect -493 840 -459 874
rect -425 840 -391 874
rect -357 840 -323 874
rect -289 840 -255 874
rect -221 840 -187 874
rect -153 840 -119 874
rect -85 840 -51 874
rect -17 840 17 874
rect 51 840 85 874
rect 119 840 153 874
rect 187 840 221 874
rect 255 840 289 874
rect 323 840 357 874
rect 391 840 425 874
rect 459 840 493 874
rect 527 840 561 874
rect 595 840 629 874
rect 663 840 697 874
rect 731 840 765 874
rect 799 840 833 874
rect 867 840 901 874
rect 935 840 969 874
rect 1003 840 1037 874
rect 1071 840 1105 874
rect 1139 840 1173 874
rect 1207 840 1241 874
rect 1275 840 1309 874
rect 1343 840 1377 874
rect 1411 840 1445 874
rect 1479 840 1513 874
rect 1547 840 1581 874
rect 1615 840 1649 874
rect 1683 840 1717 874
rect 1751 840 1785 874
rect 1819 840 1853 874
rect 1887 840 1921 874
rect 1955 840 1989 874
rect 2023 840 2057 874
rect 2091 840 2125 874
rect 2159 840 2193 874
rect 2227 840 2261 874
rect 2295 840 2329 874
rect 2363 840 2397 874
rect 2431 840 2465 874
rect 2499 840 2533 874
rect 2567 840 2601 874
rect 2635 840 2669 874
rect 2703 840 2737 874
rect 2771 840 2879 874
rect -2879 765 -2845 840
rect -2879 697 -2845 731
rect 2845 765 2879 840
rect -2879 629 -2845 663
rect -2879 561 -2845 595
rect -2879 493 -2845 527
rect -2879 425 -2845 459
rect -2879 357 -2845 391
rect -2879 289 -2845 323
rect -2879 221 -2845 255
rect -2879 153 -2845 187
rect -2879 85 -2845 119
rect -2879 17 -2845 51
rect -2879 -51 -2845 -17
rect -2879 -119 -2845 -85
rect -2879 -187 -2845 -153
rect -2879 -255 -2845 -221
rect -2879 -323 -2845 -289
rect -2879 -391 -2845 -357
rect -2879 -459 -2845 -425
rect -2879 -527 -2845 -493
rect -2879 -595 -2845 -561
rect -2879 -663 -2845 -629
rect -2879 -731 -2845 -697
rect 2845 697 2879 731
rect 2845 629 2879 663
rect 2845 561 2879 595
rect 2845 493 2879 527
rect 2845 425 2879 459
rect 2845 357 2879 391
rect 2845 289 2879 323
rect 2845 221 2879 255
rect 2845 153 2879 187
rect 2845 85 2879 119
rect 2845 17 2879 51
rect 2845 -51 2879 -17
rect 2845 -119 2879 -85
rect 2845 -187 2879 -153
rect 2845 -255 2879 -221
rect 2845 -323 2879 -289
rect 2845 -391 2879 -357
rect 2845 -459 2879 -425
rect 2845 -527 2879 -493
rect 2845 -595 2879 -561
rect 2845 -663 2879 -629
rect -2879 -840 -2845 -765
rect 2845 -731 2879 -697
rect 2845 -840 2879 -765
rect -2879 -874 -2771 -840
rect -2737 -874 -2703 -840
rect -2669 -874 -2635 -840
rect -2601 -874 -2567 -840
rect -2533 -874 -2499 -840
rect -2465 -874 -2431 -840
rect -2397 -874 -2363 -840
rect -2329 -874 -2295 -840
rect -2261 -874 -2227 -840
rect -2193 -874 -2159 -840
rect -2125 -874 -2091 -840
rect -2057 -874 -2023 -840
rect -1989 -874 -1955 -840
rect -1921 -874 -1887 -840
rect -1853 -874 -1819 -840
rect -1785 -874 -1751 -840
rect -1717 -874 -1683 -840
rect -1649 -874 -1615 -840
rect -1581 -874 -1547 -840
rect -1513 -874 -1479 -840
rect -1445 -874 -1411 -840
rect -1377 -874 -1343 -840
rect -1309 -874 -1275 -840
rect -1241 -874 -1207 -840
rect -1173 -874 -1139 -840
rect -1105 -874 -1071 -840
rect -1037 -874 -1003 -840
rect -969 -874 -935 -840
rect -901 -874 -867 -840
rect -833 -874 -799 -840
rect -765 -874 -731 -840
rect -697 -874 -663 -840
rect -629 -874 -595 -840
rect -561 -874 -527 -840
rect -493 -874 -459 -840
rect -425 -874 -391 -840
rect -357 -874 -323 -840
rect -289 -874 -255 -840
rect -221 -874 -187 -840
rect -153 -874 -119 -840
rect -85 -874 -51 -840
rect -17 -874 17 -840
rect 51 -874 85 -840
rect 119 -874 153 -840
rect 187 -874 221 -840
rect 255 -874 289 -840
rect 323 -874 357 -840
rect 391 -874 425 -840
rect 459 -874 493 -840
rect 527 -874 561 -840
rect 595 -874 629 -840
rect 663 -874 697 -840
rect 731 -874 765 -840
rect 799 -874 833 -840
rect 867 -874 901 -840
rect 935 -874 969 -840
rect 1003 -874 1037 -840
rect 1071 -874 1105 -840
rect 1139 -874 1173 -840
rect 1207 -874 1241 -840
rect 1275 -874 1309 -840
rect 1343 -874 1377 -840
rect 1411 -874 1445 -840
rect 1479 -874 1513 -840
rect 1547 -874 1581 -840
rect 1615 -874 1649 -840
rect 1683 -874 1717 -840
rect 1751 -874 1785 -840
rect 1819 -874 1853 -840
rect 1887 -874 1921 -840
rect 1955 -874 1989 -840
rect 2023 -874 2057 -840
rect 2091 -874 2125 -840
rect 2159 -874 2193 -840
rect 2227 -874 2261 -840
rect 2295 -874 2329 -840
rect 2363 -874 2397 -840
rect 2431 -874 2465 -840
rect 2499 -874 2533 -840
rect 2567 -874 2601 -840
rect 2635 -874 2669 -840
rect 2703 -874 2737 -840
rect 2771 -874 2879 -840
<< psubdiffcont >>
rect -2771 840 -2737 874
rect -2703 840 -2669 874
rect -2635 840 -2601 874
rect -2567 840 -2533 874
rect -2499 840 -2465 874
rect -2431 840 -2397 874
rect -2363 840 -2329 874
rect -2295 840 -2261 874
rect -2227 840 -2193 874
rect -2159 840 -2125 874
rect -2091 840 -2057 874
rect -2023 840 -1989 874
rect -1955 840 -1921 874
rect -1887 840 -1853 874
rect -1819 840 -1785 874
rect -1751 840 -1717 874
rect -1683 840 -1649 874
rect -1615 840 -1581 874
rect -1547 840 -1513 874
rect -1479 840 -1445 874
rect -1411 840 -1377 874
rect -1343 840 -1309 874
rect -1275 840 -1241 874
rect -1207 840 -1173 874
rect -1139 840 -1105 874
rect -1071 840 -1037 874
rect -1003 840 -969 874
rect -935 840 -901 874
rect -867 840 -833 874
rect -799 840 -765 874
rect -731 840 -697 874
rect -663 840 -629 874
rect -595 840 -561 874
rect -527 840 -493 874
rect -459 840 -425 874
rect -391 840 -357 874
rect -323 840 -289 874
rect -255 840 -221 874
rect -187 840 -153 874
rect -119 840 -85 874
rect -51 840 -17 874
rect 17 840 51 874
rect 85 840 119 874
rect 153 840 187 874
rect 221 840 255 874
rect 289 840 323 874
rect 357 840 391 874
rect 425 840 459 874
rect 493 840 527 874
rect 561 840 595 874
rect 629 840 663 874
rect 697 840 731 874
rect 765 840 799 874
rect 833 840 867 874
rect 901 840 935 874
rect 969 840 1003 874
rect 1037 840 1071 874
rect 1105 840 1139 874
rect 1173 840 1207 874
rect 1241 840 1275 874
rect 1309 840 1343 874
rect 1377 840 1411 874
rect 1445 840 1479 874
rect 1513 840 1547 874
rect 1581 840 1615 874
rect 1649 840 1683 874
rect 1717 840 1751 874
rect 1785 840 1819 874
rect 1853 840 1887 874
rect 1921 840 1955 874
rect 1989 840 2023 874
rect 2057 840 2091 874
rect 2125 840 2159 874
rect 2193 840 2227 874
rect 2261 840 2295 874
rect 2329 840 2363 874
rect 2397 840 2431 874
rect 2465 840 2499 874
rect 2533 840 2567 874
rect 2601 840 2635 874
rect 2669 840 2703 874
rect 2737 840 2771 874
rect -2879 731 -2845 765
rect 2845 731 2879 765
rect -2879 663 -2845 697
rect -2879 595 -2845 629
rect -2879 527 -2845 561
rect -2879 459 -2845 493
rect -2879 391 -2845 425
rect -2879 323 -2845 357
rect -2879 255 -2845 289
rect -2879 187 -2845 221
rect -2879 119 -2845 153
rect -2879 51 -2845 85
rect -2879 -17 -2845 17
rect -2879 -85 -2845 -51
rect -2879 -153 -2845 -119
rect -2879 -221 -2845 -187
rect -2879 -289 -2845 -255
rect -2879 -357 -2845 -323
rect -2879 -425 -2845 -391
rect -2879 -493 -2845 -459
rect -2879 -561 -2845 -527
rect -2879 -629 -2845 -595
rect -2879 -697 -2845 -663
rect 2845 663 2879 697
rect 2845 595 2879 629
rect 2845 527 2879 561
rect 2845 459 2879 493
rect 2845 391 2879 425
rect 2845 323 2879 357
rect 2845 255 2879 289
rect 2845 187 2879 221
rect 2845 119 2879 153
rect 2845 51 2879 85
rect 2845 -17 2879 17
rect 2845 -85 2879 -51
rect 2845 -153 2879 -119
rect 2845 -221 2879 -187
rect 2845 -289 2879 -255
rect 2845 -357 2879 -323
rect 2845 -425 2879 -391
rect 2845 -493 2879 -459
rect 2845 -561 2879 -527
rect 2845 -629 2879 -595
rect 2845 -697 2879 -663
rect -2879 -765 -2845 -731
rect 2845 -765 2879 -731
rect -2771 -874 -2737 -840
rect -2703 -874 -2669 -840
rect -2635 -874 -2601 -840
rect -2567 -874 -2533 -840
rect -2499 -874 -2465 -840
rect -2431 -874 -2397 -840
rect -2363 -874 -2329 -840
rect -2295 -874 -2261 -840
rect -2227 -874 -2193 -840
rect -2159 -874 -2125 -840
rect -2091 -874 -2057 -840
rect -2023 -874 -1989 -840
rect -1955 -874 -1921 -840
rect -1887 -874 -1853 -840
rect -1819 -874 -1785 -840
rect -1751 -874 -1717 -840
rect -1683 -874 -1649 -840
rect -1615 -874 -1581 -840
rect -1547 -874 -1513 -840
rect -1479 -874 -1445 -840
rect -1411 -874 -1377 -840
rect -1343 -874 -1309 -840
rect -1275 -874 -1241 -840
rect -1207 -874 -1173 -840
rect -1139 -874 -1105 -840
rect -1071 -874 -1037 -840
rect -1003 -874 -969 -840
rect -935 -874 -901 -840
rect -867 -874 -833 -840
rect -799 -874 -765 -840
rect -731 -874 -697 -840
rect -663 -874 -629 -840
rect -595 -874 -561 -840
rect -527 -874 -493 -840
rect -459 -874 -425 -840
rect -391 -874 -357 -840
rect -323 -874 -289 -840
rect -255 -874 -221 -840
rect -187 -874 -153 -840
rect -119 -874 -85 -840
rect -51 -874 -17 -840
rect 17 -874 51 -840
rect 85 -874 119 -840
rect 153 -874 187 -840
rect 221 -874 255 -840
rect 289 -874 323 -840
rect 357 -874 391 -840
rect 425 -874 459 -840
rect 493 -874 527 -840
rect 561 -874 595 -840
rect 629 -874 663 -840
rect 697 -874 731 -840
rect 765 -874 799 -840
rect 833 -874 867 -840
rect 901 -874 935 -840
rect 969 -874 1003 -840
rect 1037 -874 1071 -840
rect 1105 -874 1139 -840
rect 1173 -874 1207 -840
rect 1241 -874 1275 -840
rect 1309 -874 1343 -840
rect 1377 -874 1411 -840
rect 1445 -874 1479 -840
rect 1513 -874 1547 -840
rect 1581 -874 1615 -840
rect 1649 -874 1683 -840
rect 1717 -874 1751 -840
rect 1785 -874 1819 -840
rect 1853 -874 1887 -840
rect 1921 -874 1955 -840
rect 1989 -874 2023 -840
rect 2057 -874 2091 -840
rect 2125 -874 2159 -840
rect 2193 -874 2227 -840
rect 2261 -874 2295 -840
rect 2329 -874 2363 -840
rect 2397 -874 2431 -840
rect 2465 -874 2499 -840
rect 2533 -874 2567 -840
rect 2601 -874 2635 -840
rect 2669 -874 2703 -840
rect 2737 -874 2771 -840
<< poly >>
rect -2719 772 -2319 788
rect -2719 738 -2672 772
rect -2638 738 -2604 772
rect -2570 738 -2536 772
rect -2502 738 -2468 772
rect -2434 738 -2400 772
rect -2366 738 -2319 772
rect -2719 700 -2319 738
rect -2261 772 -1861 788
rect -2261 738 -2214 772
rect -2180 738 -2146 772
rect -2112 738 -2078 772
rect -2044 738 -2010 772
rect -1976 738 -1942 772
rect -1908 738 -1861 772
rect -2261 700 -1861 738
rect -1803 772 -1403 788
rect -1803 738 -1756 772
rect -1722 738 -1688 772
rect -1654 738 -1620 772
rect -1586 738 -1552 772
rect -1518 738 -1484 772
rect -1450 738 -1403 772
rect -1803 700 -1403 738
rect -1345 772 -945 788
rect -1345 738 -1298 772
rect -1264 738 -1230 772
rect -1196 738 -1162 772
rect -1128 738 -1094 772
rect -1060 738 -1026 772
rect -992 738 -945 772
rect -1345 700 -945 738
rect -887 772 -487 788
rect -887 738 -840 772
rect -806 738 -772 772
rect -738 738 -704 772
rect -670 738 -636 772
rect -602 738 -568 772
rect -534 738 -487 772
rect -887 700 -487 738
rect -429 772 -29 788
rect -429 738 -382 772
rect -348 738 -314 772
rect -280 738 -246 772
rect -212 738 -178 772
rect -144 738 -110 772
rect -76 738 -29 772
rect -429 700 -29 738
rect 29 772 429 788
rect 29 738 76 772
rect 110 738 144 772
rect 178 738 212 772
rect 246 738 280 772
rect 314 738 348 772
rect 382 738 429 772
rect 29 700 429 738
rect 487 772 887 788
rect 487 738 534 772
rect 568 738 602 772
rect 636 738 670 772
rect 704 738 738 772
rect 772 738 806 772
rect 840 738 887 772
rect 487 700 887 738
rect 945 772 1345 788
rect 945 738 992 772
rect 1026 738 1060 772
rect 1094 738 1128 772
rect 1162 738 1196 772
rect 1230 738 1264 772
rect 1298 738 1345 772
rect 945 700 1345 738
rect 1403 772 1803 788
rect 1403 738 1450 772
rect 1484 738 1518 772
rect 1552 738 1586 772
rect 1620 738 1654 772
rect 1688 738 1722 772
rect 1756 738 1803 772
rect 1403 700 1803 738
rect 1861 772 2261 788
rect 1861 738 1908 772
rect 1942 738 1976 772
rect 2010 738 2044 772
rect 2078 738 2112 772
rect 2146 738 2180 772
rect 2214 738 2261 772
rect 1861 700 2261 738
rect 2319 772 2719 788
rect 2319 738 2366 772
rect 2400 738 2434 772
rect 2468 738 2502 772
rect 2536 738 2570 772
rect 2604 738 2638 772
rect 2672 738 2719 772
rect 2319 700 2719 738
rect -2719 -738 -2319 -700
rect -2719 -772 -2672 -738
rect -2638 -772 -2604 -738
rect -2570 -772 -2536 -738
rect -2502 -772 -2468 -738
rect -2434 -772 -2400 -738
rect -2366 -772 -2319 -738
rect -2719 -788 -2319 -772
rect -2261 -738 -1861 -700
rect -2261 -772 -2214 -738
rect -2180 -772 -2146 -738
rect -2112 -772 -2078 -738
rect -2044 -772 -2010 -738
rect -1976 -772 -1942 -738
rect -1908 -772 -1861 -738
rect -2261 -788 -1861 -772
rect -1803 -738 -1403 -700
rect -1803 -772 -1756 -738
rect -1722 -772 -1688 -738
rect -1654 -772 -1620 -738
rect -1586 -772 -1552 -738
rect -1518 -772 -1484 -738
rect -1450 -772 -1403 -738
rect -1803 -788 -1403 -772
rect -1345 -738 -945 -700
rect -1345 -772 -1298 -738
rect -1264 -772 -1230 -738
rect -1196 -772 -1162 -738
rect -1128 -772 -1094 -738
rect -1060 -772 -1026 -738
rect -992 -772 -945 -738
rect -1345 -788 -945 -772
rect -887 -738 -487 -700
rect -887 -772 -840 -738
rect -806 -772 -772 -738
rect -738 -772 -704 -738
rect -670 -772 -636 -738
rect -602 -772 -568 -738
rect -534 -772 -487 -738
rect -887 -788 -487 -772
rect -429 -738 -29 -700
rect -429 -772 -382 -738
rect -348 -772 -314 -738
rect -280 -772 -246 -738
rect -212 -772 -178 -738
rect -144 -772 -110 -738
rect -76 -772 -29 -738
rect -429 -788 -29 -772
rect 29 -738 429 -700
rect 29 -772 76 -738
rect 110 -772 144 -738
rect 178 -772 212 -738
rect 246 -772 280 -738
rect 314 -772 348 -738
rect 382 -772 429 -738
rect 29 -788 429 -772
rect 487 -738 887 -700
rect 487 -772 534 -738
rect 568 -772 602 -738
rect 636 -772 670 -738
rect 704 -772 738 -738
rect 772 -772 806 -738
rect 840 -772 887 -738
rect 487 -788 887 -772
rect 945 -738 1345 -700
rect 945 -772 992 -738
rect 1026 -772 1060 -738
rect 1094 -772 1128 -738
rect 1162 -772 1196 -738
rect 1230 -772 1264 -738
rect 1298 -772 1345 -738
rect 945 -788 1345 -772
rect 1403 -738 1803 -700
rect 1403 -772 1450 -738
rect 1484 -772 1518 -738
rect 1552 -772 1586 -738
rect 1620 -772 1654 -738
rect 1688 -772 1722 -738
rect 1756 -772 1803 -738
rect 1403 -788 1803 -772
rect 1861 -738 2261 -700
rect 1861 -772 1908 -738
rect 1942 -772 1976 -738
rect 2010 -772 2044 -738
rect 2078 -772 2112 -738
rect 2146 -772 2180 -738
rect 2214 -772 2261 -738
rect 1861 -788 2261 -772
rect 2319 -738 2719 -700
rect 2319 -772 2366 -738
rect 2400 -772 2434 -738
rect 2468 -772 2502 -738
rect 2536 -772 2570 -738
rect 2604 -772 2638 -738
rect 2672 -772 2719 -738
rect 2319 -788 2719 -772
<< polycont >>
rect -2672 738 -2638 772
rect -2604 738 -2570 772
rect -2536 738 -2502 772
rect -2468 738 -2434 772
rect -2400 738 -2366 772
rect -2214 738 -2180 772
rect -2146 738 -2112 772
rect -2078 738 -2044 772
rect -2010 738 -1976 772
rect -1942 738 -1908 772
rect -1756 738 -1722 772
rect -1688 738 -1654 772
rect -1620 738 -1586 772
rect -1552 738 -1518 772
rect -1484 738 -1450 772
rect -1298 738 -1264 772
rect -1230 738 -1196 772
rect -1162 738 -1128 772
rect -1094 738 -1060 772
rect -1026 738 -992 772
rect -840 738 -806 772
rect -772 738 -738 772
rect -704 738 -670 772
rect -636 738 -602 772
rect -568 738 -534 772
rect -382 738 -348 772
rect -314 738 -280 772
rect -246 738 -212 772
rect -178 738 -144 772
rect -110 738 -76 772
rect 76 738 110 772
rect 144 738 178 772
rect 212 738 246 772
rect 280 738 314 772
rect 348 738 382 772
rect 534 738 568 772
rect 602 738 636 772
rect 670 738 704 772
rect 738 738 772 772
rect 806 738 840 772
rect 992 738 1026 772
rect 1060 738 1094 772
rect 1128 738 1162 772
rect 1196 738 1230 772
rect 1264 738 1298 772
rect 1450 738 1484 772
rect 1518 738 1552 772
rect 1586 738 1620 772
rect 1654 738 1688 772
rect 1722 738 1756 772
rect 1908 738 1942 772
rect 1976 738 2010 772
rect 2044 738 2078 772
rect 2112 738 2146 772
rect 2180 738 2214 772
rect 2366 738 2400 772
rect 2434 738 2468 772
rect 2502 738 2536 772
rect 2570 738 2604 772
rect 2638 738 2672 772
rect -2672 -772 -2638 -738
rect -2604 -772 -2570 -738
rect -2536 -772 -2502 -738
rect -2468 -772 -2434 -738
rect -2400 -772 -2366 -738
rect -2214 -772 -2180 -738
rect -2146 -772 -2112 -738
rect -2078 -772 -2044 -738
rect -2010 -772 -1976 -738
rect -1942 -772 -1908 -738
rect -1756 -772 -1722 -738
rect -1688 -772 -1654 -738
rect -1620 -772 -1586 -738
rect -1552 -772 -1518 -738
rect -1484 -772 -1450 -738
rect -1298 -772 -1264 -738
rect -1230 -772 -1196 -738
rect -1162 -772 -1128 -738
rect -1094 -772 -1060 -738
rect -1026 -772 -992 -738
rect -840 -772 -806 -738
rect -772 -772 -738 -738
rect -704 -772 -670 -738
rect -636 -772 -602 -738
rect -568 -772 -534 -738
rect -382 -772 -348 -738
rect -314 -772 -280 -738
rect -246 -772 -212 -738
rect -178 -772 -144 -738
rect -110 -772 -76 -738
rect 76 -772 110 -738
rect 144 -772 178 -738
rect 212 -772 246 -738
rect 280 -772 314 -738
rect 348 -772 382 -738
rect 534 -772 568 -738
rect 602 -772 636 -738
rect 670 -772 704 -738
rect 738 -772 772 -738
rect 806 -772 840 -738
rect 992 -772 1026 -738
rect 1060 -772 1094 -738
rect 1128 -772 1162 -738
rect 1196 -772 1230 -738
rect 1264 -772 1298 -738
rect 1450 -772 1484 -738
rect 1518 -772 1552 -738
rect 1586 -772 1620 -738
rect 1654 -772 1688 -738
rect 1722 -772 1756 -738
rect 1908 -772 1942 -738
rect 1976 -772 2010 -738
rect 2044 -772 2078 -738
rect 2112 -772 2146 -738
rect 2180 -772 2214 -738
rect 2366 -772 2400 -738
rect 2434 -772 2468 -738
rect 2502 -772 2536 -738
rect 2570 -772 2604 -738
rect 2638 -772 2672 -738
<< locali >>
rect -2879 840 -2771 874
rect -2737 840 -2703 874
rect -2669 840 -2635 874
rect -2601 840 -2567 874
rect -2533 840 -2499 874
rect -2465 840 -2431 874
rect -2397 840 -2363 874
rect -2329 840 -2295 874
rect -2261 840 -2227 874
rect -2193 840 -2159 874
rect -2125 840 -2091 874
rect -2057 840 -2023 874
rect -1989 840 -1955 874
rect -1921 840 -1887 874
rect -1853 840 -1819 874
rect -1785 840 -1751 874
rect -1717 840 -1683 874
rect -1649 840 -1615 874
rect -1581 840 -1547 874
rect -1513 840 -1479 874
rect -1445 840 -1411 874
rect -1377 840 -1343 874
rect -1309 840 -1275 874
rect -1241 840 -1207 874
rect -1173 840 -1139 874
rect -1105 840 -1071 874
rect -1037 840 -1003 874
rect -969 840 -935 874
rect -901 840 -867 874
rect -833 840 -799 874
rect -765 840 -731 874
rect -697 840 -663 874
rect -629 840 -595 874
rect -561 840 -527 874
rect -493 840 -459 874
rect -425 840 -391 874
rect -357 840 -323 874
rect -289 840 -255 874
rect -221 840 -187 874
rect -153 840 -119 874
rect -85 840 -51 874
rect -17 840 17 874
rect 51 840 85 874
rect 119 840 153 874
rect 187 840 221 874
rect 255 840 289 874
rect 323 840 357 874
rect 391 840 425 874
rect 459 840 493 874
rect 527 840 561 874
rect 595 840 629 874
rect 663 840 697 874
rect 731 840 765 874
rect 799 840 833 874
rect 867 840 901 874
rect 935 840 969 874
rect 1003 840 1037 874
rect 1071 840 1105 874
rect 1139 840 1173 874
rect 1207 840 1241 874
rect 1275 840 1309 874
rect 1343 840 1377 874
rect 1411 840 1445 874
rect 1479 840 1513 874
rect 1547 840 1581 874
rect 1615 840 1649 874
rect 1683 840 1717 874
rect 1751 840 1785 874
rect 1819 840 1853 874
rect 1887 840 1921 874
rect 1955 840 1989 874
rect 2023 840 2057 874
rect 2091 840 2125 874
rect 2159 840 2193 874
rect 2227 840 2261 874
rect 2295 840 2329 874
rect 2363 840 2397 874
rect 2431 840 2465 874
rect 2499 840 2533 874
rect 2567 840 2601 874
rect 2635 840 2669 874
rect 2703 840 2737 874
rect 2771 840 2879 874
rect -2879 765 -2845 840
rect -2719 738 -2672 772
rect -2638 738 -2604 772
rect -2570 738 -2536 772
rect -2502 738 -2468 772
rect -2434 738 -2400 772
rect -2366 738 -2319 772
rect -2261 738 -2214 772
rect -2180 738 -2146 772
rect -2112 738 -2078 772
rect -2044 738 -2010 772
rect -1976 738 -1942 772
rect -1908 738 -1861 772
rect -1803 738 -1756 772
rect -1722 738 -1688 772
rect -1654 738 -1620 772
rect -1586 738 -1552 772
rect -1518 738 -1484 772
rect -1450 738 -1403 772
rect -1345 738 -1298 772
rect -1264 738 -1230 772
rect -1196 738 -1162 772
rect -1128 738 -1094 772
rect -1060 738 -1026 772
rect -992 738 -945 772
rect -887 738 -840 772
rect -806 738 -772 772
rect -738 738 -704 772
rect -670 738 -636 772
rect -602 738 -568 772
rect -534 738 -487 772
rect -429 738 -382 772
rect -348 738 -314 772
rect -280 738 -246 772
rect -212 738 -178 772
rect -144 738 -110 772
rect -76 738 -29 772
rect 29 738 76 772
rect 110 738 144 772
rect 178 738 212 772
rect 246 738 280 772
rect 314 738 348 772
rect 382 738 429 772
rect 487 738 534 772
rect 568 738 602 772
rect 636 738 670 772
rect 704 738 738 772
rect 772 738 806 772
rect 840 738 887 772
rect 945 738 992 772
rect 1026 738 1060 772
rect 1094 738 1128 772
rect 1162 738 1196 772
rect 1230 738 1264 772
rect 1298 738 1345 772
rect 1403 738 1450 772
rect 1484 738 1518 772
rect 1552 738 1586 772
rect 1620 738 1654 772
rect 1688 738 1722 772
rect 1756 738 1803 772
rect 1861 738 1908 772
rect 1942 738 1976 772
rect 2010 738 2044 772
rect 2078 738 2112 772
rect 2146 738 2180 772
rect 2214 738 2261 772
rect 2319 738 2366 772
rect 2400 738 2434 772
rect 2468 738 2502 772
rect 2536 738 2570 772
rect 2604 738 2638 772
rect 2672 738 2719 772
rect 2845 765 2879 840
rect -2879 697 -2845 731
rect -2879 629 -2845 663
rect -2879 561 -2845 595
rect -2879 493 -2845 527
rect -2879 425 -2845 459
rect -2879 357 -2845 391
rect -2879 289 -2845 323
rect -2879 221 -2845 255
rect -2879 153 -2845 187
rect -2879 85 -2845 119
rect -2879 17 -2845 51
rect -2879 -51 -2845 -17
rect -2879 -119 -2845 -85
rect -2879 -187 -2845 -153
rect -2879 -255 -2845 -221
rect -2879 -323 -2845 -289
rect -2879 -391 -2845 -357
rect -2879 -459 -2845 -425
rect -2879 -527 -2845 -493
rect -2879 -595 -2845 -561
rect -2879 -663 -2845 -629
rect -2879 -731 -2845 -697
rect -2765 663 -2731 704
rect -2765 595 -2731 629
rect -2765 527 -2731 561
rect -2765 459 -2731 493
rect -2765 391 -2731 425
rect -2765 323 -2731 357
rect -2765 255 -2731 289
rect -2765 187 -2731 221
rect -2765 119 -2731 153
rect -2765 51 -2731 85
rect -2765 -17 -2731 17
rect -2765 -85 -2731 -51
rect -2765 -153 -2731 -119
rect -2765 -221 -2731 -187
rect -2765 -289 -2731 -255
rect -2765 -357 -2731 -323
rect -2765 -425 -2731 -391
rect -2765 -493 -2731 -459
rect -2765 -561 -2731 -527
rect -2765 -629 -2731 -595
rect -2765 -704 -2731 -663
rect -2307 663 -2273 704
rect -2307 595 -2273 629
rect -2307 527 -2273 561
rect -2307 459 -2273 493
rect -2307 391 -2273 425
rect -2307 323 -2273 357
rect -2307 255 -2273 289
rect -2307 187 -2273 221
rect -2307 119 -2273 153
rect -2307 51 -2273 85
rect -2307 -17 -2273 17
rect -2307 -85 -2273 -51
rect -2307 -153 -2273 -119
rect -2307 -221 -2273 -187
rect -2307 -289 -2273 -255
rect -2307 -357 -2273 -323
rect -2307 -425 -2273 -391
rect -2307 -493 -2273 -459
rect -2307 -561 -2273 -527
rect -2307 -629 -2273 -595
rect -2307 -704 -2273 -663
rect -1849 663 -1815 704
rect -1849 595 -1815 629
rect -1849 527 -1815 561
rect -1849 459 -1815 493
rect -1849 391 -1815 425
rect -1849 323 -1815 357
rect -1849 255 -1815 289
rect -1849 187 -1815 221
rect -1849 119 -1815 153
rect -1849 51 -1815 85
rect -1849 -17 -1815 17
rect -1849 -85 -1815 -51
rect -1849 -153 -1815 -119
rect -1849 -221 -1815 -187
rect -1849 -289 -1815 -255
rect -1849 -357 -1815 -323
rect -1849 -425 -1815 -391
rect -1849 -493 -1815 -459
rect -1849 -561 -1815 -527
rect -1849 -629 -1815 -595
rect -1849 -704 -1815 -663
rect -1391 663 -1357 704
rect -1391 595 -1357 629
rect -1391 527 -1357 561
rect -1391 459 -1357 493
rect -1391 391 -1357 425
rect -1391 323 -1357 357
rect -1391 255 -1357 289
rect -1391 187 -1357 221
rect -1391 119 -1357 153
rect -1391 51 -1357 85
rect -1391 -17 -1357 17
rect -1391 -85 -1357 -51
rect -1391 -153 -1357 -119
rect -1391 -221 -1357 -187
rect -1391 -289 -1357 -255
rect -1391 -357 -1357 -323
rect -1391 -425 -1357 -391
rect -1391 -493 -1357 -459
rect -1391 -561 -1357 -527
rect -1391 -629 -1357 -595
rect -1391 -704 -1357 -663
rect -933 663 -899 704
rect -933 595 -899 629
rect -933 527 -899 561
rect -933 459 -899 493
rect -933 391 -899 425
rect -933 323 -899 357
rect -933 255 -899 289
rect -933 187 -899 221
rect -933 119 -899 153
rect -933 51 -899 85
rect -933 -17 -899 17
rect -933 -85 -899 -51
rect -933 -153 -899 -119
rect -933 -221 -899 -187
rect -933 -289 -899 -255
rect -933 -357 -899 -323
rect -933 -425 -899 -391
rect -933 -493 -899 -459
rect -933 -561 -899 -527
rect -933 -629 -899 -595
rect -933 -704 -899 -663
rect -475 663 -441 704
rect -475 595 -441 629
rect -475 527 -441 561
rect -475 459 -441 493
rect -475 391 -441 425
rect -475 323 -441 357
rect -475 255 -441 289
rect -475 187 -441 221
rect -475 119 -441 153
rect -475 51 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -51
rect -475 -153 -441 -119
rect -475 -221 -441 -187
rect -475 -289 -441 -255
rect -475 -357 -441 -323
rect -475 -425 -441 -391
rect -475 -493 -441 -459
rect -475 -561 -441 -527
rect -475 -629 -441 -595
rect -475 -704 -441 -663
rect -17 663 17 704
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -704 17 -663
rect 441 663 475 704
rect 441 595 475 629
rect 441 527 475 561
rect 441 459 475 493
rect 441 391 475 425
rect 441 323 475 357
rect 441 255 475 289
rect 441 187 475 221
rect 441 119 475 153
rect 441 51 475 85
rect 441 -17 475 17
rect 441 -85 475 -51
rect 441 -153 475 -119
rect 441 -221 475 -187
rect 441 -289 475 -255
rect 441 -357 475 -323
rect 441 -425 475 -391
rect 441 -493 475 -459
rect 441 -561 475 -527
rect 441 -629 475 -595
rect 441 -704 475 -663
rect 899 663 933 704
rect 899 595 933 629
rect 899 527 933 561
rect 899 459 933 493
rect 899 391 933 425
rect 899 323 933 357
rect 899 255 933 289
rect 899 187 933 221
rect 899 119 933 153
rect 899 51 933 85
rect 899 -17 933 17
rect 899 -85 933 -51
rect 899 -153 933 -119
rect 899 -221 933 -187
rect 899 -289 933 -255
rect 899 -357 933 -323
rect 899 -425 933 -391
rect 899 -493 933 -459
rect 899 -561 933 -527
rect 899 -629 933 -595
rect 899 -704 933 -663
rect 1357 663 1391 704
rect 1357 595 1391 629
rect 1357 527 1391 561
rect 1357 459 1391 493
rect 1357 391 1391 425
rect 1357 323 1391 357
rect 1357 255 1391 289
rect 1357 187 1391 221
rect 1357 119 1391 153
rect 1357 51 1391 85
rect 1357 -17 1391 17
rect 1357 -85 1391 -51
rect 1357 -153 1391 -119
rect 1357 -221 1391 -187
rect 1357 -289 1391 -255
rect 1357 -357 1391 -323
rect 1357 -425 1391 -391
rect 1357 -493 1391 -459
rect 1357 -561 1391 -527
rect 1357 -629 1391 -595
rect 1357 -704 1391 -663
rect 1815 663 1849 704
rect 1815 595 1849 629
rect 1815 527 1849 561
rect 1815 459 1849 493
rect 1815 391 1849 425
rect 1815 323 1849 357
rect 1815 255 1849 289
rect 1815 187 1849 221
rect 1815 119 1849 153
rect 1815 51 1849 85
rect 1815 -17 1849 17
rect 1815 -85 1849 -51
rect 1815 -153 1849 -119
rect 1815 -221 1849 -187
rect 1815 -289 1849 -255
rect 1815 -357 1849 -323
rect 1815 -425 1849 -391
rect 1815 -493 1849 -459
rect 1815 -561 1849 -527
rect 1815 -629 1849 -595
rect 1815 -704 1849 -663
rect 2273 663 2307 704
rect 2273 595 2307 629
rect 2273 527 2307 561
rect 2273 459 2307 493
rect 2273 391 2307 425
rect 2273 323 2307 357
rect 2273 255 2307 289
rect 2273 187 2307 221
rect 2273 119 2307 153
rect 2273 51 2307 85
rect 2273 -17 2307 17
rect 2273 -85 2307 -51
rect 2273 -153 2307 -119
rect 2273 -221 2307 -187
rect 2273 -289 2307 -255
rect 2273 -357 2307 -323
rect 2273 -425 2307 -391
rect 2273 -493 2307 -459
rect 2273 -561 2307 -527
rect 2273 -629 2307 -595
rect 2273 -704 2307 -663
rect 2731 663 2765 704
rect 2731 595 2765 629
rect 2731 527 2765 561
rect 2731 459 2765 493
rect 2731 391 2765 425
rect 2731 323 2765 357
rect 2731 255 2765 289
rect 2731 187 2765 221
rect 2731 119 2765 153
rect 2731 51 2765 85
rect 2731 -17 2765 17
rect 2731 -85 2765 -51
rect 2731 -153 2765 -119
rect 2731 -221 2765 -187
rect 2731 -289 2765 -255
rect 2731 -357 2765 -323
rect 2731 -425 2765 -391
rect 2731 -493 2765 -459
rect 2731 -561 2765 -527
rect 2731 -629 2765 -595
rect 2731 -704 2765 -663
rect 2845 697 2879 731
rect 2845 629 2879 663
rect 2845 561 2879 595
rect 2845 493 2879 527
rect 2845 425 2879 459
rect 2845 357 2879 391
rect 2845 289 2879 323
rect 2845 221 2879 255
rect 2845 153 2879 187
rect 2845 85 2879 119
rect 2845 17 2879 51
rect 2845 -51 2879 -17
rect 2845 -119 2879 -85
rect 2845 -187 2879 -153
rect 2845 -255 2879 -221
rect 2845 -323 2879 -289
rect 2845 -391 2879 -357
rect 2845 -459 2879 -425
rect 2845 -527 2879 -493
rect 2845 -595 2879 -561
rect 2845 -663 2879 -629
rect 2845 -731 2879 -697
rect -2879 -840 -2845 -765
rect -2719 -772 -2672 -738
rect -2638 -772 -2604 -738
rect -2570 -772 -2536 -738
rect -2502 -772 -2468 -738
rect -2434 -772 -2400 -738
rect -2366 -772 -2319 -738
rect -2261 -772 -2214 -738
rect -2180 -772 -2146 -738
rect -2112 -772 -2078 -738
rect -2044 -772 -2010 -738
rect -1976 -772 -1942 -738
rect -1908 -772 -1861 -738
rect -1803 -772 -1756 -738
rect -1722 -772 -1688 -738
rect -1654 -772 -1620 -738
rect -1586 -772 -1552 -738
rect -1518 -772 -1484 -738
rect -1450 -772 -1403 -738
rect -1345 -772 -1298 -738
rect -1264 -772 -1230 -738
rect -1196 -772 -1162 -738
rect -1128 -772 -1094 -738
rect -1060 -772 -1026 -738
rect -992 -772 -945 -738
rect -887 -772 -840 -738
rect -806 -772 -772 -738
rect -738 -772 -704 -738
rect -670 -772 -636 -738
rect -602 -772 -568 -738
rect -534 -772 -487 -738
rect -429 -772 -382 -738
rect -348 -772 -314 -738
rect -280 -772 -246 -738
rect -212 -772 -178 -738
rect -144 -772 -110 -738
rect -76 -772 -29 -738
rect 29 -772 76 -738
rect 110 -772 144 -738
rect 178 -772 212 -738
rect 246 -772 280 -738
rect 314 -772 348 -738
rect 382 -772 429 -738
rect 487 -772 534 -738
rect 568 -772 602 -738
rect 636 -772 670 -738
rect 704 -772 738 -738
rect 772 -772 806 -738
rect 840 -772 887 -738
rect 945 -772 992 -738
rect 1026 -772 1060 -738
rect 1094 -772 1128 -738
rect 1162 -772 1196 -738
rect 1230 -772 1264 -738
rect 1298 -772 1345 -738
rect 1403 -772 1450 -738
rect 1484 -772 1518 -738
rect 1552 -772 1586 -738
rect 1620 -772 1654 -738
rect 1688 -772 1722 -738
rect 1756 -772 1803 -738
rect 1861 -772 1908 -738
rect 1942 -772 1976 -738
rect 2010 -772 2044 -738
rect 2078 -772 2112 -738
rect 2146 -772 2180 -738
rect 2214 -772 2261 -738
rect 2319 -772 2366 -738
rect 2400 -772 2434 -738
rect 2468 -772 2502 -738
rect 2536 -772 2570 -738
rect 2604 -772 2638 -738
rect 2672 -772 2719 -738
rect 2845 -840 2879 -765
rect -2879 -874 -2771 -840
rect -2737 -874 -2703 -840
rect -2669 -874 -2635 -840
rect -2601 -874 -2567 -840
rect -2533 -874 -2499 -840
rect -2465 -874 -2431 -840
rect -2397 -874 -2363 -840
rect -2329 -874 -2295 -840
rect -2261 -874 -2227 -840
rect -2193 -874 -2159 -840
rect -2125 -874 -2091 -840
rect -2057 -874 -2023 -840
rect -1989 -874 -1955 -840
rect -1921 -874 -1887 -840
rect -1853 -874 -1819 -840
rect -1785 -874 -1751 -840
rect -1717 -874 -1683 -840
rect -1649 -874 -1615 -840
rect -1581 -874 -1547 -840
rect -1513 -874 -1479 -840
rect -1445 -874 -1411 -840
rect -1377 -874 -1343 -840
rect -1309 -874 -1275 -840
rect -1241 -874 -1207 -840
rect -1173 -874 -1139 -840
rect -1105 -874 -1071 -840
rect -1037 -874 -1003 -840
rect -969 -874 -935 -840
rect -901 -874 -867 -840
rect -833 -874 -799 -840
rect -765 -874 -731 -840
rect -697 -874 -663 -840
rect -629 -874 -595 -840
rect -561 -874 -527 -840
rect -493 -874 -459 -840
rect -425 -874 -391 -840
rect -357 -874 -323 -840
rect -289 -874 -255 -840
rect -221 -874 -187 -840
rect -153 -874 -119 -840
rect -85 -874 -51 -840
rect -17 -874 17 -840
rect 51 -874 85 -840
rect 119 -874 153 -840
rect 187 -874 221 -840
rect 255 -874 289 -840
rect 323 -874 357 -840
rect 391 -874 425 -840
rect 459 -874 493 -840
rect 527 -874 561 -840
rect 595 -874 629 -840
rect 663 -874 697 -840
rect 731 -874 765 -840
rect 799 -874 833 -840
rect 867 -874 901 -840
rect 935 -874 969 -840
rect 1003 -874 1037 -840
rect 1071 -874 1105 -840
rect 1139 -874 1173 -840
rect 1207 -874 1241 -840
rect 1275 -874 1309 -840
rect 1343 -874 1377 -840
rect 1411 -874 1445 -840
rect 1479 -874 1513 -840
rect 1547 -874 1581 -840
rect 1615 -874 1649 -840
rect 1683 -874 1717 -840
rect 1751 -874 1785 -840
rect 1819 -874 1853 -840
rect 1887 -874 1921 -840
rect 1955 -874 1989 -840
rect 2023 -874 2057 -840
rect 2091 -874 2125 -840
rect 2159 -874 2193 -840
rect 2227 -874 2261 -840
rect 2295 -874 2329 -840
rect 2363 -874 2397 -840
rect 2431 -874 2465 -840
rect 2499 -874 2533 -840
rect 2567 -874 2601 -840
rect 2635 -874 2669 -840
rect 2703 -874 2737 -840
rect 2771 -874 2879 -840
<< properties >>
string FIXED_BBOX -2862 -857 2862 857
<< end >>
