magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect 5184 2660 5398 2676
rect -152 2404 5398 2660
rect -152 2384 5370 2404
<< nsubdiff >>
rect -84 2547 5344 2612
rect -84 2513 209 2547
rect 243 2543 1223 2547
rect 243 2513 517 2543
rect -84 2509 517 2513
rect 551 2509 859 2543
rect 893 2513 1223 2543
rect 1257 2543 1953 2547
rect 1257 2513 1575 2543
rect 893 2509 1575 2513
rect 1609 2513 1953 2543
rect 1987 2543 2647 2547
rect 1987 2513 2273 2543
rect 1609 2509 2273 2513
rect 2307 2513 2647 2543
rect 2681 2513 2993 2547
rect 3027 2543 4861 2547
rect 3027 2537 4371 2543
rect 3027 2513 3709 2537
rect 2307 2509 3709 2513
rect -84 2503 3709 2509
rect 3743 2509 4371 2537
rect 4405 2513 4861 2543
rect 4895 2513 5344 2547
rect 4405 2509 5344 2513
rect 3743 2503 5344 2509
rect -84 2452 5344 2503
<< nsubdiffcont >>
rect 209 2513 243 2547
rect 517 2509 551 2543
rect 859 2509 893 2543
rect 1223 2513 1257 2547
rect 1575 2509 1609 2543
rect 1953 2513 1987 2547
rect 2273 2509 2307 2543
rect 2647 2513 2681 2547
rect 2993 2513 3027 2547
rect 3709 2503 3743 2537
rect 4371 2509 4405 2543
rect 4861 2513 4895 2547
<< locali >>
rect 3882 2576 3966 2580
rect -20 2560 5316 2576
rect -20 2554 3907 2560
rect -20 2550 1771 2554
rect -20 2547 369 2550
rect -20 2544 209 2547
rect -20 2510 81 2544
rect 115 2513 209 2544
rect 243 2516 369 2547
rect 403 2543 693 2550
rect 403 2516 517 2543
rect 243 2513 517 2516
rect 115 2510 517 2513
rect -20 2509 517 2510
rect 551 2516 693 2543
rect 727 2543 1041 2550
rect 727 2516 859 2543
rect 551 2509 859 2516
rect 893 2516 1041 2543
rect 1075 2547 1415 2550
rect 1075 2516 1223 2547
rect 893 2513 1223 2516
rect 1257 2516 1415 2547
rect 1449 2543 1771 2550
rect 1449 2516 1575 2543
rect 1257 2513 1575 2516
rect 893 2509 1575 2513
rect 1609 2520 1771 2543
rect 1805 2550 2829 2554
rect 1805 2547 2509 2550
rect 1805 2520 1953 2547
rect 1609 2513 1953 2520
rect 1987 2544 2509 2547
rect 1987 2513 2087 2544
rect 1609 2510 2087 2513
rect 2121 2543 2509 2544
rect 2121 2510 2273 2543
rect 1609 2509 2273 2510
rect 2307 2516 2509 2543
rect 2543 2547 2829 2550
rect 2543 2516 2647 2547
rect 2307 2513 2647 2516
rect 2681 2520 2829 2547
rect 2863 2550 3907 2554
rect 2863 2547 3143 2550
rect 2863 2520 2993 2547
rect 2681 2513 2993 2520
rect 3027 2516 3143 2547
rect 3177 2516 3495 2550
rect 3529 2537 3907 2550
rect 3529 2516 3709 2537
rect 3027 2513 3709 2516
rect 2307 2509 3709 2513
rect -20 2503 3709 2509
rect 3743 2526 3907 2537
rect 3941 2554 5316 2560
rect 3941 2550 4745 2554
rect 3941 2526 4237 2550
rect 3743 2516 4237 2526
rect 4271 2543 4477 2550
rect 4271 2516 4371 2543
rect 3743 2509 4371 2516
rect 4405 2516 4477 2543
rect 4511 2520 4745 2550
rect 4779 2550 5316 2554
rect 4779 2547 4969 2550
rect 4779 2520 4861 2547
rect 4511 2516 4861 2520
rect 4405 2513 4861 2516
rect 4895 2516 4969 2547
rect 5003 2516 5316 2550
rect 4895 2513 5316 2516
rect 4405 2509 5316 2513
rect 3743 2503 5316 2509
rect -20 2474 5316 2503
rect 1204 2470 3808 2474
rect 1204 2314 1264 2470
rect 3746 2322 3806 2470
rect 159 2213 176 2247
rect 210 2213 227 2247
rect 317 2213 334 2247
rect 368 2213 385 2247
rect 475 2213 492 2247
rect 526 2213 543 2247
rect 633 2213 650 2247
rect 684 2213 701 2247
rect 791 2213 808 2247
rect 842 2213 859 2247
rect 949 2213 966 2247
rect 1000 2213 1017 2247
rect 1107 2213 1124 2247
rect 1158 2213 1175 2247
rect 1265 2213 1282 2247
rect 1316 2213 1333 2247
rect 1423 2213 1440 2247
rect 1474 2213 1491 2247
rect 1581 2213 1598 2247
rect 1632 2213 1649 2247
rect 1739 2213 1756 2247
rect 1790 2213 1807 2247
rect 1897 2213 1914 2247
rect 1948 2213 1965 2247
rect 2055 2213 2072 2247
rect 2106 2213 2123 2247
rect 2213 2213 2230 2247
rect 2264 2213 2281 2247
rect 2371 2213 2388 2247
rect 2422 2213 2439 2247
rect 2860 2218 2877 2252
rect 2911 2218 2928 2252
rect 3018 2218 3035 2252
rect 3069 2218 3086 2252
rect 3176 2218 3193 2252
rect 3227 2218 3244 2252
rect 3334 2218 3351 2252
rect 3385 2218 3402 2252
rect 3492 2218 3509 2252
rect 3543 2218 3560 2252
rect 3650 2218 3667 2252
rect 3701 2218 3718 2252
rect 3808 2218 3825 2252
rect 3859 2218 3876 2252
rect 3966 2218 3983 2252
rect 4017 2218 4034 2252
rect 4124 2218 4141 2252
rect 4175 2218 4192 2252
rect 4282 2218 4299 2252
rect 4333 2218 4350 2252
rect 4440 2218 4457 2252
rect 4491 2218 4508 2252
rect 4598 2218 4615 2252
rect 4649 2218 4666 2252
rect 4756 2218 4773 2252
rect 4807 2218 4824 2252
rect 4914 2218 4931 2252
rect 4965 2218 4982 2252
rect 5072 2218 5089 2252
rect 5123 2218 5140 2252
rect 98 2052 136 2070
rect 98 2018 100 2052
rect 134 2018 136 2052
rect 98 2000 136 2018
rect 414 2060 452 2078
rect 414 2026 416 2060
rect 450 2026 452 2060
rect 414 2008 452 2026
rect 726 2060 764 2078
rect 726 2026 728 2060
rect 762 2026 764 2060
rect 726 2008 764 2026
rect 1044 2066 1082 2084
rect 1044 2032 1046 2066
rect 1080 2032 1082 2066
rect 1044 2014 1082 2032
rect 1358 2058 1396 2076
rect 1358 2024 1360 2058
rect 1394 2024 1396 2058
rect 1358 2006 1396 2024
rect 1676 2054 1714 2072
rect 1676 2020 1678 2054
rect 1712 2020 1714 2054
rect 1676 2002 1714 2020
rect 1992 2060 2030 2078
rect 1992 2026 1994 2060
rect 2028 2026 2030 2060
rect 1992 2008 2030 2026
rect 2308 2064 2346 2082
rect 2308 2030 2310 2064
rect 2344 2030 2346 2064
rect 2308 2012 2346 2030
rect 2796 2026 2832 2060
rect 2796 1992 2797 2026
rect 2831 1992 2832 2026
rect 2796 1958 2832 1992
rect 3110 2040 3146 2074
rect 3110 2006 3111 2040
rect 3145 2006 3146 2040
rect 3110 1972 3146 2006
rect 3270 2004 3304 2088
rect 3428 2040 3464 2074
rect 3428 2006 3429 2040
rect 3463 2006 3464 2040
rect 3586 2012 3620 2096
rect 3746 2036 3782 2070
rect 3428 1972 3464 2006
rect 3746 2002 3747 2036
rect 3781 2002 3782 2036
rect 3902 2016 3936 2100
rect 4058 2042 4094 2076
rect 3746 1968 3782 2002
rect 4058 2008 4059 2042
rect 4093 2008 4094 2042
rect 4058 1974 4094 2008
rect 4374 2044 4410 2078
rect 4374 2010 4375 2044
rect 4409 2010 4410 2044
rect 4374 1976 4410 2010
rect 4690 2036 4726 2070
rect 4690 2002 4691 2036
rect 4725 2002 4726 2036
rect 4690 1968 4726 2002
rect 5012 2040 5048 2074
rect 5012 2006 5013 2040
rect 5047 2006 5048 2040
rect 5012 1972 5048 2006
rect 3268 1857 3302 1858
rect 2956 1849 2990 1850
rect 252 1798 290 1816
rect 252 1764 254 1798
rect 288 1764 290 1798
rect 252 1746 290 1764
rect 566 1802 604 1820
rect 566 1768 568 1802
rect 602 1768 604 1802
rect 566 1750 604 1768
rect 888 1800 926 1818
rect 888 1766 890 1800
rect 924 1766 926 1800
rect 888 1748 926 1766
rect 1204 1804 1242 1822
rect 1204 1770 1206 1804
rect 1240 1770 1242 1804
rect 1204 1752 1242 1770
rect 1522 1808 1560 1826
rect 1522 1774 1524 1808
rect 1558 1774 1560 1808
rect 1522 1756 1560 1774
rect 1834 1808 1872 1826
rect 1834 1774 1836 1808
rect 1870 1774 1872 1808
rect 1834 1756 1872 1774
rect 2156 1808 2194 1826
rect 2156 1774 2158 1808
rect 2192 1774 2194 1808
rect 2156 1756 2194 1774
rect 2466 1804 2504 1822
rect 2466 1770 2468 1804
rect 2502 1770 2504 1804
rect 2466 1752 2504 1770
rect 2956 1777 2990 1815
rect 3902 1855 3936 1856
rect 3268 1785 3302 1823
rect 3268 1750 3302 1751
rect 3586 1853 3620 1854
rect 3586 1781 3620 1819
rect 3902 1783 3936 1821
rect 3902 1748 3936 1749
rect 4222 1855 4256 1856
rect 4222 1783 4256 1821
rect 4222 1748 4256 1749
rect 4536 1849 4570 1850
rect 4536 1777 4570 1815
rect 3586 1746 3620 1747
rect 2956 1742 2990 1743
rect 4536 1742 4570 1743
rect 4852 1849 4886 1850
rect 4852 1777 4886 1815
rect 4852 1742 4886 1743
rect 5168 1849 5202 1850
rect 5168 1777 5202 1815
rect 5168 1742 5202 1743
rect 2371 85 2388 119
rect 2422 85 2439 119
rect 2274 -412 2342 -396
rect 2392 -402 2405 -368
rect 2439 -402 2452 -368
rect 2894 -404 2907 -370
rect 2941 -404 2954 -370
rect 2274 -446 2289 -412
rect 2323 -446 2342 -412
rect 2274 -462 2342 -446
rect 3004 -414 3072 -398
rect 3004 -448 3029 -414
rect 3063 -448 3072 -414
rect 2392 -490 2405 -456
rect 2439 -490 2452 -456
rect 2894 -492 2907 -458
rect 2941 -492 2954 -458
rect 3004 -464 3072 -448
rect 2396 -602 2412 -568
rect 2446 -602 2462 -568
rect 2892 -606 2908 -572
rect 2942 -606 2958 -572
rect 2642 -1016 2648 -982
rect 2682 -1016 2688 -982
rect 1372 -1067 1406 -1044
rect 1372 -1139 1406 -1101
rect 1372 -1211 1406 -1173
rect 1372 -1283 1406 -1245
rect 1372 -1355 1406 -1317
rect 1372 -1412 1406 -1389
rect 1456 -1474 1463 -1440
rect 1497 -1474 1535 -1440
rect 1569 -1474 1607 -1440
rect 1641 -1474 1679 -1440
rect 1713 -1474 1751 -1440
rect 1785 -1474 1823 -1440
rect 1857 -1474 1895 -1440
rect 1929 -1474 1967 -1440
rect 2001 -1474 2039 -1440
rect 2073 -1474 2111 -1440
rect 2145 -1474 2183 -1440
rect 2217 -1474 2255 -1440
rect 2289 -1474 2327 -1440
rect 2361 -1474 2399 -1440
rect 2433 -1474 2471 -1440
rect 2505 -1474 2543 -1440
rect 2577 -1474 2615 -1440
rect 2649 -1474 2687 -1440
rect 2721 -1474 2759 -1440
rect 2793 -1474 2831 -1440
rect 2865 -1474 2903 -1440
rect 2937 -1474 2975 -1440
rect 3009 -1474 3047 -1440
rect 3081 -1474 3119 -1440
rect 3153 -1474 3191 -1440
rect 3225 -1474 3263 -1440
rect 3297 -1474 3335 -1440
rect 3369 -1474 3407 -1440
rect 3441 -1474 3479 -1440
rect 3513 -1474 3551 -1440
rect 3585 -1474 3623 -1440
rect 3657 -1474 3695 -1440
rect 3729 -1474 3767 -1440
rect 3801 -1474 3839 -1440
rect 3873 -1474 3911 -1440
rect 3945 -1474 3952 -1440
rect 1478 -1586 1487 -1552
rect 1521 -1586 1530 -1552
rect 1810 -1592 1819 -1558
rect 1853 -1592 1862 -1558
rect 2292 -1592 2301 -1558
rect 2335 -1592 2344 -1558
rect 2944 -1586 2953 -1552
rect 2987 -1586 2996 -1552
rect 3530 -1590 3539 -1556
rect 3573 -1590 3582 -1556
rect 3848 -1588 3857 -1554
rect 3891 -1588 3900 -1554
<< viali >>
rect 81 2510 115 2544
rect 369 2516 403 2550
rect 693 2516 727 2550
rect 1041 2516 1075 2550
rect 1415 2516 1449 2550
rect 1771 2520 1805 2554
rect 2087 2510 2121 2544
rect 2509 2516 2543 2550
rect 2829 2520 2863 2554
rect 3143 2516 3177 2550
rect 3495 2516 3529 2550
rect 3907 2526 3941 2560
rect 4237 2516 4271 2550
rect 4477 2516 4511 2550
rect 4745 2520 4779 2554
rect 4969 2516 5003 2550
rect 176 2213 210 2247
rect 334 2213 368 2247
rect 492 2213 526 2247
rect 650 2213 684 2247
rect 808 2213 842 2247
rect 966 2213 1000 2247
rect 1124 2213 1158 2247
rect 1282 2213 1316 2247
rect 1440 2213 1474 2247
rect 1598 2213 1632 2247
rect 1756 2213 1790 2247
rect 1914 2213 1948 2247
rect 2072 2213 2106 2247
rect 2230 2213 2264 2247
rect 2388 2213 2422 2247
rect 2877 2218 2911 2252
rect 3035 2218 3069 2252
rect 3193 2218 3227 2252
rect 3351 2218 3385 2252
rect 3509 2218 3543 2252
rect 3667 2218 3701 2252
rect 3825 2218 3859 2252
rect 3983 2218 4017 2252
rect 4141 2218 4175 2252
rect 4299 2218 4333 2252
rect 4457 2218 4491 2252
rect 4615 2218 4649 2252
rect 4773 2218 4807 2252
rect 4931 2218 4965 2252
rect 5089 2218 5123 2252
rect 100 2018 134 2052
rect 416 2026 450 2060
rect 728 2026 762 2060
rect 1046 2032 1080 2066
rect 1360 2024 1394 2058
rect 1678 2020 1712 2054
rect 1994 2026 2028 2060
rect 2310 2030 2344 2064
rect 2797 1992 2831 2026
rect 3111 2006 3145 2040
rect 3429 2006 3463 2040
rect 3747 2002 3781 2036
rect 4059 2008 4093 2042
rect 4375 2010 4409 2044
rect 4691 2002 4725 2036
rect 5013 2006 5047 2040
rect 254 1764 288 1798
rect 568 1768 602 1802
rect 890 1766 924 1800
rect 1206 1770 1240 1804
rect 1524 1774 1558 1808
rect 1836 1774 1870 1808
rect 2158 1774 2192 1808
rect 2468 1770 2502 1804
rect 2956 1815 2990 1849
rect 2956 1743 2990 1777
rect 3268 1823 3302 1857
rect 3268 1751 3302 1785
rect 3586 1819 3620 1853
rect 3586 1747 3620 1781
rect 3902 1821 3936 1855
rect 3902 1749 3936 1783
rect 4222 1821 4256 1855
rect 4222 1749 4256 1783
rect 4536 1815 4570 1849
rect 4536 1743 4570 1777
rect 4852 1815 4886 1849
rect 4852 1743 4886 1777
rect 5168 1815 5202 1849
rect 5168 1743 5202 1777
rect 2388 85 2422 119
rect 2405 -402 2439 -368
rect 2907 -404 2941 -370
rect 2289 -446 2323 -412
rect 3029 -448 3063 -414
rect 2405 -490 2439 -456
rect 2907 -492 2941 -458
rect 2412 -602 2446 -568
rect 2908 -606 2942 -572
rect 2648 -1016 2682 -982
rect 1372 -1101 1406 -1067
rect 1372 -1173 1406 -1139
rect 1372 -1245 1406 -1211
rect 1372 -1317 1406 -1283
rect 1372 -1389 1406 -1355
rect 1463 -1474 1497 -1440
rect 1535 -1474 1569 -1440
rect 1607 -1474 1641 -1440
rect 1679 -1474 1713 -1440
rect 1751 -1474 1785 -1440
rect 1823 -1474 1857 -1440
rect 1895 -1474 1929 -1440
rect 1967 -1474 2001 -1440
rect 2039 -1474 2073 -1440
rect 2111 -1474 2145 -1440
rect 2183 -1474 2217 -1440
rect 2255 -1474 2289 -1440
rect 2327 -1474 2361 -1440
rect 2399 -1474 2433 -1440
rect 2471 -1474 2505 -1440
rect 2543 -1474 2577 -1440
rect 2615 -1474 2649 -1440
rect 2687 -1474 2721 -1440
rect 2759 -1474 2793 -1440
rect 2831 -1474 2865 -1440
rect 2903 -1474 2937 -1440
rect 2975 -1474 3009 -1440
rect 3047 -1474 3081 -1440
rect 3119 -1474 3153 -1440
rect 3191 -1474 3225 -1440
rect 3263 -1474 3297 -1440
rect 3335 -1474 3369 -1440
rect 3407 -1474 3441 -1440
rect 3479 -1474 3513 -1440
rect 3551 -1474 3585 -1440
rect 3623 -1474 3657 -1440
rect 3695 -1474 3729 -1440
rect 3767 -1474 3801 -1440
rect 3839 -1474 3873 -1440
rect 3911 -1474 3945 -1440
rect 1487 -1586 1521 -1552
rect 1819 -1592 1853 -1558
rect 2301 -1592 2335 -1558
rect 2953 -1586 2987 -1552
rect 3539 -1590 3573 -1556
rect 3857 -1588 3891 -1554
<< metal1 >>
rect 1739 4741 3642 4973
rect 1739 3473 1988 4741
rect 3384 3473 3642 4741
rect 1739 3396 3642 3473
rect -122 2583 5343 3396
rect -122 2544 93 2583
rect 145 2560 5343 2583
rect 145 2554 3907 2560
rect 145 2550 1771 2554
rect -122 2510 81 2544
rect 145 2531 369 2550
rect 115 2519 369 2531
rect 145 2516 369 2519
rect 403 2516 693 2550
rect 727 2516 1041 2550
rect 1075 2516 1415 2550
rect 1449 2520 1771 2550
rect 1805 2550 2829 2554
rect 1805 2544 2509 2550
rect 1805 2520 2087 2544
rect 1449 2516 2087 2520
rect 145 2510 2087 2516
rect 2121 2516 2509 2544
rect 2543 2520 2829 2550
rect 2863 2550 3907 2554
rect 2863 2520 3143 2550
rect 2543 2516 3143 2520
rect 3177 2516 3495 2550
rect 3529 2526 3907 2550
rect 3941 2554 5343 2560
rect 3941 2550 4745 2554
rect 3941 2526 4237 2550
rect 3529 2516 4237 2526
rect 4271 2516 4477 2550
rect 4511 2520 4745 2550
rect 4779 2550 5343 2554
rect 4779 2520 4969 2550
rect 4511 2516 4969 2520
rect 5003 2546 5343 2550
rect 5003 2516 5157 2546
rect 2121 2510 5157 2516
rect -122 2467 93 2510
rect 145 2494 5157 2510
rect 5209 2494 5343 2546
rect 145 2467 5343 2494
rect -122 2437 5343 2467
rect -110 2436 5338 2437
rect 2830 2274 5170 2278
rect 132 2252 5170 2274
rect 132 2247 2877 2252
rect 132 2213 176 2247
rect 210 2213 334 2247
rect 368 2213 492 2247
rect 526 2213 650 2247
rect 684 2213 808 2247
rect 842 2213 966 2247
rect 1000 2213 1124 2247
rect 1158 2213 1282 2247
rect 1316 2213 1440 2247
rect 1474 2213 1598 2247
rect 1632 2213 1756 2247
rect 1790 2213 1914 2247
rect 1948 2213 2072 2247
rect 2106 2213 2230 2247
rect 2264 2213 2388 2247
rect 2422 2218 2877 2247
rect 2911 2218 3035 2252
rect 3069 2218 3193 2252
rect 3227 2218 3351 2252
rect 3385 2218 3509 2252
rect 3543 2218 3667 2252
rect 3701 2218 3825 2252
rect 3859 2218 3983 2252
rect 4017 2218 4141 2252
rect 4175 2218 4299 2252
rect 4333 2218 4457 2252
rect 4491 2218 4615 2252
rect 4649 2218 4773 2252
rect 4807 2218 4931 2252
rect 4965 2218 5089 2252
rect 5123 2218 5170 2252
rect 2422 2213 5170 2218
rect 132 2200 5170 2213
rect 2350 2196 3320 2200
rect 26 2110 234 2124
rect 26 2103 2356 2110
rect 26 2051 93 2103
rect 145 2066 2356 2103
rect 145 2060 1046 2066
rect 145 2051 416 2060
rect 26 2039 100 2051
rect 134 2039 416 2051
rect 26 1987 93 2039
rect 145 2026 416 2039
rect 450 2026 728 2060
rect 762 2032 1046 2060
rect 1080 2064 2356 2066
rect 1080 2060 2310 2064
rect 1080 2058 1994 2060
rect 1080 2032 1360 2058
rect 762 2026 1360 2032
rect 145 2024 1360 2026
rect 1394 2054 1994 2058
rect 1394 2024 1678 2054
rect 145 2020 1678 2024
rect 1712 2026 1994 2054
rect 2028 2030 2310 2060
rect 2344 2030 2356 2064
rect 2028 2026 2356 2030
rect 1712 2020 2356 2026
rect 145 1987 2356 2020
rect 26 1962 2356 1987
rect 26 1944 234 1962
rect 2750 2084 2874 2086
rect 2750 2044 5062 2084
rect 2750 2042 4375 2044
rect 2750 2040 4059 2042
rect 2750 2026 3111 2040
rect 2750 1992 2797 2026
rect 2831 2006 3111 2026
rect 3145 2006 3429 2040
rect 3463 2036 4059 2040
rect 3463 2006 3747 2036
rect 2831 2002 3747 2006
rect 3781 2008 4059 2036
rect 4093 2010 4375 2042
rect 4409 2040 5062 2044
rect 4409 2036 5013 2040
rect 4409 2010 4691 2036
rect 4093 2008 4691 2010
rect 3781 2002 4691 2008
rect 4725 2006 5013 2036
rect 5047 2006 5062 2040
rect 4725 2002 5062 2006
rect 2831 1992 5062 2002
rect 2750 1950 5062 1992
rect 2426 1864 2546 1870
rect 238 1808 2546 1864
rect 2750 1832 2874 1950
rect 5108 1864 5260 1878
rect 238 1804 1524 1808
rect 238 1802 1206 1804
rect 238 1798 568 1802
rect 238 1764 254 1798
rect 288 1768 568 1798
rect 602 1800 1206 1802
rect 602 1768 890 1800
rect 288 1766 890 1768
rect 924 1770 1206 1800
rect 1240 1774 1524 1804
rect 1558 1774 1836 1808
rect 1870 1774 2158 1808
rect 2192 1804 2546 1808
rect 2192 1774 2468 1804
rect 1240 1770 2468 1774
rect 2502 1770 2546 1804
rect 924 1766 2546 1770
rect 288 1764 2546 1766
rect 238 1700 2546 1764
rect -631 42 -269 190
rect 2426 134 2546 1700
rect 2352 119 2546 134
rect 2352 85 2388 119
rect 2422 85 2546 119
rect 2352 64 2546 85
rect -631 -74 -495 42
rect -379 -74 -269 42
rect -631 -119 -269 -74
rect 2426 -119 2546 64
rect -631 -196 2546 -119
rect 2738 62 2874 1832
rect 2944 1857 5260 1864
rect 2944 1849 3268 1857
rect 2944 1815 2956 1849
rect 2990 1823 3268 1849
rect 3302 1855 5260 1857
rect 3302 1853 3902 1855
rect 3302 1823 3586 1853
rect 2990 1819 3586 1823
rect 3620 1821 3902 1853
rect 3936 1821 4222 1855
rect 4256 1849 5260 1855
rect 4256 1821 4536 1849
rect 3620 1819 4536 1821
rect 2990 1815 4536 1819
rect 4570 1815 4852 1849
rect 4886 1815 5168 1849
rect 5202 1820 5260 1849
rect 2944 1785 5175 1815
rect 2944 1777 3268 1785
rect 2944 1743 2956 1777
rect 2990 1751 3268 1777
rect 3302 1783 5175 1785
rect 3302 1781 3902 1783
rect 3302 1751 3586 1781
rect 2990 1747 3586 1751
rect 3620 1749 3902 1781
rect 3936 1749 4222 1783
rect 4256 1777 5175 1783
rect 4256 1749 4536 1777
rect 3620 1747 4536 1749
rect 2990 1743 4536 1747
rect 4570 1743 4852 1777
rect 4886 1743 5168 1777
rect 5227 1768 5260 1820
rect 5202 1743 5260 1768
rect 2944 1734 5260 1743
rect 5108 1724 5260 1734
rect 2738 -119 2862 62
rect 5594 42 5956 190
rect 5594 -74 5704 42
rect 5820 -74 5956 42
rect 5594 -119 5956 -74
rect 2738 -196 5956 -119
rect 2372 -352 2474 -196
rect 2372 -368 2478 -352
rect -373 -398 2342 -396
rect -631 -412 2342 -398
rect 2372 -402 2405 -368
rect 2439 -402 2478 -368
rect 2372 -406 2478 -402
rect 2378 -410 2478 -406
rect 2874 -370 2976 -196
rect 2874 -404 2907 -370
rect 2941 -404 2976 -370
rect 2874 -410 2976 -404
rect -631 -446 2289 -412
rect 2323 -446 2342 -412
rect -631 -462 2342 -446
rect 3016 -414 5956 -398
rect 3016 -448 3029 -414
rect 3063 -448 5956 -414
rect 2370 -456 2476 -450
rect -631 -641 -269 -462
rect 2370 -490 2405 -456
rect 2439 -490 2476 -456
rect 2366 -558 2476 -490
rect 2872 -458 2982 -452
rect 2872 -492 2907 -458
rect 2941 -492 2982 -458
rect 3016 -464 5956 -448
rect 2872 -558 2982 -492
rect 2362 -568 2982 -558
rect 2362 -602 2412 -568
rect 2446 -572 2982 -568
rect 2446 -602 2908 -572
rect 2362 -606 2908 -602
rect 2942 -606 2982 -572
rect 2362 -620 2982 -606
rect -631 -757 -495 -641
rect -379 -757 -269 -641
rect -631 -905 -269 -757
rect 2622 -728 2708 -620
rect 5594 -641 5956 -464
rect 2622 -982 2706 -728
rect 5594 -757 5704 -641
rect 5820 -757 5956 -641
rect 5594 -905 5956 -757
rect 2622 -1016 2648 -982
rect 2682 -1016 2706 -982
rect 2622 -1018 2706 -1016
rect 1069 -1067 1421 -1019
rect 2626 -1022 2706 -1018
rect 1069 -1101 1372 -1067
rect 1406 -1101 1421 -1067
rect 1069 -1139 1421 -1101
rect 1069 -1173 1372 -1139
rect 1406 -1173 1421 -1139
rect 1069 -1211 1421 -1173
rect 1069 -1222 1372 -1211
rect -694 -1245 1372 -1222
rect 1406 -1245 1421 -1211
rect -694 -1283 1421 -1245
rect -694 -1317 1372 -1283
rect 1406 -1317 1421 -1283
rect -694 -1343 1421 -1317
rect -631 -1465 -269 -1343
rect 1069 -1355 1421 -1343
rect 1069 -1389 1372 -1355
rect 1406 -1389 1421 -1355
rect 1069 -1411 1421 -1389
rect 1069 -1434 1412 -1411
rect -631 -1581 -495 -1465
rect -379 -1581 -269 -1465
rect 1441 -1440 3970 -1432
rect 1441 -1474 1463 -1440
rect 1497 -1474 1535 -1440
rect 1569 -1474 1607 -1440
rect 1641 -1474 1679 -1440
rect 1713 -1474 1751 -1440
rect 1785 -1474 1823 -1440
rect 1857 -1474 1895 -1440
rect 1929 -1474 1967 -1440
rect 2001 -1474 2039 -1440
rect 2073 -1474 2111 -1440
rect 2145 -1474 2183 -1440
rect 2217 -1474 2255 -1440
rect 2289 -1474 2327 -1440
rect 2361 -1474 2399 -1440
rect 2433 -1474 2471 -1440
rect 2505 -1474 2543 -1440
rect 2577 -1474 2615 -1440
rect 2649 -1474 2687 -1440
rect 2721 -1474 2759 -1440
rect 2793 -1474 2831 -1440
rect 2865 -1474 2903 -1440
rect 2937 -1474 2975 -1440
rect 3009 -1474 3047 -1440
rect 3081 -1474 3119 -1440
rect 3153 -1474 3191 -1440
rect 3225 -1474 3263 -1440
rect 3297 -1474 3335 -1440
rect 3369 -1474 3407 -1440
rect 3441 -1474 3479 -1440
rect 3513 -1474 3551 -1440
rect 3585 -1474 3623 -1440
rect 3657 -1474 3695 -1440
rect 3729 -1474 3767 -1440
rect 3801 -1474 3839 -1440
rect 3873 -1474 3911 -1440
rect 3945 -1474 3970 -1440
rect 1441 -1522 3970 -1474
rect -631 -1729 -269 -1581
rect 1170 -1552 4300 -1522
rect 1170 -1586 1487 -1552
rect 1521 -1558 2953 -1552
rect 1521 -1586 1819 -1558
rect 1170 -1592 1819 -1586
rect 1853 -1592 2301 -1558
rect 2335 -1586 2953 -1558
rect 2987 -1554 4300 -1552
rect 2987 -1556 3857 -1554
rect 2987 -1586 3539 -1556
rect 2335 -1590 3539 -1586
rect 3573 -1588 3857 -1556
rect 3891 -1588 4300 -1554
rect 3573 -1590 4300 -1588
rect 2335 -1592 4300 -1590
rect 1170 -1748 4300 -1592
rect 1848 -1939 3912 -1748
rect 1848 -2003 2305 -1939
rect 1848 -3207 2113 -2003
rect 3637 -3143 3912 -1939
rect 3445 -3207 3912 -3143
rect 1848 -3461 3912 -3207
rect 1848 -3510 3751 -3461
<< rmetal1 >>
rect 234 1960 2356 1962
<< via1 >>
rect 1988 3473 3384 4741
rect 93 2544 145 2583
rect 93 2531 115 2544
rect 115 2531 145 2544
rect 93 2510 115 2519
rect 115 2510 145 2519
rect 93 2467 145 2510
rect 5157 2494 5209 2546
rect 93 2052 145 2103
rect 93 2051 100 2052
rect 100 2051 134 2052
rect 134 2051 145 2052
rect 93 2018 100 2039
rect 100 2018 134 2039
rect 134 2018 145 2039
rect 93 1987 145 2018
rect -495 -74 -379 42
rect 5175 1815 5202 1820
rect 5202 1815 5227 1820
rect 5175 1777 5227 1815
rect 5175 1768 5202 1777
rect 5202 1768 5227 1777
rect 5704 -74 5820 42
rect -495 -757 -379 -641
rect 5704 -757 5820 -641
rect -495 -1581 -379 -1465
rect 2305 -2003 3637 -1939
rect 2113 -3143 3637 -2003
rect 2113 -3207 3445 -3143
<< metal2 >>
rect 1739 4774 3642 4973
rect 1739 3438 1945 4774
rect 3441 3438 3642 4774
rect 1739 3195 3642 3438
rect 44 2583 194 2618
rect 44 2531 93 2583
rect 145 2531 194 2583
rect 44 2519 194 2531
rect 44 2467 93 2519
rect 145 2467 194 2519
rect 44 2103 194 2467
rect 44 2051 93 2103
rect 145 2051 194 2103
rect 44 2039 194 2051
rect 44 1987 93 2039
rect 145 1987 194 2039
rect 44 1938 194 1987
rect 5116 2546 5276 2584
rect 5116 2494 5157 2546
rect 5209 2494 5276 2546
rect 5116 1820 5276 2494
rect 5116 1768 5175 1820
rect 5227 1768 5276 1820
rect 5116 1724 5276 1768
rect -631 51 -269 190
rect -631 -85 -503 51
rect -367 -85 -269 51
rect -631 -196 -269 -85
rect 5594 51 5956 190
rect 5594 -85 5692 51
rect 5828 -85 5956 51
rect 5594 -196 5956 -85
rect -631 -631 -269 -519
rect -631 -767 -503 -631
rect -367 -767 -269 -631
rect -631 -905 -269 -767
rect 5594 -631 5956 -519
rect 5594 -767 5692 -631
rect 5828 -767 5956 -631
rect 5594 -905 5956 -767
rect -631 -1455 -269 -1343
rect -631 -1591 -503 -1455
rect -367 -1591 -269 -1455
rect -631 -1729 -269 -1591
rect 2009 -1732 3912 -1683
rect 1848 -1867 3912 -1732
rect 1848 -1947 2215 -1867
rect 1848 -3283 2055 -1947
rect 3711 -3203 3912 -1867
rect 3551 -3283 3912 -3203
rect 1848 -3461 3912 -3283
rect 1848 -3510 3751 -3461
<< via2 >>
rect 1945 4741 3441 4774
rect 1945 3473 1988 4741
rect 1988 3473 3384 4741
rect 3384 3473 3441 4741
rect 1945 3438 3441 3473
rect -503 42 -367 51
rect -503 -74 -495 42
rect -495 -74 -379 42
rect -379 -74 -367 42
rect -503 -85 -367 -74
rect 5692 42 5828 51
rect 5692 -74 5704 42
rect 5704 -74 5820 42
rect 5820 -74 5828 42
rect 5692 -85 5828 -74
rect -503 -641 -367 -631
rect -503 -757 -495 -641
rect -495 -757 -379 -641
rect -379 -757 -367 -641
rect -503 -767 -367 -757
rect 5692 -641 5828 -631
rect 5692 -757 5704 -641
rect 5704 -757 5820 -641
rect 5820 -757 5828 -641
rect 5692 -767 5828 -757
rect -503 -1465 -367 -1455
rect -503 -1581 -495 -1465
rect -495 -1581 -379 -1465
rect -379 -1581 -367 -1465
rect -503 -1591 -367 -1581
rect 2215 -1939 3711 -1867
rect 2215 -1947 2305 -1939
rect 2055 -2003 2305 -1947
rect 2305 -2003 3637 -1939
rect 2055 -3207 2113 -2003
rect 2113 -3143 3637 -2003
rect 3637 -3143 3711 -1939
rect 2113 -3207 3445 -3143
rect 3445 -3203 3711 -3143
rect 3445 -3207 3551 -3203
rect 2055 -3283 3551 -3207
<< metal3 >>
rect 1739 4857 3642 4973
rect 1739 3353 1905 4857
rect 3489 3353 3642 4857
rect 1739 3195 3642 3353
rect -631 97 -269 190
rect -631 -127 -510 97
rect -366 -127 -269 97
rect -631 -196 -269 -127
rect 5594 97 5956 190
rect 5594 -127 5690 97
rect 5834 -127 5956 97
rect 5594 -196 5956 -127
rect -631 -589 -269 -519
rect -631 -813 -510 -589
rect -366 -813 -269 -589
rect -631 -905 -269 -813
rect 5594 -589 5956 -519
rect 5594 -813 5690 -589
rect 5834 -813 5956 -589
rect 5594 -905 5956 -813
rect -631 -1413 -269 -1343
rect -631 -1637 -510 -1413
rect -366 -1637 -269 -1413
rect -631 -1729 -269 -1637
rect 2009 -1732 3912 -1683
rect 1848 -1823 3912 -1732
rect 1848 -1903 2174 -1823
rect 1848 -3327 2014 -1903
rect 3758 -3247 3912 -1823
rect 3598 -3327 3912 -3247
rect 1848 -3461 3912 -3327
rect 1848 -3510 3751 -3461
<< via3 >>
rect 1905 4774 3489 4857
rect 1905 3438 1945 4774
rect 1945 3438 3441 4774
rect 3441 3438 3489 4774
rect 1905 3353 3489 3438
rect -510 51 -366 97
rect -510 -85 -503 51
rect -503 -85 -367 51
rect -367 -85 -366 51
rect -510 -127 -366 -85
rect 5690 51 5834 97
rect 5690 -85 5692 51
rect 5692 -85 5828 51
rect 5828 -85 5834 51
rect 5690 -127 5834 -85
rect -510 -631 -366 -589
rect -510 -767 -503 -631
rect -503 -767 -367 -631
rect -367 -767 -366 -631
rect -510 -813 -366 -767
rect 5690 -631 5834 -589
rect 5690 -767 5692 -631
rect 5692 -767 5828 -631
rect 5828 -767 5834 -631
rect 5690 -813 5834 -767
rect -510 -1455 -366 -1413
rect -510 -1591 -503 -1455
rect -503 -1591 -367 -1455
rect -367 -1591 -366 -1455
rect -510 -1637 -366 -1591
rect 2174 -1867 3758 -1823
rect 2174 -1903 2215 -1867
rect 2014 -1947 2215 -1903
rect 2215 -1947 3711 -1867
rect 2014 -3283 2055 -1947
rect 2055 -3203 3711 -1947
rect 3711 -3203 3758 -1867
rect 2055 -3283 3551 -3203
rect 3551 -3247 3758 -3203
rect 3551 -3283 3598 -3247
rect 2014 -3327 3598 -3283
<< metal4 >>
rect 1739 4857 3642 4973
rect 1739 3353 1905 4857
rect 3489 3353 3642 4857
rect 1739 3338 1934 3353
rect 3450 3338 3642 3353
rect 1739 3195 3642 3338
rect -631 103 -269 190
rect -631 -133 -555 103
rect -319 -133 -269 103
rect -631 -196 -269 -133
rect 5594 103 5956 190
rect 5594 -133 5644 103
rect 5880 -133 5956 103
rect 5594 -196 5956 -133
rect -631 -582 -269 -519
rect -631 -818 -555 -582
rect -319 -818 -269 -582
rect -631 -905 -269 -818
rect 5594 -582 5956 -519
rect 5594 -818 5644 -582
rect 5880 -818 5956 -582
rect 5594 -905 5956 -818
rect -631 -1406 -269 -1343
rect -631 -1642 -555 -1406
rect -319 -1642 -269 -1406
rect -631 -1729 -269 -1642
rect 2009 -1732 3912 -1683
rect 1848 -1823 3912 -1732
rect 1848 -1826 2174 -1823
rect 3758 -1826 3912 -1823
rect 1848 -3342 1964 -1826
rect 3800 -3342 3912 -1826
rect 1848 -3461 3912 -3342
rect 1848 -3510 3751 -3461
<< via4 >>
rect 1934 3353 3450 4854
rect 1934 3338 3450 3353
rect -555 97 -319 103
rect -555 -127 -510 97
rect -510 -127 -366 97
rect -366 -127 -319 97
rect -555 -133 -319 -127
rect 5644 97 5880 103
rect 5644 -127 5690 97
rect 5690 -127 5834 97
rect 5834 -127 5880 97
rect 5644 -133 5880 -127
rect -555 -589 -319 -582
rect -555 -813 -510 -589
rect -510 -813 -366 -589
rect -366 -813 -319 -589
rect -555 -818 -319 -813
rect 5644 -589 5880 -582
rect 5644 -813 5690 -589
rect 5690 -813 5834 -589
rect 5834 -813 5880 -589
rect 5644 -818 5880 -813
rect -555 -1413 -319 -1406
rect -555 -1637 -510 -1413
rect -510 -1637 -366 -1413
rect -366 -1637 -319 -1413
rect -555 -1642 -319 -1637
rect 1964 -1903 2174 -1826
rect 2174 -1903 3758 -1826
rect 1964 -3327 2014 -1903
rect 2014 -3247 3758 -1903
rect 3758 -3247 3800 -1826
rect 2014 -3327 3598 -3247
rect 3598 -3327 3800 -3247
rect 1964 -3342 3800 -3327
<< metal5 >>
rect 1739 4854 3642 4973
rect 1739 3338 1934 4854
rect 3450 3338 3642 4854
rect 1739 3195 3642 3338
rect -694 103 -269 213
rect -694 -133 -555 103
rect -319 -133 -269 103
rect -694 -196 -269 -133
rect 5594 103 6019 213
rect 5594 -133 5644 103
rect 5880 -133 6019 103
rect 5594 -196 6019 -133
rect -694 -582 -269 -519
rect -694 -818 -555 -582
rect -319 -818 -269 -582
rect -694 -928 -269 -818
rect 5594 -582 6019 -519
rect 5594 -818 5644 -582
rect 5880 -818 6019 -582
rect 5594 -928 6019 -818
rect -694 -1406 -269 -1343
rect -694 -1642 -555 -1406
rect -319 -1642 -269 -1406
rect -694 -1752 -269 -1642
rect 2009 -1732 3912 -1683
rect 1848 -1826 3912 -1732
rect 1848 -3342 1964 -1826
rect 3800 -3342 3912 -1826
rect 1848 -3461 3912 -3342
rect 1848 -3510 3751 -3461
use sky130_fd_pr__nfet_01v8_lvt_D42ZUM  sky130_fd_pr__nfet_01v8_lvt_D42ZUM_0
timestamp 1611881054
transform 0 1 2924 -1 0 -431
box -175 -216 175 216
use sky130_fd_pr__nfet_01v8_lvt_D42ZUM  sky130_fd_pr__nfet_01v8_lvt_D42ZUM_1
timestamp 1611881054
transform 0 1 2422 -1 0 -429
box -175 -216 175 216
use sky130_fd_pr__pfet_01v8_NC6LGM  sky130_fd_pr__pfet_01v8_NC6LGM_0
timestamp 1611881054
transform 1 0 1299 0 1 1166
box -1352 -1219 1352 1219
use sky130_fd_pr__pfet_01v8_NC6LGM  sky130_fd_pr__pfet_01v8_NC6LGM_1
timestamp 1611881054
transform 1 0 4000 0 1 1171
box -1352 -1219 1352 1219
use sky130_fd_pr__nfet_01v8_lvt_69NU8X  sky130_fd_pr__nfet_01v8_lvt_69NU8X_0
timestamp 1611881054
transform 0 1 2704 -1 0 -1228
box -360 -1434 360 1434
<< labels >>
rlabel metal1 s 2652 -744 2684 -700 4 Itail_b
rlabel metal1 s 2356 2494 2412 2550 4 Vdd
port 1 nsew
rlabel metal1 s 2460 -134 2516 -78 4 ON2b
port 2 nsew
rlabel metal1 s 2778 -132 2834 -76 4 ON1b
port 3 nsew
rlabel locali s 2314 -438 2330 -418 4 ON1a
port 4 nsew
rlabel locali s 3010 -442 3026 -422 4 ON2a
port 5 nsew
rlabel metal1 s 2664 -1694 2750 -1640 4 Gnd
port 6 nsew
rlabel metal1 s 1370 -1286 1410 -1216 4 vbiasn
port 7 nsew
<< end >>
