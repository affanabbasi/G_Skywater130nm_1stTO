magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect 7862 2528 11846 2532
rect 4870 2486 6072 2490
rect 7862 2486 14424 2528
rect 4870 2238 14424 2486
rect 4870 2218 11846 2238
rect 2628 2202 11846 2218
rect 2628 1796 6072 2202
rect 2628 1726 3080 1796
rect 3086 1787 6072 1796
rect 3086 1752 3101 1787
rect 4577 1752 6072 1787
rect 3086 1726 6072 1752
rect 2628 1725 6072 1726
rect 2628 796 3008 1725
rect 2544 794 3008 796
rect 524 756 3008 794
rect 3042 1040 6072 1725
rect 7862 2140 11846 2202
rect 7862 2092 11450 2140
rect 7862 2058 9501 2092
rect 7862 2040 11450 2058
rect 11494 2040 11846 2140
rect 7862 1702 11846 2040
rect 7862 1650 11506 1702
rect 11552 1650 11846 1702
rect 7862 1646 11846 1650
rect 7862 1635 11478 1646
rect 7862 1634 11453 1635
rect 11469 1634 11478 1635
rect 7862 1600 9501 1634
rect 11477 1600 11478 1634
rect 7862 1576 11478 1600
rect 7862 1568 9486 1576
rect 11436 1572 11478 1576
rect 11436 1568 11474 1572
rect 7862 1474 11474 1568
rect 11492 1474 11846 1646
rect 7862 1442 11846 1474
rect 3042 1010 6000 1040
rect 3042 1008 6070 1010
rect 3042 946 6072 1008
rect 3042 766 4906 946
rect 3042 756 3050 766
rect 524 528 3050 756
rect 4632 738 4678 766
rect 524 400 2766 528
rect 524 198 2566 400
rect 524 -10 1014 198
rect 1588 -6 2566 198
rect 6044 78 7972 568
rect 524 -26 900 -10
<< pwell >>
rect 10518 -856 13588 -842
rect 7216 -858 13588 -856
rect 4424 -860 13588 -858
rect -162 -862 762 -860
rect 2590 -862 13588 -860
rect -162 -942 13588 -862
rect 1798 -944 13588 -942
rect 1798 -946 2622 -944
rect 4424 -946 13588 -944
rect 7216 -948 9712 -946
rect 10518 -954 13588 -946
<< psubdiff >>
rect 10518 -856 13588 -842
rect 7216 -858 13588 -856
rect 4424 -860 13588 -858
rect -162 -862 762 -860
rect 2590 -862 13588 -860
rect -162 -877 13588 -862
rect -162 -879 10707 -877
rect -162 -883 5629 -879
rect -162 -886 2953 -883
rect -162 -920 -53 -886
rect -19 -920 105 -886
rect 139 -920 269 -886
rect 303 -920 421 -886
rect 455 -887 2953 -886
rect 455 -888 782 -887
rect 455 -920 559 -888
rect -162 -922 559 -920
rect 593 -921 782 -888
rect 816 -889 1626 -887
rect 816 -891 1060 -889
rect 816 -921 918 -891
rect 593 -922 918 -921
rect -162 -925 918 -922
rect 952 -923 1060 -891
rect 1094 -891 1340 -889
rect 1094 -923 1204 -891
rect 952 -925 1204 -923
rect 1238 -923 1340 -891
rect 1374 -893 1626 -889
rect 1374 -923 1472 -893
rect 1238 -925 1472 -923
rect -162 -927 1472 -925
rect 1506 -921 1626 -893
rect 1660 -889 2953 -887
rect 1660 -893 1978 -889
rect 1660 -921 1804 -893
rect 1506 -927 1804 -921
rect 1838 -923 1978 -893
rect 2012 -890 2775 -889
rect 2012 -891 2610 -890
rect 2012 -893 2264 -891
rect 2012 -923 2126 -893
rect 1838 -927 2126 -923
rect 2160 -925 2264 -893
rect 2298 -895 2610 -891
rect 2298 -925 2424 -895
rect 2160 -927 2424 -925
rect -162 -929 2424 -927
rect 2458 -924 2610 -895
rect 2644 -923 2775 -890
rect 2809 -917 2953 -889
rect 2987 -887 4323 -883
rect 2987 -917 3125 -887
rect 2809 -921 3125 -917
rect 3159 -921 3309 -887
rect 3343 -889 3827 -887
rect 3343 -921 3465 -889
rect 2809 -923 3465 -921
rect 3499 -923 3641 -889
rect 3675 -921 3827 -889
rect 3861 -921 3983 -887
rect 4017 -921 4155 -887
rect 4189 -917 4323 -887
rect 4357 -917 4455 -883
rect 4489 -887 4849 -883
rect 4489 -889 4719 -887
rect 4489 -917 4585 -889
rect 4189 -921 4585 -917
rect 3675 -923 4585 -921
rect 4619 -921 4719 -889
rect 4753 -917 4849 -887
rect 4883 -887 5135 -883
rect 4883 -917 4997 -887
rect 4753 -921 4997 -917
rect 5031 -917 5135 -887
rect 5169 -887 5461 -883
rect 5169 -917 5297 -887
rect 5031 -921 5297 -917
rect 5331 -917 5461 -887
rect 5495 -913 5629 -883
rect 5663 -883 5921 -879
rect 5663 -913 5773 -883
rect 5495 -917 5773 -913
rect 5807 -913 5921 -883
rect 5955 -883 6509 -879
rect 5955 -913 6077 -883
rect 5807 -917 6077 -913
rect 6111 -917 6223 -883
rect 6257 -917 6369 -883
rect 6403 -913 6509 -883
rect 6543 -887 6907 -879
rect 6543 -913 6653 -887
rect 6403 -917 6653 -913
rect 5331 -921 6653 -917
rect 6687 -921 6787 -887
rect 6821 -913 6907 -887
rect 6941 -883 10707 -879
rect 6941 -913 7039 -883
rect 6821 -917 7039 -913
rect 7073 -917 7171 -883
rect 7205 -885 8229 -883
rect 7205 -917 7313 -885
rect 6821 -919 7313 -917
rect 7347 -889 7791 -885
rect 7347 -919 7461 -889
rect 6821 -921 7461 -919
rect 4619 -923 7461 -921
rect 7495 -893 7791 -889
rect 7495 -923 7623 -893
rect 2644 -924 7623 -923
rect 2458 -927 7623 -924
rect 7657 -919 7791 -893
rect 7825 -919 7939 -885
rect 7973 -919 8081 -885
rect 8115 -917 8229 -885
rect 8263 -885 8651 -883
rect 8263 -917 8381 -885
rect 8115 -919 8381 -917
rect 8415 -919 8511 -885
rect 8545 -917 8651 -885
rect 8685 -885 9699 -883
rect 8685 -917 8839 -885
rect 8545 -919 8839 -917
rect 8873 -919 9019 -885
rect 9053 -919 9187 -885
rect 9221 -889 9543 -885
rect 9221 -919 9381 -889
rect 7657 -923 9381 -919
rect 9415 -919 9543 -889
rect 9577 -917 9699 -885
rect 9733 -917 9857 -883
rect 9891 -885 10707 -883
rect 9891 -917 10041 -885
rect 9577 -919 10041 -917
rect 10075 -919 10225 -885
rect 10259 -919 10389 -885
rect 10423 -887 10707 -885
rect 10423 -919 10545 -887
rect 9415 -921 10545 -919
rect 10579 -911 10707 -887
rect 10741 -911 10901 -877
rect 10935 -881 11301 -877
rect 10935 -911 11091 -881
rect 10579 -915 11091 -911
rect 11125 -911 11301 -881
rect 11335 -881 11867 -877
rect 11335 -911 11495 -881
rect 11125 -915 11495 -911
rect 11529 -887 11867 -881
rect 11529 -915 11681 -887
rect 10579 -921 11681 -915
rect 11715 -911 11867 -887
rect 11901 -881 12631 -877
rect 11901 -887 12221 -881
rect 11901 -911 12047 -887
rect 11715 -921 12047 -911
rect 12081 -915 12221 -887
rect 12255 -915 12431 -881
rect 12465 -911 12631 -881
rect 12665 -911 12831 -877
rect 12865 -911 13065 -877
rect 13099 -881 13588 -877
rect 13099 -911 13323 -881
rect 12465 -915 13323 -911
rect 13357 -915 13588 -881
rect 12081 -921 13588 -915
rect 9415 -923 13588 -921
rect 7657 -927 13588 -923
rect 2458 -929 13588 -927
rect -162 -942 13588 -929
rect 1798 -944 13588 -942
rect 1798 -946 2622 -944
rect 4424 -946 13588 -944
rect 7216 -948 9712 -946
rect 10518 -954 13588 -946
<< nsubdiff >>
rect 11790 2442 14300 2448
rect 11746 2436 14300 2442
rect 8046 2426 14300 2436
rect 5736 2413 14300 2426
rect 5736 2409 9531 2413
rect 5736 2407 8405 2409
rect 5736 2405 6873 2407
rect 5736 2371 5857 2405
rect 5891 2401 6299 2405
rect 5891 2371 6005 2401
rect 5736 2367 6005 2371
rect 6039 2367 6133 2401
rect 6167 2371 6299 2401
rect 6333 2403 6873 2405
rect 6333 2371 6437 2403
rect 6167 2369 6437 2371
rect 6471 2401 6725 2403
rect 6471 2369 6587 2401
rect 6167 2367 6587 2369
rect 6621 2369 6725 2401
rect 6759 2373 6873 2403
rect 6907 2405 8405 2407
rect 6907 2403 7293 2405
rect 6907 2401 7157 2403
rect 6907 2373 7011 2401
rect 6759 2369 7011 2373
rect 6621 2367 7011 2369
rect 7045 2369 7157 2401
rect 7191 2371 7293 2403
rect 7327 2403 7559 2405
rect 7327 2371 7421 2403
rect 7191 2369 7421 2371
rect 7455 2371 7559 2403
rect 7593 2371 7691 2405
rect 7725 2403 8405 2405
rect 7725 2401 7991 2403
rect 7725 2371 7831 2401
rect 7455 2369 7831 2371
rect 7045 2367 7831 2369
rect 7865 2369 7991 2401
rect 8025 2369 8143 2403
rect 8177 2369 8279 2403
rect 8313 2375 8405 2403
rect 8439 2375 8569 2409
rect 8603 2407 8837 2409
rect 8603 2375 8713 2407
rect 8313 2373 8713 2375
rect 8747 2375 8837 2407
rect 8871 2375 9001 2409
rect 9035 2407 9327 2409
rect 9035 2375 9159 2407
rect 8747 2373 9159 2375
rect 9193 2375 9327 2407
rect 9361 2379 9531 2409
rect 9565 2379 9685 2413
rect 9719 2379 9859 2413
rect 9893 2379 10059 2413
rect 10093 2379 10209 2413
rect 10243 2379 10373 2413
rect 10407 2379 10523 2413
rect 10557 2409 10869 2413
rect 10557 2379 10661 2409
rect 9361 2375 10661 2379
rect 10695 2379 10869 2409
rect 10903 2379 11017 2413
rect 11051 2407 11461 2413
rect 11051 2379 11229 2407
rect 10695 2375 11229 2379
rect 9193 2373 11229 2375
rect 11263 2379 11461 2407
rect 11495 2410 14300 2413
rect 11495 2409 11818 2410
rect 11495 2379 11645 2409
rect 11263 2375 11645 2379
rect 11679 2376 11818 2409
rect 11852 2376 11886 2410
rect 11920 2376 11954 2410
rect 11988 2376 12022 2410
rect 12056 2376 12090 2410
rect 12124 2376 12158 2410
rect 12192 2376 12226 2410
rect 12260 2376 12294 2410
rect 12328 2376 12362 2410
rect 12396 2376 12430 2410
rect 12464 2376 12498 2410
rect 12532 2376 12566 2410
rect 12600 2376 12634 2410
rect 12668 2376 12702 2410
rect 12736 2376 12770 2410
rect 12804 2376 12838 2410
rect 12872 2376 12906 2410
rect 12940 2376 12974 2410
rect 13008 2376 13042 2410
rect 13076 2376 13110 2410
rect 13144 2376 13178 2410
rect 13212 2376 13246 2410
rect 13280 2376 13314 2410
rect 13348 2376 13382 2410
rect 13416 2376 13450 2410
rect 13484 2376 13518 2410
rect 13552 2376 13586 2410
rect 13620 2376 13654 2410
rect 13688 2376 13722 2410
rect 13756 2376 13790 2410
rect 13824 2376 13858 2410
rect 13892 2376 13926 2410
rect 13960 2376 13994 2410
rect 14028 2376 14062 2410
rect 14096 2376 14130 2410
rect 14164 2376 14198 2410
rect 14232 2376 14300 2410
rect 11679 2375 14300 2376
rect 11263 2373 14300 2375
rect 8313 2369 14300 2373
rect 7865 2367 14300 2369
rect 5736 2350 14300 2367
rect 5736 2344 8054 2350
rect 11746 2348 14300 2350
rect 11746 2346 11986 2348
rect 2700 2135 4864 2166
rect 2700 2131 4033 2135
rect 2700 2125 3133 2131
rect 2700 2091 2819 2125
rect 2853 2091 2969 2125
rect 3003 2097 3133 2125
rect 3167 2129 4033 2131
rect 3167 2125 3737 2129
rect 3167 2097 3293 2125
rect 3003 2091 3293 2097
rect 3327 2091 3449 2125
rect 3483 2091 3591 2125
rect 3625 2095 3737 2125
rect 3771 2095 3875 2129
rect 3909 2101 4033 2129
rect 4067 2131 4864 2135
rect 4067 2101 4183 2131
rect 3909 2097 4183 2101
rect 4217 2097 4355 2131
rect 4389 2097 4511 2131
rect 4545 2097 4693 2131
rect 4727 2097 4864 2131
rect 3909 2095 4864 2097
rect 3625 2091 4864 2095
rect 2700 2058 4864 2091
rect 700 610 770 612
rect 1694 610 2720 612
rect 700 598 2720 610
rect 700 596 1945 598
rect 700 594 1701 596
rect 700 560 748 594
rect 782 560 864 594
rect 898 560 986 594
rect 1020 560 1106 594
rect 1140 560 1222 594
rect 1256 590 1452 594
rect 1256 560 1326 590
rect 700 556 1326 560
rect 1360 560 1452 590
rect 1486 560 1570 594
rect 1604 562 1701 594
rect 1735 594 1945 596
rect 1735 562 1817 594
rect 1604 560 1817 562
rect 1851 564 1945 594
rect 1979 596 2451 598
rect 1979 594 2189 596
rect 1979 564 2075 594
rect 1851 560 2075 564
rect 2109 562 2189 594
rect 2223 562 2313 596
rect 2347 564 2451 596
rect 2485 564 2577 598
rect 2611 564 2720 598
rect 2347 562 2720 564
rect 2109 560 2720 562
rect 1360 556 2720 560
rect 700 546 2720 556
rect 700 540 770 546
rect 1694 544 2720 546
<< psubdiffcont >>
rect -53 -920 -19 -886
rect 105 -920 139 -886
rect 269 -920 303 -886
rect 421 -920 455 -886
rect 559 -922 593 -888
rect 782 -921 816 -887
rect 918 -925 952 -891
rect 1060 -923 1094 -889
rect 1204 -925 1238 -891
rect 1340 -923 1374 -889
rect 1472 -927 1506 -893
rect 1626 -921 1660 -887
rect 1804 -927 1838 -893
rect 1978 -923 2012 -889
rect 2126 -927 2160 -893
rect 2264 -925 2298 -891
rect 2424 -929 2458 -895
rect 2610 -924 2644 -890
rect 2775 -923 2809 -889
rect 2953 -917 2987 -883
rect 3125 -921 3159 -887
rect 3309 -921 3343 -887
rect 3465 -923 3499 -889
rect 3641 -923 3675 -889
rect 3827 -921 3861 -887
rect 3983 -921 4017 -887
rect 4155 -921 4189 -887
rect 4323 -917 4357 -883
rect 4455 -917 4489 -883
rect 4585 -923 4619 -889
rect 4719 -921 4753 -887
rect 4849 -917 4883 -883
rect 4997 -921 5031 -887
rect 5135 -917 5169 -883
rect 5297 -921 5331 -887
rect 5461 -917 5495 -883
rect 5629 -913 5663 -879
rect 5773 -917 5807 -883
rect 5921 -913 5955 -879
rect 6077 -917 6111 -883
rect 6223 -917 6257 -883
rect 6369 -917 6403 -883
rect 6509 -913 6543 -879
rect 6653 -921 6687 -887
rect 6787 -921 6821 -887
rect 6907 -913 6941 -879
rect 7039 -917 7073 -883
rect 7171 -917 7205 -883
rect 7313 -919 7347 -885
rect 7461 -923 7495 -889
rect 7623 -927 7657 -893
rect 7791 -919 7825 -885
rect 7939 -919 7973 -885
rect 8081 -919 8115 -885
rect 8229 -917 8263 -883
rect 8381 -919 8415 -885
rect 8511 -919 8545 -885
rect 8651 -917 8685 -883
rect 8839 -919 8873 -885
rect 9019 -919 9053 -885
rect 9187 -919 9221 -885
rect 9381 -923 9415 -889
rect 9543 -919 9577 -885
rect 9699 -917 9733 -883
rect 9857 -917 9891 -883
rect 10041 -919 10075 -885
rect 10225 -919 10259 -885
rect 10389 -919 10423 -885
rect 10545 -921 10579 -887
rect 10707 -911 10741 -877
rect 10901 -911 10935 -877
rect 11091 -915 11125 -881
rect 11301 -911 11335 -877
rect 11495 -915 11529 -881
rect 11681 -921 11715 -887
rect 11867 -911 11901 -877
rect 12047 -921 12081 -887
rect 12221 -915 12255 -881
rect 12431 -915 12465 -881
rect 12631 -911 12665 -877
rect 12831 -911 12865 -877
rect 13065 -911 13099 -877
rect 13323 -915 13357 -881
<< nsubdiffcont >>
rect 5857 2371 5891 2405
rect 6005 2367 6039 2401
rect 6133 2367 6167 2401
rect 6299 2371 6333 2405
rect 6437 2369 6471 2403
rect 6587 2367 6621 2401
rect 6725 2369 6759 2403
rect 6873 2373 6907 2407
rect 7011 2367 7045 2401
rect 7157 2369 7191 2403
rect 7293 2371 7327 2405
rect 7421 2369 7455 2403
rect 7559 2371 7593 2405
rect 7691 2371 7725 2405
rect 7831 2367 7865 2401
rect 7991 2369 8025 2403
rect 8143 2369 8177 2403
rect 8279 2369 8313 2403
rect 8405 2375 8439 2409
rect 8569 2375 8603 2409
rect 8713 2373 8747 2407
rect 8837 2375 8871 2409
rect 9001 2375 9035 2409
rect 9159 2373 9193 2407
rect 9327 2375 9361 2409
rect 9531 2379 9565 2413
rect 9685 2379 9719 2413
rect 9859 2379 9893 2413
rect 10059 2379 10093 2413
rect 10209 2379 10243 2413
rect 10373 2379 10407 2413
rect 10523 2379 10557 2413
rect 10661 2375 10695 2409
rect 10869 2379 10903 2413
rect 11017 2379 11051 2413
rect 11229 2373 11263 2407
rect 11461 2379 11495 2413
rect 11645 2375 11679 2409
rect 11818 2376 11852 2410
rect 11886 2376 11920 2410
rect 11954 2376 11988 2410
rect 12022 2376 12056 2410
rect 12090 2376 12124 2410
rect 12158 2376 12192 2410
rect 12226 2376 12260 2410
rect 12294 2376 12328 2410
rect 12362 2376 12396 2410
rect 12430 2376 12464 2410
rect 12498 2376 12532 2410
rect 12566 2376 12600 2410
rect 12634 2376 12668 2410
rect 12702 2376 12736 2410
rect 12770 2376 12804 2410
rect 12838 2376 12872 2410
rect 12906 2376 12940 2410
rect 12974 2376 13008 2410
rect 13042 2376 13076 2410
rect 13110 2376 13144 2410
rect 13178 2376 13212 2410
rect 13246 2376 13280 2410
rect 13314 2376 13348 2410
rect 13382 2376 13416 2410
rect 13450 2376 13484 2410
rect 13518 2376 13552 2410
rect 13586 2376 13620 2410
rect 13654 2376 13688 2410
rect 13722 2376 13756 2410
rect 13790 2376 13824 2410
rect 13858 2376 13892 2410
rect 13926 2376 13960 2410
rect 13994 2376 14028 2410
rect 14062 2376 14096 2410
rect 14130 2376 14164 2410
rect 14198 2376 14232 2410
rect 2819 2091 2853 2125
rect 2969 2091 3003 2125
rect 3133 2097 3167 2131
rect 3293 2091 3327 2125
rect 3449 2091 3483 2125
rect 3591 2091 3625 2125
rect 3737 2095 3771 2129
rect 3875 2095 3909 2129
rect 4033 2101 4067 2135
rect 4183 2097 4217 2131
rect 4355 2097 4389 2131
rect 4511 2097 4545 2131
rect 4693 2097 4727 2131
rect 748 560 782 594
rect 864 560 898 594
rect 986 560 1020 594
rect 1106 560 1140 594
rect 1222 560 1256 594
rect 1326 556 1360 590
rect 1452 560 1486 594
rect 1570 560 1604 594
rect 1701 562 1735 596
rect 1817 560 1851 594
rect 1945 564 1979 598
rect 2075 560 2109 594
rect 2189 562 2223 596
rect 2313 562 2347 596
rect 2451 564 2485 598
rect 2577 564 2611 598
<< locali >>
rect 9412 2421 9464 2426
rect 9412 2420 9421 2421
rect 8320 2416 8372 2418
rect 8846 2416 9421 2420
rect 8022 2414 9421 2416
rect 5764 2413 9421 2414
rect 5764 2409 8329 2413
rect 5764 2407 6659 2409
rect 5764 2405 6219 2407
rect 5764 2401 5857 2405
rect 5764 2367 5797 2401
rect 5831 2371 5857 2401
rect 5891 2371 5927 2405
rect 5961 2401 6071 2405
rect 5961 2371 6005 2401
rect 5831 2367 6005 2371
rect 6039 2371 6071 2401
rect 6105 2401 6219 2405
rect 6105 2371 6133 2401
rect 6039 2367 6133 2371
rect 6167 2373 6219 2401
rect 6253 2405 6363 2407
rect 6253 2373 6299 2405
rect 6167 2371 6299 2373
rect 6333 2373 6363 2405
rect 6397 2405 6659 2407
rect 6397 2403 6503 2405
rect 6397 2373 6437 2403
rect 6333 2371 6437 2373
rect 6167 2369 6437 2371
rect 6471 2371 6503 2403
rect 6537 2401 6659 2405
rect 6537 2371 6587 2401
rect 6471 2369 6587 2371
rect 6167 2367 6587 2369
rect 6621 2375 6659 2401
rect 6693 2407 6947 2409
rect 6693 2405 6873 2407
rect 6693 2403 6799 2405
rect 6693 2375 6725 2403
rect 6621 2369 6725 2375
rect 6759 2371 6799 2403
rect 6833 2373 6873 2405
rect 6907 2375 6947 2407
rect 6981 2407 8065 2409
rect 6981 2405 7357 2407
rect 6981 2401 7085 2405
rect 6981 2375 7011 2401
rect 6907 2373 7011 2375
rect 6833 2371 7011 2373
rect 6759 2369 7011 2371
rect 6621 2367 7011 2369
rect 7045 2371 7085 2401
rect 7119 2403 7215 2405
rect 7119 2371 7157 2403
rect 7045 2369 7157 2371
rect 7191 2371 7215 2403
rect 7249 2371 7293 2405
rect 7327 2373 7357 2405
rect 7391 2403 7485 2407
rect 7391 2373 7421 2403
rect 7327 2371 7421 2373
rect 7191 2369 7421 2371
rect 7455 2373 7485 2403
rect 7519 2405 7913 2407
rect 7519 2373 7559 2405
rect 7455 2371 7559 2373
rect 7593 2371 7623 2405
rect 7657 2371 7691 2405
rect 7725 2403 7913 2405
rect 7725 2371 7755 2403
rect 7455 2369 7755 2371
rect 7789 2401 7913 2403
rect 7789 2369 7831 2401
rect 7045 2367 7831 2369
rect 7865 2373 7913 2401
rect 7947 2403 8065 2407
rect 7947 2373 7991 2403
rect 7865 2369 7991 2373
rect 8025 2375 8065 2403
rect 8099 2407 8329 2409
rect 8099 2403 8215 2407
rect 8099 2375 8143 2403
rect 8025 2369 8143 2375
rect 8177 2373 8215 2403
rect 8249 2403 8329 2407
rect 8249 2373 8279 2403
rect 8177 2369 8279 2373
rect 8313 2379 8329 2403
rect 8363 2409 9225 2413
rect 8363 2379 8405 2409
rect 8313 2375 8405 2379
rect 8439 2375 8479 2409
rect 8513 2375 8569 2409
rect 8603 2375 8623 2409
rect 8657 2407 8763 2409
rect 8657 2375 8713 2407
rect 8313 2373 8713 2375
rect 8747 2375 8763 2407
rect 8797 2375 8837 2409
rect 8871 2375 8907 2409
rect 8941 2375 9001 2409
rect 9035 2375 9065 2409
rect 9099 2407 9225 2409
rect 9099 2375 9159 2407
rect 8747 2373 9159 2375
rect 9193 2379 9225 2407
rect 9259 2409 9421 2413
rect 9259 2379 9327 2409
rect 9193 2375 9327 2379
rect 9361 2387 9421 2409
rect 9455 2420 9464 2421
rect 9600 2423 9652 2428
rect 9600 2420 9609 2423
rect 9455 2413 9609 2420
rect 9455 2387 9531 2413
rect 9361 2379 9531 2387
rect 9565 2389 9609 2413
rect 9643 2420 9652 2423
rect 9764 2420 9816 2422
rect 9942 2420 9994 2422
rect 10110 2421 10162 2426
rect 10110 2420 10119 2421
rect 9643 2417 10119 2420
rect 9643 2413 9773 2417
rect 9643 2389 9685 2413
rect 9565 2379 9685 2389
rect 9719 2383 9773 2413
rect 9807 2413 9951 2417
rect 9807 2383 9859 2413
rect 9719 2379 9859 2383
rect 9893 2383 9951 2413
rect 9985 2413 10119 2417
rect 9985 2383 10059 2413
rect 9893 2379 10059 2383
rect 10093 2387 10119 2413
rect 10153 2420 10162 2421
rect 10278 2421 10330 2426
rect 10278 2420 10287 2421
rect 10153 2413 10287 2420
rect 10153 2387 10209 2413
rect 10093 2379 10209 2387
rect 10243 2387 10287 2413
rect 10321 2420 10330 2421
rect 10442 2423 10494 2428
rect 11124 2427 11176 2432
rect 10442 2420 10451 2423
rect 10321 2413 10451 2420
rect 10321 2387 10373 2413
rect 10243 2379 10373 2387
rect 10407 2389 10451 2413
rect 10485 2420 10494 2423
rect 10578 2421 10630 2426
rect 10578 2420 10587 2421
rect 10485 2413 10587 2420
rect 10485 2389 10523 2413
rect 10407 2379 10523 2389
rect 10557 2387 10587 2413
rect 10621 2420 10630 2421
rect 10760 2421 10812 2426
rect 10760 2420 10769 2421
rect 10621 2409 10769 2420
rect 10621 2387 10661 2409
rect 10557 2379 10661 2387
rect 9361 2375 10661 2379
rect 10695 2387 10769 2409
rect 10803 2420 10812 2421
rect 11124 2420 11133 2427
rect 10803 2413 11133 2420
rect 10803 2387 10869 2413
rect 10695 2379 10869 2387
rect 10903 2407 11017 2413
rect 10903 2379 10921 2407
rect 10695 2375 10921 2379
rect 9193 2373 10921 2375
rect 10955 2379 11017 2407
rect 11051 2393 11133 2413
rect 11167 2420 11176 2427
rect 11348 2431 11400 2436
rect 11348 2420 11357 2431
rect 11167 2407 11357 2420
rect 11167 2393 11229 2407
rect 11051 2379 11229 2393
rect 10955 2373 11229 2379
rect 11263 2397 11357 2407
rect 11391 2420 11400 2431
rect 11538 2431 11590 2436
rect 11538 2420 11547 2431
rect 11391 2413 11547 2420
rect 11391 2397 11461 2413
rect 11263 2379 11461 2397
rect 11495 2397 11547 2413
rect 11581 2420 11590 2431
rect 11716 2420 14266 2422
rect 11581 2417 14266 2420
rect 11581 2409 11725 2417
rect 11581 2397 11645 2409
rect 11495 2379 11645 2397
rect 11263 2375 11645 2379
rect 11679 2383 11725 2409
rect 11759 2410 14266 2417
rect 11759 2383 11818 2410
rect 11679 2376 11818 2383
rect 11854 2376 11886 2410
rect 11926 2376 11954 2410
rect 11998 2376 12022 2410
rect 12070 2376 12090 2410
rect 12142 2376 12158 2410
rect 12214 2376 12226 2410
rect 12286 2376 12294 2410
rect 12358 2376 12362 2410
rect 12464 2376 12468 2410
rect 12532 2376 12540 2410
rect 12600 2376 12612 2410
rect 12668 2376 12684 2410
rect 12736 2376 12756 2410
rect 12804 2376 12828 2410
rect 12872 2376 12900 2410
rect 12940 2376 12972 2410
rect 13008 2376 13042 2410
rect 13078 2376 13110 2410
rect 13150 2376 13178 2410
rect 13222 2376 13246 2410
rect 13294 2376 13314 2410
rect 13366 2376 13382 2410
rect 13438 2376 13450 2410
rect 13510 2376 13518 2410
rect 13582 2376 13586 2410
rect 13688 2376 13692 2410
rect 13756 2376 13764 2410
rect 13824 2376 13836 2410
rect 13892 2376 13908 2410
rect 13960 2376 13980 2410
rect 14028 2376 14052 2410
rect 14096 2376 14124 2410
rect 14164 2376 14196 2410
rect 14232 2376 14266 2410
rect 11679 2375 14266 2376
rect 11263 2373 14266 2375
rect 8313 2369 14266 2373
rect 7865 2368 14266 2369
rect 7865 2367 11304 2368
rect 5764 2364 11304 2367
rect 5764 2362 8032 2364
rect 6122 2150 6150 2184
rect 6184 2150 6222 2184
rect 6256 2150 6294 2184
rect 6328 2150 6366 2184
rect 6400 2150 6438 2184
rect 6472 2150 6510 2184
rect 6544 2150 6582 2184
rect 6616 2150 6654 2184
rect 6688 2150 6726 2184
rect 6760 2150 6798 2184
rect 6832 2150 6870 2184
rect 6904 2150 6942 2184
rect 6976 2150 7014 2184
rect 7048 2150 7086 2184
rect 7120 2150 7158 2184
rect 7192 2150 7230 2184
rect 7264 2150 7302 2184
rect 7336 2150 7374 2184
rect 7408 2150 7446 2184
rect 7480 2150 7518 2184
rect 7552 2150 7590 2184
rect 7624 2150 7662 2184
rect 7696 2150 7734 2184
rect 7768 2150 7796 2184
rect 9402 2172 9428 2206
rect 9462 2172 9500 2206
rect 9534 2172 9572 2206
rect 9606 2172 9644 2206
rect 9678 2172 9716 2206
rect 9750 2172 9788 2206
rect 9822 2172 9860 2206
rect 9894 2172 9932 2206
rect 9966 2172 10004 2206
rect 10038 2172 10076 2206
rect 10110 2172 10148 2206
rect 10182 2172 10220 2206
rect 10254 2172 10292 2206
rect 10326 2172 10364 2206
rect 10398 2172 10436 2206
rect 10470 2172 10508 2206
rect 10542 2172 10580 2206
rect 10614 2172 10652 2206
rect 10686 2172 10724 2206
rect 10758 2172 10796 2206
rect 10830 2172 10868 2206
rect 10902 2172 10940 2206
rect 10974 2172 11012 2206
rect 11046 2172 11084 2206
rect 11118 2172 11156 2206
rect 11190 2172 11228 2206
rect 11262 2172 11300 2206
rect 11334 2172 11372 2206
rect 11406 2172 11444 2206
rect 11478 2172 11516 2206
rect 11550 2172 11576 2206
rect 11976 2170 12002 2204
rect 12036 2170 12074 2204
rect 12108 2170 12146 2204
rect 12180 2170 12218 2204
rect 12252 2170 12290 2204
rect 12324 2170 12362 2204
rect 12396 2170 12434 2204
rect 12468 2170 12506 2204
rect 12540 2170 12578 2204
rect 12612 2170 12650 2204
rect 12684 2170 12722 2204
rect 12756 2170 12794 2204
rect 12828 2170 12866 2204
rect 12900 2170 12938 2204
rect 12972 2170 13010 2204
rect 13044 2170 13082 2204
rect 13116 2170 13154 2204
rect 13188 2170 13226 2204
rect 13260 2170 13298 2204
rect 13332 2170 13370 2204
rect 13404 2170 13442 2204
rect 13476 2170 13514 2204
rect 13548 2170 13586 2204
rect 13620 2170 13658 2204
rect 13692 2170 13730 2204
rect 13764 2170 13802 2204
rect 13836 2170 13874 2204
rect 13908 2170 13946 2204
rect 13980 2170 14018 2204
rect 14052 2170 14090 2204
rect 14124 2170 14150 2204
rect 2722 2135 4842 2150
rect 2722 2131 4033 2135
rect 2722 2129 2885 2131
rect 2722 2095 2751 2129
rect 2785 2125 2885 2129
rect 2785 2095 2819 2125
rect 2722 2091 2819 2095
rect 2853 2097 2885 2125
rect 2919 2129 3133 2131
rect 2919 2125 3045 2129
rect 2919 2097 2969 2125
rect 2853 2091 2969 2097
rect 3003 2095 3045 2125
rect 3079 2097 3133 2129
rect 3167 2097 3219 2131
rect 3253 2129 3519 2131
rect 3253 2125 3367 2129
rect 3253 2097 3293 2125
rect 3079 2095 3293 2097
rect 3003 2091 3293 2095
rect 3327 2095 3367 2125
rect 3401 2125 3519 2129
rect 3401 2095 3449 2125
rect 3327 2091 3449 2095
rect 3483 2097 3519 2125
rect 3553 2129 3791 2131
rect 3553 2125 3655 2129
rect 3553 2097 3591 2125
rect 3483 2091 3591 2097
rect 3625 2095 3655 2125
rect 3689 2095 3737 2129
rect 3771 2097 3791 2129
rect 3825 2129 4033 2131
rect 3825 2097 3875 2129
rect 3771 2095 3875 2097
rect 3909 2095 3943 2129
rect 3977 2101 4033 2129
rect 4067 2131 4269 2135
rect 4067 2101 4101 2131
rect 3977 2097 4101 2101
rect 4135 2097 4183 2131
rect 4217 2101 4269 2131
rect 4303 2131 4842 2135
rect 4303 2101 4355 2131
rect 4217 2097 4355 2101
rect 4389 2097 4427 2131
rect 4461 2097 4511 2131
rect 4545 2129 4693 2131
rect 4545 2097 4603 2129
rect 3977 2095 4603 2097
rect 4637 2097 4693 2129
rect 4727 2097 4765 2131
rect 4799 2097 4842 2131
rect 4637 2095 4842 2097
rect 3625 2091 4842 2095
rect 2722 2078 4842 2091
rect 3002 1866 3030 1900
rect 3064 1866 3102 1900
rect 3136 1866 3174 1900
rect 3208 1866 3246 1900
rect 3280 1866 3318 1900
rect 3352 1866 3390 1900
rect 3424 1866 3462 1900
rect 3496 1866 3534 1900
rect 3568 1866 3606 1900
rect 3640 1866 3678 1900
rect 3712 1866 3750 1900
rect 3784 1866 3822 1900
rect 3856 1866 3894 1900
rect 3928 1866 3966 1900
rect 4000 1866 4038 1900
rect 4072 1866 4110 1900
rect 4144 1866 4182 1900
rect 4216 1866 4254 1900
rect 4288 1866 4326 1900
rect 4360 1866 4398 1900
rect 4432 1866 4470 1900
rect 4504 1866 4542 1900
rect 4576 1866 4614 1900
rect 4648 1866 4676 1900
rect 2244 600 2292 602
rect 704 598 2251 600
rect 704 596 1274 598
rect 704 594 800 596
rect 704 560 748 594
rect 782 562 800 594
rect 834 594 1042 596
rect 834 562 864 594
rect 782 560 864 562
rect 898 592 986 594
rect 898 560 922 592
rect 704 558 922 560
rect 956 560 986 592
rect 1020 562 1042 594
rect 1076 594 1274 596
rect 1076 562 1106 594
rect 1020 560 1106 562
rect 1140 592 1222 594
rect 1140 560 1164 592
rect 956 558 1164 560
rect 1198 560 1222 592
rect 1256 564 1274 594
rect 1308 596 1945 598
rect 1308 594 1701 596
rect 1308 590 1384 594
rect 1308 564 1326 590
rect 1256 560 1326 564
rect 1198 558 1326 560
rect 704 556 1326 558
rect 1360 560 1384 590
rect 1418 560 1452 594
rect 1486 560 1506 594
rect 1540 560 1570 594
rect 1604 560 1638 594
rect 1672 562 1701 594
rect 1735 562 1757 596
rect 1791 594 1881 596
rect 1791 562 1817 594
rect 1672 560 1817 562
rect 1851 562 1881 594
rect 1915 564 1945 596
rect 1979 596 2123 598
rect 1979 564 2007 596
rect 1915 562 2007 564
rect 2041 594 2123 596
rect 2041 562 2075 594
rect 1851 560 2075 562
rect 2109 564 2123 594
rect 2157 596 2251 598
rect 2157 564 2189 596
rect 2109 562 2189 564
rect 2223 566 2251 596
rect 2285 598 2710 600
rect 2285 596 2451 598
rect 2285 566 2313 596
rect 2223 562 2313 566
rect 2347 594 2451 596
rect 2347 562 2383 594
rect 2109 560 2383 562
rect 2417 564 2451 594
rect 2485 564 2521 598
rect 2555 564 2577 598
rect 2611 594 2710 598
rect 2611 564 2623 594
rect 2417 560 2623 564
rect 2657 560 2710 594
rect 1360 558 2710 560
rect 1360 556 1702 558
rect 704 554 1702 556
rect 704 552 766 554
rect 5568 484 5594 518
rect 5628 484 5666 518
rect 5700 484 5738 518
rect 5772 484 5810 518
rect 5844 484 5882 518
rect 5916 484 5942 518
rect 8020 498 8046 532
rect 8080 498 8118 532
rect 8152 498 8190 532
rect 8224 498 8262 532
rect 8296 498 8334 532
rect 8368 498 8394 532
rect 1132 344 1158 378
rect 1192 344 1230 378
rect 1264 344 1302 378
rect 1336 344 1374 378
rect 1408 344 1446 378
rect 1480 344 1506 378
rect 5667 370 5702 404
rect 5736 370 5774 404
rect 5808 370 5843 404
rect 8119 384 8154 418
rect 8188 384 8226 418
rect 8260 384 8295 418
rect 11084 410 11101 444
rect 11135 410 11173 444
rect 11207 410 11245 444
rect 11279 410 11317 444
rect 11351 410 11389 444
rect 11423 410 11461 444
rect 11495 410 11533 444
rect 11567 410 11605 444
rect 11639 410 11677 444
rect 11711 410 11749 444
rect 11783 410 11821 444
rect 11855 410 11893 444
rect 11927 410 11965 444
rect 11999 410 12037 444
rect 12071 410 12109 444
rect 12143 410 12181 444
rect 12215 410 12253 444
rect 12287 410 12325 444
rect 12359 410 12397 444
rect 12431 410 12469 444
rect 12503 410 12541 444
rect 12575 410 12613 444
rect 12647 410 12685 444
rect 12719 410 12757 444
rect 12791 410 12829 444
rect 12863 410 12901 444
rect 12935 410 12973 444
rect 13007 410 13045 444
rect 13079 410 13117 444
rect 13151 410 13189 444
rect 13223 410 13240 444
rect 2102 336 2128 370
rect 2162 336 2200 370
rect 2234 336 2272 370
rect 2306 336 2344 370
rect 2378 336 2416 370
rect 2450 336 2476 370
rect 8354 354 8388 356
rect 5902 340 5936 342
rect 8354 318 8388 320
rect 5902 304 5936 306
rect 1231 230 1266 264
rect 1300 230 1338 264
rect 1372 230 1407 264
rect 2201 222 2236 256
rect 2270 222 2308 256
rect 2342 222 2377 256
rect 3498 216 3511 250
rect 3545 216 3558 250
rect 5667 242 5702 276
rect 5736 242 5774 276
rect 5808 242 5843 276
rect 8119 256 8154 290
rect 8188 256 8226 290
rect 8260 256 8295 290
rect 1231 142 1266 176
rect 1300 142 1338 176
rect 1372 142 1407 176
rect 2201 134 2236 168
rect 2270 134 2308 168
rect 2342 134 2377 168
rect 3498 128 3511 162
rect 3545 128 3558 162
rect 3408 14 3439 48
rect 3473 14 3511 48
rect 3545 14 3583 48
rect 3617 14 3648 48
rect 11030 -142 11049 -108
rect 11083 -142 11121 -108
rect 11155 -142 11193 -108
rect 11227 -142 11265 -108
rect 11299 -142 11337 -108
rect 11371 -142 11409 -108
rect 11443 -142 11481 -108
rect 11515 -142 11553 -108
rect 11587 -142 11625 -108
rect 11659 -142 11697 -108
rect 11731 -142 11769 -108
rect 11803 -142 11841 -108
rect 11875 -142 11913 -108
rect 11947 -142 11985 -108
rect 12019 -142 12057 -108
rect 12091 -142 12129 -108
rect 12163 -142 12201 -108
rect 12235 -142 12273 -108
rect 12307 -142 12345 -108
rect 12379 -142 12417 -108
rect 12451 -142 12489 -108
rect 12523 -142 12561 -108
rect 12595 -142 12633 -108
rect 12667 -142 12705 -108
rect 12739 -142 12777 -108
rect 12811 -142 12849 -108
rect 12883 -142 12921 -108
rect 12955 -142 12993 -108
rect 13027 -142 13065 -108
rect 13099 -142 13137 -108
rect 13171 -142 13209 -108
rect 13243 -142 13281 -108
rect 13315 -142 13353 -108
rect 13387 -142 13406 -108
rect 10946 -193 10980 -170
rect 10946 -265 10980 -227
rect 10946 -337 10980 -299
rect 10946 -409 10980 -371
rect 306 -482 319 -448
rect 353 -482 366 -448
rect 2296 -470 2334 -436
rect 3932 -456 3945 -422
rect 3979 -456 3992 -422
rect 4710 -448 4713 -414
rect 4747 -448 4785 -414
rect 4819 -448 4857 -414
rect 4891 -448 4929 -414
rect 4963 -448 5001 -414
rect 5035 -448 5073 -414
rect 5107 -448 5145 -414
rect 5179 -448 5217 -414
rect 5251 -448 5289 -414
rect 5323 -448 5361 -414
rect 5395 -448 5433 -414
rect 5467 -448 5505 -414
rect 5539 -448 5577 -414
rect 5611 -448 5649 -414
rect 5683 -448 5686 -414
rect 5928 -448 5931 -414
rect 5965 -448 6003 -414
rect 6037 -448 6075 -414
rect 6109 -448 6147 -414
rect 6181 -448 6219 -414
rect 6253 -448 6291 -414
rect 6325 -448 6363 -414
rect 6397 -448 6435 -414
rect 6469 -448 6507 -414
rect 6541 -448 6579 -414
rect 6613 -448 6651 -414
rect 6685 -448 6723 -414
rect 6757 -448 6795 -414
rect 6829 -448 6867 -414
rect 6901 -448 6904 -414
rect 7828 -446 7831 -412
rect 7865 -446 7903 -412
rect 7937 -446 7975 -412
rect 8009 -446 8047 -412
rect 8081 -446 8119 -412
rect 8153 -446 8191 -412
rect 8225 -446 8263 -412
rect 8297 -446 8335 -412
rect 8369 -446 8407 -412
rect 8441 -446 8479 -412
rect 8513 -446 8551 -412
rect 8585 -446 8623 -412
rect 8657 -446 8695 -412
rect 8729 -446 8767 -412
rect 8801 -446 8804 -412
rect 9046 -446 9049 -412
rect 9083 -446 9121 -412
rect 9155 -446 9193 -412
rect 9227 -446 9265 -412
rect 9299 -446 9337 -412
rect 9371 -446 9409 -412
rect 9443 -446 9481 -412
rect 9515 -446 9553 -412
rect 9587 -446 9625 -412
rect 9659 -446 9697 -412
rect 9731 -446 9769 -412
rect 9803 -446 9841 -412
rect 9875 -446 9913 -412
rect 9947 -446 9985 -412
rect 10019 -446 10022 -412
rect 3078 -508 3082 -474
rect 5748 -476 5790 -460
rect 5742 -493 5790 -476
rect 306 -570 319 -536
rect 353 -570 366 -536
rect 2296 -558 2334 -524
rect 3932 -544 3945 -510
rect 3979 -544 3992 -510
rect 5776 -527 5790 -493
rect 5742 -544 5790 -527
rect 5748 -560 5790 -544
rect 5830 -493 5872 -462
rect 5830 -527 5838 -493
rect 5830 -562 5872 -527
rect 6954 -493 6988 -476
rect 6954 -544 6988 -527
rect 7744 -491 7778 -474
rect 7744 -542 7778 -525
rect 8854 -491 8888 -474
rect 8854 -542 8888 -525
rect 8962 -491 8996 -474
rect 8962 -542 8996 -525
rect 10946 -481 10980 -443
rect 10946 -538 10980 -515
rect 4710 -606 4713 -572
rect 4747 -606 4785 -572
rect 4819 -606 4857 -572
rect 4891 -606 4929 -572
rect 4963 -606 5001 -572
rect 5035 -606 5073 -572
rect 5107 -606 5145 -572
rect 5179 -606 5217 -572
rect 5251 -606 5289 -572
rect 5323 -606 5361 -572
rect 5395 -606 5433 -572
rect 5467 -606 5505 -572
rect 5539 -606 5577 -572
rect 5611 -606 5649 -572
rect 5683 -606 5686 -572
rect 5928 -606 5931 -572
rect 5965 -606 6003 -572
rect 6037 -606 6075 -572
rect 6109 -606 6147 -572
rect 6181 -606 6219 -572
rect 6253 -606 6291 -572
rect 6325 -606 6363 -572
rect 6397 -606 6435 -572
rect 6469 -606 6507 -572
rect 6541 -606 6579 -572
rect 6613 -606 6651 -572
rect 6685 -606 6723 -572
rect 6757 -606 6795 -572
rect 6829 -606 6867 -572
rect 6901 -606 6904 -572
rect 7828 -604 7831 -570
rect 7865 -604 7903 -570
rect 7937 -604 7975 -570
rect 8009 -604 8047 -570
rect 8081 -604 8119 -570
rect 8153 -604 8191 -570
rect 8225 -604 8263 -570
rect 8297 -604 8335 -570
rect 8369 -604 8407 -570
rect 8441 -604 8479 -570
rect 8513 -604 8551 -570
rect 8585 -604 8623 -570
rect 8657 -604 8695 -570
rect 8729 -604 8767 -570
rect 8801 -604 8804 -570
rect 9046 -604 9049 -570
rect 9083 -604 9121 -570
rect 9155 -604 9193 -570
rect 9227 -604 9265 -570
rect 9299 -604 9337 -570
rect 9371 -604 9409 -570
rect 9443 -604 9481 -570
rect 9515 -604 9553 -570
rect 9587 -604 9625 -570
rect 9659 -604 9697 -570
rect 9731 -604 9769 -570
rect 9803 -604 9841 -570
rect 9875 -604 9913 -570
rect 9947 -604 9985 -570
rect 10019 -604 10022 -570
rect 11030 -600 11049 -566
rect 11083 -600 11121 -566
rect 11155 -600 11193 -566
rect 11227 -600 11265 -566
rect 11299 -600 11337 -566
rect 11371 -600 11409 -566
rect 11443 -600 11481 -566
rect 11515 -600 11553 -566
rect 11587 -600 11625 -566
rect 11659 -600 11697 -566
rect 11731 -600 11769 -566
rect 11803 -600 11841 -566
rect 11875 -600 11913 -566
rect 11947 -600 11985 -566
rect 12019 -600 12057 -566
rect 12091 -600 12129 -566
rect 12163 -600 12201 -566
rect 12235 -600 12273 -566
rect 12307 -600 12345 -566
rect 12379 -600 12417 -566
rect 12451 -600 12489 -566
rect 12523 -600 12561 -566
rect 12595 -600 12633 -566
rect 12667 -600 12705 -566
rect 12739 -600 12777 -566
rect 12811 -600 12849 -566
rect 12883 -600 12921 -566
rect 12955 -600 12993 -566
rect 13027 -600 13065 -566
rect 13099 -600 13137 -566
rect 13171 -600 13209 -566
rect 13243 -600 13281 -566
rect 13315 -600 13353 -566
rect 13387 -600 13406 -566
rect 216 -684 247 -650
rect 281 -684 319 -650
rect 353 -684 391 -650
rect 425 -684 456 -650
rect 1192 -676 1210 -642
rect 1244 -676 1282 -642
rect 1316 -676 1354 -642
rect 1388 -676 1426 -642
rect 1460 -676 1478 -642
rect 2172 -672 2190 -638
rect 2224 -672 2262 -638
rect 2296 -672 2334 -638
rect 2368 -672 2406 -638
rect 2440 -672 2458 -638
rect 3052 -666 3083 -632
rect 3117 -666 3155 -632
rect 3189 -666 3227 -632
rect 3261 -666 3292 -632
rect 3842 -658 3873 -624
rect 3907 -658 3945 -624
rect 3979 -658 4017 -624
rect 4051 -658 4082 -624
rect 4620 -720 4638 -686
rect 4672 -720 4710 -686
rect 4744 -720 4782 -686
rect 4816 -720 4854 -686
rect 4888 -720 4926 -686
rect 4960 -720 4998 -686
rect 5032 -720 5070 -686
rect 5104 -720 5142 -686
rect 5176 -720 5214 -686
rect 5248 -720 5286 -686
rect 5320 -720 5358 -686
rect 5392 -720 5430 -686
rect 5464 -720 5502 -686
rect 5536 -720 5574 -686
rect 5608 -720 5646 -686
rect 5680 -720 5718 -686
rect 5752 -720 5790 -686
rect 5824 -720 5862 -686
rect 5896 -720 5934 -686
rect 5968 -720 6006 -686
rect 6040 -720 6078 -686
rect 6112 -720 6150 -686
rect 6184 -720 6222 -686
rect 6256 -720 6294 -686
rect 6328 -720 6366 -686
rect 6400 -720 6438 -686
rect 6472 -720 6510 -686
rect 6544 -720 6582 -686
rect 6616 -720 6654 -686
rect 6688 -720 6726 -686
rect 6760 -720 6798 -686
rect 6832 -720 6870 -686
rect 6904 -720 6942 -686
rect 6976 -720 6994 -686
rect 7738 -718 7756 -684
rect 7790 -718 7828 -684
rect 7862 -718 7900 -684
rect 7934 -718 7972 -684
rect 8006 -718 8044 -684
rect 8078 -718 8116 -684
rect 8150 -718 8188 -684
rect 8222 -718 8260 -684
rect 8294 -718 8332 -684
rect 8366 -718 8404 -684
rect 8438 -718 8476 -684
rect 8510 -718 8548 -684
rect 8582 -718 8620 -684
rect 8654 -718 8692 -684
rect 8726 -718 8764 -684
rect 8798 -718 8836 -684
rect 8870 -718 8908 -684
rect 8942 -718 8980 -684
rect 9014 -718 9052 -684
rect 9086 -718 9124 -684
rect 9158 -718 9196 -684
rect 9230 -718 9268 -684
rect 9302 -718 9340 -684
rect 9374 -718 9412 -684
rect 9446 -718 9484 -684
rect 9518 -718 9556 -684
rect 9590 -718 9628 -684
rect 9662 -718 9700 -684
rect 9734 -718 9772 -684
rect 9806 -718 9844 -684
rect 9878 -718 9916 -684
rect 9950 -718 9988 -684
rect 10022 -718 10060 -684
rect 10094 -718 10112 -684
rect 10940 -714 10941 -680
rect 10975 -714 11013 -680
rect 11047 -714 11085 -680
rect 11119 -714 11157 -680
rect 11191 -714 11229 -680
rect 11263 -714 11301 -680
rect 11335 -714 11373 -680
rect 11407 -714 11445 -680
rect 11479 -714 11517 -680
rect 11551 -714 11589 -680
rect 11623 -714 11661 -680
rect 11695 -714 11733 -680
rect 11767 -714 11805 -680
rect 11839 -714 11877 -680
rect 11911 -714 11949 -680
rect 11983 -714 12021 -680
rect 12055 -714 12093 -680
rect 12127 -714 12165 -680
rect 12199 -714 12237 -680
rect 12271 -714 12309 -680
rect 12343 -714 12381 -680
rect 12415 -714 12453 -680
rect 12487 -714 12525 -680
rect 12559 -714 12597 -680
rect 12631 -714 12669 -680
rect 12703 -714 12741 -680
rect 12775 -714 12813 -680
rect 12847 -714 12885 -680
rect 12919 -714 12957 -680
rect 12991 -714 13029 -680
rect 13063 -714 13101 -680
rect 13135 -714 13173 -680
rect 13207 -714 13245 -680
rect 13279 -714 13317 -680
rect 13351 -714 13389 -680
rect 13423 -714 13461 -680
rect 13495 -714 13496 -680
rect 11586 -862 11646 -856
rect 4638 -872 4690 -870
rect 4776 -872 4828 -870
rect 4912 -872 4964 -870
rect 5054 -872 5106 -870
rect 5542 -872 5594 -870
rect 5992 -872 6044 -870
rect 7650 -872 9262 -870
rect 10470 -871 13554 -862
rect 10470 -872 11599 -871
rect 4402 -874 9262 -872
rect 10454 -874 11599 -872
rect 2690 -876 2748 -874
rect 2858 -876 2916 -874
rect 3030 -876 3088 -874
rect 3208 -876 3266 -874
rect 4060 -876 4118 -874
rect 4240 -876 4298 -874
rect 4402 -876 11599 -874
rect 2584 -877 11599 -876
rect 2584 -878 4647 -877
rect 742 -880 4647 -878
rect -144 -883 4647 -880
rect -144 -884 2953 -883
rect -144 -886 2702 -884
rect -144 -888 -53 -886
rect -144 -922 -123 -888
rect -89 -920 -53 -888
rect -19 -888 105 -886
rect -19 -920 27 -888
rect -89 -922 27 -920
rect 61 -920 105 -888
rect 139 -920 185 -886
rect 219 -920 269 -886
rect 303 -888 421 -886
rect 303 -920 333 -888
rect 61 -922 333 -920
rect 367 -920 421 -888
rect 455 -887 2702 -886
rect 455 -888 716 -887
rect 455 -920 483 -888
rect 367 -922 483 -920
rect 517 -922 559 -888
rect 593 -922 629 -888
rect 663 -921 716 -888
rect 750 -921 782 -887
rect 816 -891 984 -887
rect 816 -921 846 -891
rect 663 -922 846 -921
rect -144 -925 846 -922
rect 880 -925 918 -891
rect 952 -921 984 -891
rect 1018 -889 1556 -887
rect 1018 -921 1060 -889
rect 952 -923 1060 -921
rect 1094 -923 1126 -889
rect 1160 -891 1340 -889
rect 1160 -923 1204 -891
rect 952 -925 1204 -923
rect 1238 -893 1340 -891
rect 1238 -925 1268 -893
rect -144 -927 1268 -925
rect 1302 -923 1340 -893
rect 1374 -923 1414 -889
rect 1448 -893 1556 -889
rect 1448 -923 1472 -893
rect 1302 -927 1472 -923
rect 1506 -921 1556 -893
rect 1590 -921 1626 -887
rect 1660 -921 1728 -887
rect 1762 -889 2702 -887
rect 1762 -891 1978 -889
rect 1762 -893 1896 -891
rect 1762 -921 1804 -893
rect 1506 -927 1804 -921
rect 1838 -925 1896 -893
rect 1930 -923 1978 -891
rect 2012 -923 2050 -889
rect 2084 -893 2198 -889
rect 2084 -923 2126 -893
rect 1930 -925 2126 -923
rect 1838 -927 2126 -925
rect 2160 -923 2198 -893
rect 2232 -891 2340 -889
rect 2232 -923 2264 -891
rect 2160 -925 2264 -923
rect 2298 -923 2340 -891
rect 2374 -895 2510 -889
rect 2374 -923 2424 -895
rect 2298 -925 2424 -923
rect 2160 -927 2424 -925
rect -144 -929 2424 -927
rect 2458 -923 2510 -895
rect 2544 -890 2702 -889
rect 2544 -923 2610 -890
rect 2458 -924 2610 -923
rect 2644 -918 2702 -890
rect 2736 -889 2870 -884
rect 2736 -918 2775 -889
rect 2644 -923 2775 -918
rect 2809 -918 2870 -889
rect 2904 -917 2953 -884
rect 2987 -884 4323 -883
rect 2987 -917 3042 -884
rect 2904 -918 3042 -917
rect 3076 -887 3220 -884
rect 3076 -918 3125 -887
rect 2809 -921 3125 -918
rect 3159 -918 3220 -887
rect 3254 -886 4072 -884
rect 3254 -887 3392 -886
rect 3254 -918 3309 -887
rect 3159 -921 3309 -918
rect 3343 -920 3392 -887
rect 3426 -889 3742 -886
rect 3426 -920 3465 -889
rect 3343 -921 3465 -920
rect 2809 -923 3465 -921
rect 3499 -890 3641 -889
rect 3499 -923 3558 -890
rect 2644 -924 3558 -923
rect 3592 -923 3641 -890
rect 3675 -920 3742 -889
rect 3776 -887 3912 -886
rect 3776 -920 3827 -887
rect 3675 -921 3827 -920
rect 3861 -920 3912 -887
rect 3946 -887 4072 -886
rect 3946 -920 3983 -887
rect 3861 -921 3983 -920
rect 4017 -918 4072 -887
rect 4106 -887 4252 -884
rect 4106 -918 4155 -887
rect 4017 -921 4155 -918
rect 4189 -918 4252 -887
rect 4286 -917 4323 -884
rect 4357 -917 4393 -883
rect 4427 -917 4455 -883
rect 4489 -917 4517 -883
rect 4551 -889 4647 -883
rect 4551 -917 4585 -889
rect 4286 -918 4585 -917
rect 4189 -921 4585 -918
rect 3675 -923 4585 -921
rect 4619 -911 4647 -889
rect 4681 -887 4785 -877
rect 4681 -911 4719 -887
rect 4619 -921 4719 -911
rect 4753 -911 4785 -887
rect 4819 -883 4921 -877
rect 4819 -911 4849 -883
rect 4753 -917 4849 -911
rect 4883 -911 4921 -883
rect 4955 -887 5063 -877
rect 4955 -911 4997 -887
rect 4883 -917 4997 -911
rect 4753 -921 4997 -917
rect 5031 -911 5063 -887
rect 5097 -883 5551 -877
rect 5097 -911 5135 -883
rect 5031 -917 5135 -911
rect 5169 -917 5221 -883
rect 5255 -887 5389 -883
rect 5255 -917 5297 -887
rect 5031 -921 5297 -917
rect 5331 -917 5389 -887
rect 5423 -917 5461 -883
rect 5495 -911 5551 -883
rect 5585 -879 6001 -877
rect 5585 -911 5629 -879
rect 5495 -913 5629 -911
rect 5663 -883 5845 -879
rect 5663 -913 5691 -883
rect 5495 -917 5691 -913
rect 5725 -917 5773 -883
rect 5807 -913 5845 -883
rect 5879 -913 5921 -879
rect 5955 -911 6001 -879
rect 6035 -879 10707 -877
rect 6035 -883 6293 -879
rect 6035 -911 6077 -883
rect 5955 -913 6077 -911
rect 5807 -917 6077 -913
rect 6111 -917 6151 -883
rect 6185 -917 6223 -883
rect 6257 -913 6293 -883
rect 6327 -883 6441 -879
rect 6327 -913 6369 -883
rect 6257 -917 6369 -913
rect 6403 -913 6441 -883
rect 6475 -913 6509 -879
rect 6543 -883 6907 -879
rect 6543 -913 6585 -883
rect 6403 -917 6585 -913
rect 6619 -887 6719 -883
rect 6619 -917 6653 -887
rect 5331 -921 6653 -917
rect 6687 -917 6719 -887
rect 6753 -887 6907 -883
rect 6753 -917 6787 -887
rect 6687 -921 6787 -917
rect 6821 -889 6907 -887
rect 6821 -921 6849 -889
rect 4619 -923 6849 -921
rect 6883 -913 6907 -889
rect 6941 -881 10707 -879
rect 6941 -883 10619 -881
rect 6941 -889 7039 -883
rect 6941 -913 6967 -889
rect 6883 -923 6967 -913
rect 7001 -917 7039 -889
rect 7073 -889 7171 -883
rect 7073 -917 7101 -889
rect 7001 -923 7101 -917
rect 7135 -917 7171 -889
rect 7205 -885 7541 -883
rect 7205 -917 7239 -885
rect 7135 -919 7239 -917
rect 7273 -919 7313 -885
rect 7347 -919 7385 -885
rect 7419 -889 7541 -885
rect 7419 -919 7461 -889
rect 7135 -923 7461 -919
rect 7495 -917 7541 -889
rect 7575 -893 7711 -883
rect 7575 -917 7623 -893
rect 7495 -923 7623 -917
rect 3592 -924 7623 -923
rect 2458 -927 7623 -924
rect 7657 -917 7711 -893
rect 7745 -885 8007 -883
rect 7745 -917 7791 -885
rect 7657 -919 7791 -917
rect 7825 -887 7939 -885
rect 7825 -919 7869 -887
rect 7657 -921 7869 -919
rect 7903 -919 7939 -887
rect 7973 -917 8007 -885
rect 8041 -885 8229 -883
rect 8041 -917 8081 -885
rect 7973 -919 8081 -917
rect 8115 -919 8151 -885
rect 8185 -917 8229 -885
rect 8263 -885 8651 -883
rect 8263 -887 8381 -885
rect 8263 -917 8307 -887
rect 8185 -919 8307 -917
rect 7903 -921 8307 -919
rect 8341 -919 8381 -887
rect 8415 -887 8511 -885
rect 8415 -919 8443 -887
rect 8341 -921 8443 -919
rect 8477 -919 8511 -887
rect 8545 -887 8651 -885
rect 8545 -919 8585 -887
rect 8477 -921 8585 -919
rect 8619 -917 8651 -887
rect 8685 -885 9273 -883
rect 8685 -893 8839 -885
rect 8685 -917 8733 -893
rect 8619 -921 8733 -917
rect 7657 -927 8733 -921
rect 8767 -919 8839 -893
rect 8873 -887 9019 -885
rect 8873 -919 8937 -887
rect 8767 -921 8937 -919
rect 8971 -919 9019 -887
rect 9053 -893 9187 -885
rect 9053 -919 9109 -893
rect 8971 -921 9109 -919
rect 8767 -927 9109 -921
rect 9143 -919 9187 -893
rect 9221 -917 9273 -885
rect 9307 -889 9471 -883
rect 9307 -917 9381 -889
rect 9221 -919 9381 -917
rect 9143 -923 9381 -919
rect 9415 -917 9471 -889
rect 9505 -885 9699 -883
rect 9505 -917 9543 -885
rect 9415 -919 9543 -917
rect 9577 -887 9699 -885
rect 9577 -919 9639 -887
rect 9415 -921 9639 -919
rect 9673 -917 9699 -887
rect 9733 -885 9857 -883
rect 9733 -917 9777 -885
rect 9673 -919 9777 -917
rect 9811 -917 9857 -885
rect 9891 -917 9943 -883
rect 9977 -885 10619 -883
rect 9977 -917 10041 -885
rect 9811 -919 10041 -917
rect 10075 -919 10137 -885
rect 10171 -919 10225 -885
rect 10259 -889 10389 -885
rect 10259 -919 10299 -889
rect 9673 -921 10299 -919
rect 9415 -923 10299 -921
rect 10333 -919 10389 -889
rect 10423 -887 10619 -885
rect 10423 -919 10467 -887
rect 10333 -921 10467 -919
rect 10501 -921 10545 -887
rect 10579 -915 10619 -887
rect 10653 -911 10707 -881
rect 10741 -911 10803 -877
rect 10837 -911 10901 -877
rect 10935 -911 11013 -877
rect 11047 -881 11209 -877
rect 11047 -911 11091 -881
rect 10653 -915 11091 -911
rect 11125 -911 11209 -881
rect 11243 -911 11301 -877
rect 11335 -911 11399 -877
rect 11433 -881 11599 -877
rect 11433 -911 11495 -881
rect 11125 -915 11495 -911
rect 11529 -905 11599 -881
rect 11633 -877 13554 -871
rect 11633 -881 11867 -877
rect 11633 -887 11783 -881
rect 11633 -905 11681 -887
rect 11529 -915 11681 -905
rect 10579 -921 11681 -915
rect 11715 -915 11783 -887
rect 11817 -911 11867 -881
rect 11901 -911 11959 -877
rect 11993 -881 12631 -877
rect 11993 -887 12221 -881
rect 11993 -911 12047 -887
rect 11817 -915 12047 -911
rect 11715 -921 12047 -915
rect 12081 -921 12129 -887
rect 12163 -915 12221 -887
rect 12255 -915 12343 -881
rect 12377 -915 12431 -881
rect 12465 -915 12539 -881
rect 12573 -911 12631 -881
rect 12665 -891 12831 -877
rect 12665 -911 12723 -891
rect 12573 -915 12723 -911
rect 12163 -921 12723 -915
rect 10333 -923 12723 -921
rect 9143 -925 12723 -923
rect 12757 -911 12831 -891
rect 12865 -911 12963 -877
rect 12997 -911 13065 -877
rect 13099 -881 13445 -877
rect 13099 -911 13187 -881
rect 12757 -915 13187 -911
rect 13221 -915 13323 -881
rect 13357 -911 13445 -881
rect 13479 -911 13554 -877
rect 13357 -915 13554 -911
rect 12757 -925 13554 -915
rect 9143 -927 13554 -925
rect 2458 -929 13554 -927
rect -144 -932 13554 -929
rect 742 -934 4410 -932
rect 6056 -934 13554 -932
rect 742 -936 2592 -934
rect 10454 -936 13554 -934
rect 12710 -940 12770 -936
<< viali >>
rect 5797 2367 5831 2401
rect 5927 2371 5961 2405
rect 6071 2371 6105 2405
rect 6219 2373 6253 2407
rect 6363 2373 6397 2407
rect 6503 2371 6537 2405
rect 6659 2375 6693 2409
rect 6799 2371 6833 2405
rect 6947 2375 6981 2409
rect 7085 2371 7119 2405
rect 7215 2371 7249 2405
rect 7357 2373 7391 2407
rect 7485 2373 7519 2407
rect 7623 2371 7657 2405
rect 7755 2369 7789 2403
rect 7913 2373 7947 2407
rect 8065 2375 8099 2409
rect 8215 2373 8249 2407
rect 8329 2379 8363 2413
rect 8479 2375 8513 2409
rect 8623 2375 8657 2409
rect 8763 2375 8797 2409
rect 8907 2375 8941 2409
rect 9065 2375 9099 2409
rect 9225 2379 9259 2413
rect 9421 2387 9455 2421
rect 9609 2389 9643 2423
rect 9773 2383 9807 2417
rect 9951 2383 9985 2417
rect 10119 2387 10153 2421
rect 10287 2387 10321 2421
rect 10451 2389 10485 2423
rect 10587 2387 10621 2421
rect 10769 2387 10803 2421
rect 10921 2373 10955 2407
rect 11133 2393 11167 2427
rect 11357 2397 11391 2431
rect 11547 2397 11581 2431
rect 11725 2383 11759 2417
rect 11820 2376 11852 2410
rect 11852 2376 11854 2410
rect 11892 2376 11920 2410
rect 11920 2376 11926 2410
rect 11964 2376 11988 2410
rect 11988 2376 11998 2410
rect 12036 2376 12056 2410
rect 12056 2376 12070 2410
rect 12108 2376 12124 2410
rect 12124 2376 12142 2410
rect 12180 2376 12192 2410
rect 12192 2376 12214 2410
rect 12252 2376 12260 2410
rect 12260 2376 12286 2410
rect 12324 2376 12328 2410
rect 12328 2376 12358 2410
rect 12396 2376 12430 2410
rect 12468 2376 12498 2410
rect 12498 2376 12502 2410
rect 12540 2376 12566 2410
rect 12566 2376 12574 2410
rect 12612 2376 12634 2410
rect 12634 2376 12646 2410
rect 12684 2376 12702 2410
rect 12702 2376 12718 2410
rect 12756 2376 12770 2410
rect 12770 2376 12790 2410
rect 12828 2376 12838 2410
rect 12838 2376 12862 2410
rect 12900 2376 12906 2410
rect 12906 2376 12934 2410
rect 12972 2376 12974 2410
rect 12974 2376 13006 2410
rect 13044 2376 13076 2410
rect 13076 2376 13078 2410
rect 13116 2376 13144 2410
rect 13144 2376 13150 2410
rect 13188 2376 13212 2410
rect 13212 2376 13222 2410
rect 13260 2376 13280 2410
rect 13280 2376 13294 2410
rect 13332 2376 13348 2410
rect 13348 2376 13366 2410
rect 13404 2376 13416 2410
rect 13416 2376 13438 2410
rect 13476 2376 13484 2410
rect 13484 2376 13510 2410
rect 13548 2376 13552 2410
rect 13552 2376 13582 2410
rect 13620 2376 13654 2410
rect 13692 2376 13722 2410
rect 13722 2376 13726 2410
rect 13764 2376 13790 2410
rect 13790 2376 13798 2410
rect 13836 2376 13858 2410
rect 13858 2376 13870 2410
rect 13908 2376 13926 2410
rect 13926 2376 13942 2410
rect 13980 2376 13994 2410
rect 13994 2376 14014 2410
rect 14052 2376 14062 2410
rect 14062 2376 14086 2410
rect 14124 2376 14130 2410
rect 14130 2376 14158 2410
rect 14196 2376 14198 2410
rect 14198 2376 14230 2410
rect 6150 2150 6184 2184
rect 6222 2150 6256 2184
rect 6294 2150 6328 2184
rect 6366 2150 6400 2184
rect 6438 2150 6472 2184
rect 6510 2150 6544 2184
rect 6582 2150 6616 2184
rect 6654 2150 6688 2184
rect 6726 2150 6760 2184
rect 6798 2150 6832 2184
rect 6870 2150 6904 2184
rect 6942 2150 6976 2184
rect 7014 2150 7048 2184
rect 7086 2150 7120 2184
rect 7158 2150 7192 2184
rect 7230 2150 7264 2184
rect 7302 2150 7336 2184
rect 7374 2150 7408 2184
rect 7446 2150 7480 2184
rect 7518 2150 7552 2184
rect 7590 2150 7624 2184
rect 7662 2150 7696 2184
rect 7734 2150 7768 2184
rect 9428 2172 9462 2206
rect 9500 2172 9534 2206
rect 9572 2172 9606 2206
rect 9644 2172 9678 2206
rect 9716 2172 9750 2206
rect 9788 2172 9822 2206
rect 9860 2172 9894 2206
rect 9932 2172 9966 2206
rect 10004 2172 10038 2206
rect 10076 2172 10110 2206
rect 10148 2172 10182 2206
rect 10220 2172 10254 2206
rect 10292 2172 10326 2206
rect 10364 2172 10398 2206
rect 10436 2172 10470 2206
rect 10508 2172 10542 2206
rect 10580 2172 10614 2206
rect 10652 2172 10686 2206
rect 10724 2172 10758 2206
rect 10796 2172 10830 2206
rect 10868 2172 10902 2206
rect 10940 2172 10974 2206
rect 11012 2172 11046 2206
rect 11084 2172 11118 2206
rect 11156 2172 11190 2206
rect 11228 2172 11262 2206
rect 11300 2172 11334 2206
rect 11372 2172 11406 2206
rect 11444 2172 11478 2206
rect 11516 2172 11550 2206
rect 12002 2170 12036 2204
rect 12074 2170 12108 2204
rect 12146 2170 12180 2204
rect 12218 2170 12252 2204
rect 12290 2170 12324 2204
rect 12362 2170 12396 2204
rect 12434 2170 12468 2204
rect 12506 2170 12540 2204
rect 12578 2170 12612 2204
rect 12650 2170 12684 2204
rect 12722 2170 12756 2204
rect 12794 2170 12828 2204
rect 12866 2170 12900 2204
rect 12938 2170 12972 2204
rect 13010 2170 13044 2204
rect 13082 2170 13116 2204
rect 13154 2170 13188 2204
rect 13226 2170 13260 2204
rect 13298 2170 13332 2204
rect 13370 2170 13404 2204
rect 13442 2170 13476 2204
rect 13514 2170 13548 2204
rect 13586 2170 13620 2204
rect 13658 2170 13692 2204
rect 13730 2170 13764 2204
rect 13802 2170 13836 2204
rect 13874 2170 13908 2204
rect 13946 2170 13980 2204
rect 14018 2170 14052 2204
rect 14090 2170 14124 2204
rect 2751 2095 2785 2129
rect 2885 2097 2919 2131
rect 3045 2095 3079 2129
rect 3219 2097 3253 2131
rect 3367 2095 3401 2129
rect 3519 2097 3553 2131
rect 3655 2095 3689 2129
rect 3791 2097 3825 2131
rect 3943 2095 3977 2129
rect 4101 2097 4135 2131
rect 4269 2101 4303 2135
rect 4427 2097 4461 2131
rect 4603 2095 4637 2129
rect 4765 2097 4799 2131
rect 3030 1866 3064 1900
rect 3102 1866 3136 1900
rect 3174 1866 3208 1900
rect 3246 1866 3280 1900
rect 3318 1866 3352 1900
rect 3390 1866 3424 1900
rect 3462 1866 3496 1900
rect 3534 1866 3568 1900
rect 3606 1866 3640 1900
rect 3678 1866 3712 1900
rect 3750 1866 3784 1900
rect 3822 1866 3856 1900
rect 3894 1866 3928 1900
rect 3966 1866 4000 1900
rect 4038 1866 4072 1900
rect 4110 1866 4144 1900
rect 4182 1866 4216 1900
rect 4254 1866 4288 1900
rect 4326 1866 4360 1900
rect 4398 1866 4432 1900
rect 4470 1866 4504 1900
rect 4542 1866 4576 1900
rect 4614 1866 4648 1900
rect 800 562 834 596
rect 922 558 956 592
rect 1042 562 1076 596
rect 1164 558 1198 592
rect 1274 564 1308 598
rect 1384 560 1418 594
rect 1506 560 1540 594
rect 1638 560 1672 594
rect 1757 562 1791 596
rect 1881 562 1915 596
rect 2007 562 2041 596
rect 2123 564 2157 598
rect 2251 566 2285 600
rect 2383 560 2417 594
rect 2521 564 2555 598
rect 2623 560 2657 594
rect 5594 484 5628 518
rect 5666 484 5700 518
rect 5738 484 5772 518
rect 5810 484 5844 518
rect 5882 484 5916 518
rect 8046 498 8080 532
rect 8118 498 8152 532
rect 8190 498 8224 532
rect 8262 498 8296 532
rect 8334 498 8368 532
rect 1158 344 1192 378
rect 1230 344 1264 378
rect 1302 344 1336 378
rect 1374 344 1408 378
rect 1446 344 1480 378
rect 5702 370 5736 404
rect 5774 370 5808 404
rect 8154 384 8188 418
rect 8226 384 8260 418
rect 11101 410 11135 444
rect 11173 410 11207 444
rect 11245 410 11279 444
rect 11317 410 11351 444
rect 11389 410 11423 444
rect 11461 410 11495 444
rect 11533 410 11567 444
rect 11605 410 11639 444
rect 11677 410 11711 444
rect 11749 410 11783 444
rect 11821 410 11855 444
rect 11893 410 11927 444
rect 11965 410 11999 444
rect 12037 410 12071 444
rect 12109 410 12143 444
rect 12181 410 12215 444
rect 12253 410 12287 444
rect 12325 410 12359 444
rect 12397 410 12431 444
rect 12469 410 12503 444
rect 12541 410 12575 444
rect 12613 410 12647 444
rect 12685 410 12719 444
rect 12757 410 12791 444
rect 12829 410 12863 444
rect 12901 410 12935 444
rect 12973 410 13007 444
rect 13045 410 13079 444
rect 13117 410 13151 444
rect 13189 410 13223 444
rect 2128 336 2162 370
rect 2200 336 2234 370
rect 2272 336 2306 370
rect 2344 336 2378 370
rect 2416 336 2450 370
rect 5902 306 5936 340
rect 8354 320 8388 354
rect 1266 230 1300 264
rect 1338 230 1372 264
rect 2236 222 2270 256
rect 2308 222 2342 256
rect 1138 186 1172 220
rect 3511 216 3545 250
rect 5702 242 5736 276
rect 5774 242 5808 276
rect 8154 256 8188 290
rect 8226 256 8260 290
rect 2108 178 2142 212
rect 1266 142 1300 176
rect 1338 142 1372 176
rect 3414 172 3448 206
rect 2236 134 2270 168
rect 2308 134 2342 168
rect 3511 128 3545 162
rect 3439 14 3473 48
rect 3511 14 3545 48
rect 3583 14 3617 48
rect 11049 -142 11083 -108
rect 11121 -142 11155 -108
rect 11193 -142 11227 -108
rect 11265 -142 11299 -108
rect 11337 -142 11371 -108
rect 11409 -142 11443 -108
rect 11481 -142 11515 -108
rect 11553 -142 11587 -108
rect 11625 -142 11659 -108
rect 11697 -142 11731 -108
rect 11769 -142 11803 -108
rect 11841 -142 11875 -108
rect 11913 -142 11947 -108
rect 11985 -142 12019 -108
rect 12057 -142 12091 -108
rect 12129 -142 12163 -108
rect 12201 -142 12235 -108
rect 12273 -142 12307 -108
rect 12345 -142 12379 -108
rect 12417 -142 12451 -108
rect 12489 -142 12523 -108
rect 12561 -142 12595 -108
rect 12633 -142 12667 -108
rect 12705 -142 12739 -108
rect 12777 -142 12811 -108
rect 12849 -142 12883 -108
rect 12921 -142 12955 -108
rect 12993 -142 13027 -108
rect 13065 -142 13099 -108
rect 13137 -142 13171 -108
rect 13209 -142 13243 -108
rect 13281 -142 13315 -108
rect 13353 -142 13387 -108
rect 10946 -227 10980 -193
rect 10946 -299 10980 -265
rect 10946 -371 10980 -337
rect 319 -482 353 -448
rect 3945 -456 3979 -422
rect 4713 -448 4747 -414
rect 4785 -448 4819 -414
rect 4857 -448 4891 -414
rect 4929 -448 4963 -414
rect 5001 -448 5035 -414
rect 5073 -448 5107 -414
rect 5145 -448 5179 -414
rect 5217 -448 5251 -414
rect 5289 -448 5323 -414
rect 5361 -448 5395 -414
rect 5433 -448 5467 -414
rect 5505 -448 5539 -414
rect 5577 -448 5611 -414
rect 5649 -448 5683 -414
rect 5931 -448 5965 -414
rect 6003 -448 6037 -414
rect 6075 -448 6109 -414
rect 6147 -448 6181 -414
rect 6219 -448 6253 -414
rect 6291 -448 6325 -414
rect 6363 -448 6397 -414
rect 6435 -448 6469 -414
rect 6507 -448 6541 -414
rect 6579 -448 6613 -414
rect 6651 -448 6685 -414
rect 6723 -448 6757 -414
rect 6795 -448 6829 -414
rect 6867 -448 6901 -414
rect 7831 -446 7865 -412
rect 7903 -446 7937 -412
rect 7975 -446 8009 -412
rect 8047 -446 8081 -412
rect 8119 -446 8153 -412
rect 8191 -446 8225 -412
rect 8263 -446 8297 -412
rect 8335 -446 8369 -412
rect 8407 -446 8441 -412
rect 8479 -446 8513 -412
rect 8551 -446 8585 -412
rect 8623 -446 8657 -412
rect 8695 -446 8729 -412
rect 8767 -446 8801 -412
rect 9049 -446 9083 -412
rect 9121 -446 9155 -412
rect 9193 -446 9227 -412
rect 9265 -446 9299 -412
rect 9337 -446 9371 -412
rect 9409 -446 9443 -412
rect 9481 -446 9515 -412
rect 9553 -446 9587 -412
rect 9625 -446 9659 -412
rect 9697 -446 9731 -412
rect 9769 -446 9803 -412
rect 9841 -446 9875 -412
rect 9913 -446 9947 -412
rect 9985 -446 10019 -412
rect 10946 -443 10980 -409
rect 2178 -514 2212 -480
rect 319 -570 353 -536
rect 3945 -544 3979 -510
rect 5742 -527 5776 -493
rect 5838 -527 5872 -493
rect 6954 -527 6988 -493
rect 7744 -525 7778 -491
rect 8854 -525 8888 -491
rect 8962 -525 8996 -491
rect 10946 -515 10980 -481
rect 4713 -606 4747 -572
rect 4785 -606 4819 -572
rect 4857 -606 4891 -572
rect 4929 -606 4963 -572
rect 5001 -606 5035 -572
rect 5073 -606 5107 -572
rect 5145 -606 5179 -572
rect 5217 -606 5251 -572
rect 5289 -606 5323 -572
rect 5361 -606 5395 -572
rect 5433 -606 5467 -572
rect 5505 -606 5539 -572
rect 5577 -606 5611 -572
rect 5649 -606 5683 -572
rect 5931 -606 5965 -572
rect 6003 -606 6037 -572
rect 6075 -606 6109 -572
rect 6147 -606 6181 -572
rect 6219 -606 6253 -572
rect 6291 -606 6325 -572
rect 6363 -606 6397 -572
rect 6435 -606 6469 -572
rect 6507 -606 6541 -572
rect 6579 -606 6613 -572
rect 6651 -606 6685 -572
rect 6723 -606 6757 -572
rect 6795 -606 6829 -572
rect 6867 -606 6901 -572
rect 7831 -604 7865 -570
rect 7903 -604 7937 -570
rect 7975 -604 8009 -570
rect 8047 -604 8081 -570
rect 8119 -604 8153 -570
rect 8191 -604 8225 -570
rect 8263 -604 8297 -570
rect 8335 -604 8369 -570
rect 8407 -604 8441 -570
rect 8479 -604 8513 -570
rect 8551 -604 8585 -570
rect 8623 -604 8657 -570
rect 8695 -604 8729 -570
rect 8767 -604 8801 -570
rect 9049 -604 9083 -570
rect 9121 -604 9155 -570
rect 9193 -604 9227 -570
rect 9265 -604 9299 -570
rect 9337 -604 9371 -570
rect 9409 -604 9443 -570
rect 9481 -604 9515 -570
rect 9553 -604 9587 -570
rect 9625 -604 9659 -570
rect 9697 -604 9731 -570
rect 9769 -604 9803 -570
rect 9841 -604 9875 -570
rect 9913 -604 9947 -570
rect 9985 -604 10019 -570
rect 11049 -600 11083 -566
rect 11121 -600 11155 -566
rect 11193 -600 11227 -566
rect 11265 -600 11299 -566
rect 11337 -600 11371 -566
rect 11409 -600 11443 -566
rect 11481 -600 11515 -566
rect 11553 -600 11587 -566
rect 11625 -600 11659 -566
rect 11697 -600 11731 -566
rect 11769 -600 11803 -566
rect 11841 -600 11875 -566
rect 11913 -600 11947 -566
rect 11985 -600 12019 -566
rect 12057 -600 12091 -566
rect 12129 -600 12163 -566
rect 12201 -600 12235 -566
rect 12273 -600 12307 -566
rect 12345 -600 12379 -566
rect 12417 -600 12451 -566
rect 12489 -600 12523 -566
rect 12561 -600 12595 -566
rect 12633 -600 12667 -566
rect 12705 -600 12739 -566
rect 12777 -600 12811 -566
rect 12849 -600 12883 -566
rect 12921 -600 12955 -566
rect 12993 -600 13027 -566
rect 13065 -600 13099 -566
rect 13137 -600 13171 -566
rect 13209 -600 13243 -566
rect 13281 -600 13315 -566
rect 13353 -600 13387 -566
rect 247 -684 281 -650
rect 319 -684 353 -650
rect 391 -684 425 -650
rect 1210 -676 1244 -642
rect 1282 -676 1316 -642
rect 1354 -676 1388 -642
rect 1426 -676 1460 -642
rect 2190 -672 2224 -638
rect 2262 -672 2296 -638
rect 2334 -672 2368 -638
rect 2406 -672 2440 -638
rect 3083 -666 3117 -632
rect 3155 -666 3189 -632
rect 3227 -666 3261 -632
rect 3873 -658 3907 -624
rect 3945 -658 3979 -624
rect 4017 -658 4051 -624
rect 4638 -720 4672 -686
rect 4710 -720 4744 -686
rect 4782 -720 4816 -686
rect 4854 -720 4888 -686
rect 4926 -720 4960 -686
rect 4998 -720 5032 -686
rect 5070 -720 5104 -686
rect 5142 -720 5176 -686
rect 5214 -720 5248 -686
rect 5286 -720 5320 -686
rect 5358 -720 5392 -686
rect 5430 -720 5464 -686
rect 5502 -720 5536 -686
rect 5574 -720 5608 -686
rect 5646 -720 5680 -686
rect 5718 -720 5752 -686
rect 5790 -720 5824 -686
rect 5862 -720 5896 -686
rect 5934 -720 5968 -686
rect 6006 -720 6040 -686
rect 6078 -720 6112 -686
rect 6150 -720 6184 -686
rect 6222 -720 6256 -686
rect 6294 -720 6328 -686
rect 6366 -720 6400 -686
rect 6438 -720 6472 -686
rect 6510 -720 6544 -686
rect 6582 -720 6616 -686
rect 6654 -720 6688 -686
rect 6726 -720 6760 -686
rect 6798 -720 6832 -686
rect 6870 -720 6904 -686
rect 6942 -720 6976 -686
rect 7756 -718 7790 -684
rect 7828 -718 7862 -684
rect 7900 -718 7934 -684
rect 7972 -718 8006 -684
rect 8044 -718 8078 -684
rect 8116 -718 8150 -684
rect 8188 -718 8222 -684
rect 8260 -718 8294 -684
rect 8332 -718 8366 -684
rect 8404 -718 8438 -684
rect 8476 -718 8510 -684
rect 8548 -718 8582 -684
rect 8620 -718 8654 -684
rect 8692 -718 8726 -684
rect 8764 -718 8798 -684
rect 8836 -718 8870 -684
rect 8908 -718 8942 -684
rect 8980 -718 9014 -684
rect 9052 -718 9086 -684
rect 9124 -718 9158 -684
rect 9196 -718 9230 -684
rect 9268 -718 9302 -684
rect 9340 -718 9374 -684
rect 9412 -718 9446 -684
rect 9484 -718 9518 -684
rect 9556 -718 9590 -684
rect 9628 -718 9662 -684
rect 9700 -718 9734 -684
rect 9772 -718 9806 -684
rect 9844 -718 9878 -684
rect 9916 -718 9950 -684
rect 9988 -718 10022 -684
rect 10060 -718 10094 -684
rect 10941 -714 10975 -680
rect 11013 -714 11047 -680
rect 11085 -714 11119 -680
rect 11157 -714 11191 -680
rect 11229 -714 11263 -680
rect 11301 -714 11335 -680
rect 11373 -714 11407 -680
rect 11445 -714 11479 -680
rect 11517 -714 11551 -680
rect 11589 -714 11623 -680
rect 11661 -714 11695 -680
rect 11733 -714 11767 -680
rect 11805 -714 11839 -680
rect 11877 -714 11911 -680
rect 11949 -714 11983 -680
rect 12021 -714 12055 -680
rect 12093 -714 12127 -680
rect 12165 -714 12199 -680
rect 12237 -714 12271 -680
rect 12309 -714 12343 -680
rect 12381 -714 12415 -680
rect 12453 -714 12487 -680
rect 12525 -714 12559 -680
rect 12597 -714 12631 -680
rect 12669 -714 12703 -680
rect 12741 -714 12775 -680
rect 12813 -714 12847 -680
rect 12885 -714 12919 -680
rect 12957 -714 12991 -680
rect 13029 -714 13063 -680
rect 13101 -714 13135 -680
rect 13173 -714 13207 -680
rect 13245 -714 13279 -680
rect 13317 -714 13351 -680
rect 13389 -714 13423 -680
rect 13461 -714 13495 -680
rect -123 -922 -89 -888
rect 27 -922 61 -888
rect 185 -920 219 -886
rect 333 -922 367 -888
rect 483 -922 517 -888
rect 629 -922 663 -888
rect 716 -921 750 -887
rect 846 -925 880 -891
rect 984 -921 1018 -887
rect 1126 -923 1160 -889
rect 1268 -927 1302 -893
rect 1414 -923 1448 -889
rect 1556 -921 1590 -887
rect 1728 -921 1762 -887
rect 1896 -925 1930 -891
rect 2050 -923 2084 -889
rect 2198 -923 2232 -889
rect 2340 -923 2374 -889
rect 2510 -923 2544 -889
rect 2702 -918 2736 -884
rect 2870 -918 2904 -884
rect 3042 -918 3076 -884
rect 3220 -918 3254 -884
rect 3392 -920 3426 -886
rect 3558 -924 3592 -890
rect 3742 -920 3776 -886
rect 3912 -920 3946 -886
rect 4072 -918 4106 -884
rect 4252 -918 4286 -884
rect 4393 -917 4427 -883
rect 4517 -917 4551 -883
rect 4647 -911 4681 -877
rect 4785 -911 4819 -877
rect 4921 -911 4955 -877
rect 5063 -911 5097 -877
rect 5221 -917 5255 -883
rect 5389 -917 5423 -883
rect 5551 -911 5585 -877
rect 5691 -917 5725 -883
rect 5845 -913 5879 -879
rect 6001 -911 6035 -877
rect 6151 -917 6185 -883
rect 6293 -913 6327 -879
rect 6441 -913 6475 -879
rect 6585 -917 6619 -883
rect 6719 -917 6753 -883
rect 6849 -923 6883 -889
rect 6967 -923 7001 -889
rect 7101 -923 7135 -889
rect 7239 -919 7273 -885
rect 7385 -919 7419 -885
rect 7541 -917 7575 -883
rect 7711 -917 7745 -883
rect 7869 -921 7903 -887
rect 8007 -917 8041 -883
rect 8151 -919 8185 -885
rect 8307 -921 8341 -887
rect 8443 -921 8477 -887
rect 8585 -921 8619 -887
rect 8733 -927 8767 -893
rect 8937 -921 8971 -887
rect 9109 -927 9143 -893
rect 9273 -917 9307 -883
rect 9471 -917 9505 -883
rect 9639 -921 9673 -887
rect 9777 -919 9811 -885
rect 9943 -917 9977 -883
rect 10137 -919 10171 -885
rect 10299 -923 10333 -889
rect 10467 -921 10501 -887
rect 10619 -915 10653 -881
rect 10803 -911 10837 -877
rect 11013 -911 11047 -877
rect 11209 -911 11243 -877
rect 11399 -911 11433 -877
rect 11599 -905 11633 -871
rect 11783 -915 11817 -881
rect 11959 -911 11993 -877
rect 12129 -921 12163 -887
rect 12343 -915 12377 -881
rect 12539 -915 12573 -881
rect 12723 -925 12757 -891
rect 12963 -911 12997 -877
rect 13187 -915 13221 -881
rect 13445 -911 13479 -877
<< metal1 >>
rect 2518 2908 2984 3042
rect 2518 2728 2661 2908
rect 2841 2728 2984 2908
rect 2518 2188 2984 2728
rect 4296 2306 4552 2566
rect 11856 2474 14386 2476
rect 9040 2470 14386 2474
rect 5700 2466 8116 2468
rect 4866 2464 8116 2466
rect 8834 2464 14386 2470
rect 4866 2431 14386 2464
rect 4866 2427 11357 2431
rect 4866 2423 11133 2427
rect 4866 2421 9609 2423
rect 4866 2413 9421 2421
rect 4866 2409 8329 2413
rect 4866 2407 6659 2409
rect 4866 2405 6219 2407
rect 4866 2401 5927 2405
rect 4866 2367 5797 2401
rect 5831 2371 5927 2401
rect 5961 2371 6071 2405
rect 6105 2373 6219 2405
rect 6253 2373 6363 2407
rect 6397 2405 6659 2407
rect 6397 2373 6503 2405
rect 6105 2371 6503 2373
rect 6537 2375 6659 2405
rect 6693 2405 6947 2409
rect 6693 2375 6799 2405
rect 6537 2371 6799 2375
rect 6833 2375 6947 2405
rect 6981 2407 8065 2409
rect 6981 2405 7357 2407
rect 6981 2375 7085 2405
rect 6833 2371 7085 2375
rect 7119 2371 7215 2405
rect 7249 2373 7357 2405
rect 7391 2373 7485 2407
rect 7519 2405 7913 2407
rect 7519 2373 7623 2405
rect 7249 2371 7623 2373
rect 7657 2403 7913 2405
rect 7657 2371 7755 2403
rect 5831 2369 7755 2371
rect 7789 2373 7913 2403
rect 7947 2375 8065 2407
rect 8099 2407 8329 2409
rect 8099 2375 8215 2407
rect 7947 2373 8215 2375
rect 8249 2379 8329 2407
rect 8363 2409 9225 2413
rect 8363 2379 8479 2409
rect 8249 2375 8479 2379
rect 8513 2375 8623 2409
rect 8657 2375 8763 2409
rect 8797 2375 8907 2409
rect 8941 2375 9065 2409
rect 9099 2379 9225 2409
rect 9259 2387 9421 2413
rect 9455 2389 9609 2421
rect 9643 2421 10451 2423
rect 9643 2417 10119 2421
rect 9643 2389 9773 2417
rect 9455 2387 9773 2389
rect 9259 2383 9773 2387
rect 9807 2383 9951 2417
rect 9985 2387 10119 2417
rect 10153 2387 10287 2421
rect 10321 2389 10451 2421
rect 10485 2421 11133 2423
rect 10485 2389 10587 2421
rect 10321 2387 10587 2389
rect 10621 2387 10769 2421
rect 10803 2407 11133 2421
rect 10803 2387 10921 2407
rect 9985 2383 10921 2387
rect 9259 2379 10921 2383
rect 9099 2375 10921 2379
rect 8249 2373 10921 2375
rect 10955 2393 11133 2407
rect 11167 2397 11357 2427
rect 11391 2397 11547 2431
rect 11581 2417 14386 2431
rect 11581 2397 11725 2417
rect 11167 2393 11725 2397
rect 10955 2383 11725 2393
rect 11759 2410 14386 2417
rect 11759 2383 11820 2410
rect 10955 2376 11820 2383
rect 11854 2376 11892 2410
rect 11926 2376 11964 2410
rect 11998 2376 12036 2410
rect 12070 2376 12108 2410
rect 12142 2376 12180 2410
rect 12214 2376 12252 2410
rect 12286 2376 12324 2410
rect 12358 2376 12396 2410
rect 12430 2376 12468 2410
rect 12502 2376 12540 2410
rect 12574 2376 12612 2410
rect 12646 2376 12684 2410
rect 12718 2376 12756 2410
rect 12790 2376 12828 2410
rect 12862 2376 12900 2410
rect 12934 2376 12972 2410
rect 13006 2376 13044 2410
rect 13078 2376 13116 2410
rect 13150 2376 13188 2410
rect 13222 2376 13260 2410
rect 13294 2376 13332 2410
rect 13366 2376 13404 2410
rect 13438 2376 13476 2410
rect 13510 2376 13548 2410
rect 13582 2376 13620 2410
rect 13654 2376 13692 2410
rect 13726 2376 13764 2410
rect 13798 2376 13836 2410
rect 13870 2376 13908 2410
rect 13942 2376 13980 2410
rect 14014 2376 14052 2410
rect 14086 2376 14124 2410
rect 14158 2376 14196 2410
rect 14230 2376 14386 2410
rect 10955 2373 14386 2376
rect 7789 2369 14386 2373
rect 5831 2367 14386 2369
rect 4866 2312 14386 2367
rect 4866 2308 8116 2312
rect 8834 2310 14386 2312
rect 8834 2308 9144 2310
rect 4866 2188 5734 2308
rect 2518 2178 5734 2188
rect 2668 2168 5734 2178
rect 6100 2184 7810 2308
rect 2668 2135 4898 2168
rect 6100 2150 6150 2184
rect 6184 2150 6222 2184
rect 6256 2150 6294 2184
rect 6328 2150 6366 2184
rect 6400 2150 6438 2184
rect 6472 2150 6510 2184
rect 6544 2150 6582 2184
rect 6616 2150 6654 2184
rect 6688 2150 6726 2184
rect 6760 2150 6798 2184
rect 6832 2150 6870 2184
rect 6904 2150 6942 2184
rect 6976 2150 7014 2184
rect 7048 2150 7086 2184
rect 7120 2150 7158 2184
rect 7192 2150 7230 2184
rect 7264 2150 7302 2184
rect 7336 2150 7374 2184
rect 7408 2150 7446 2184
rect 7480 2150 7518 2184
rect 7552 2150 7590 2184
rect 7624 2150 7662 2184
rect 7696 2150 7734 2184
rect 7768 2150 7810 2184
rect 6100 2138 7810 2150
rect 2668 2131 4269 2135
rect 2668 2129 2885 2131
rect 2668 2095 2751 2129
rect 2785 2097 2885 2129
rect 2919 2129 3219 2131
rect 2919 2097 3045 2129
rect 2785 2095 3045 2097
rect 3079 2097 3219 2129
rect 3253 2129 3519 2131
rect 3253 2097 3367 2129
rect 3079 2095 3367 2097
rect 3401 2097 3519 2129
rect 3553 2129 3791 2131
rect 3553 2097 3655 2129
rect 3401 2095 3655 2097
rect 3689 2097 3791 2129
rect 3825 2129 4101 2131
rect 3825 2097 3943 2129
rect 3689 2095 3943 2097
rect 3977 2097 4101 2129
rect 4135 2101 4269 2131
rect 4303 2131 4898 2135
rect 4303 2101 4427 2131
rect 4135 2097 4427 2101
rect 4461 2129 4765 2131
rect 4461 2097 4603 2129
rect 3977 2095 4603 2097
rect 4637 2097 4765 2129
rect 4799 2097 4898 2131
rect 6206 2104 7714 2138
rect 4637 2095 4898 2097
rect 2668 2026 4898 2095
rect 6192 2074 7714 2104
rect 6210 2070 7714 2074
rect 6210 2035 6221 2070
rect 7690 2048 7714 2070
rect 7690 2036 7704 2048
rect 7679 2035 7704 2036
rect -740 1715 -274 1849
rect -740 1535 -597 1715
rect -417 1535 -274 1715
rect -740 1383 -274 1535
rect -740 700 382 834
rect -740 520 -597 700
rect -417 520 382 700
rect 694 626 1746 628
rect 2668 626 2744 2026
rect 2988 1900 4694 2026
rect 2988 1866 3030 1900
rect 3064 1866 3102 1900
rect 3136 1866 3174 1900
rect 3208 1866 3246 1900
rect 3280 1866 3318 1900
rect 3352 1866 3390 1900
rect 3424 1866 3462 1900
rect 3496 1866 3534 1900
rect 3568 1866 3606 1900
rect 3640 1866 3678 1900
rect 3712 1866 3750 1900
rect 3784 1866 3822 1900
rect 3856 1866 3894 1900
rect 3928 1866 3966 1900
rect 4000 1866 4038 1900
rect 4072 1866 4110 1900
rect 4144 1866 4182 1900
rect 4216 1866 4254 1900
rect 4288 1866 4326 1900
rect 4360 1866 4398 1900
rect 4432 1866 4470 1900
rect 4504 1866 4542 1900
rect 4576 1866 4614 1900
rect 4648 1866 4694 1900
rect 2988 1852 4694 1866
rect 3086 1796 4588 1852
rect 2982 1724 3054 1758
rect 3086 1726 4596 1796
rect 2982 756 3008 1724
rect 3042 756 3054 1724
rect 2982 740 3054 756
rect 4630 1154 4716 1756
rect 5768 1702 6152 2030
rect 6210 2028 7704 2035
rect 6210 2026 6722 2028
rect 6220 2022 6722 2026
rect 7500 2024 7704 2028
rect 5730 1154 6152 1702
rect 4630 1040 6152 1154
rect 4630 1010 6000 1040
rect 6082 1038 6152 1040
rect 7472 1020 7704 1024
rect 6208 1012 7704 1020
rect 6208 1011 6221 1012
rect 4630 746 4994 1010
rect 6208 977 6210 1011
rect 7662 977 7704 1012
rect 6208 974 7704 977
rect 4584 740 4994 746
rect 2982 732 4994 740
rect 6204 958 7704 974
rect 5558 736 5962 738
rect 6204 736 7712 958
rect 2982 728 4680 732
rect 2982 694 3101 728
rect 4577 694 4680 728
rect 2982 682 4680 694
rect 2982 658 4604 682
rect 694 600 2784 626
rect 694 598 2251 600
rect 694 596 1274 598
rect 694 562 800 596
rect 834 592 1042 596
rect 834 562 922 592
rect 694 558 922 562
rect 956 562 1042 592
rect 1076 592 1274 596
rect 1076 562 1164 592
rect 956 558 1164 562
rect 1198 564 1274 592
rect 1308 596 2123 598
rect 1308 594 1757 596
rect 1308 564 1384 594
rect 1198 560 1384 564
rect 1418 560 1506 594
rect 1540 560 1638 594
rect 1672 562 1757 594
rect 1791 562 1881 596
rect 1915 562 2007 596
rect 2041 564 2123 596
rect 2157 566 2251 598
rect 2285 598 2784 600
rect 2285 594 2521 598
rect 2285 566 2383 594
rect 2157 564 2383 566
rect 2041 562 2383 564
rect 1672 560 2383 562
rect 2417 564 2521 594
rect 2555 594 2784 598
rect 2555 564 2623 594
rect 2417 560 2623 564
rect 2657 560 2784 594
rect 1198 558 2784 560
rect 694 526 2784 558
rect 694 524 776 526
rect 694 520 764 524
rect -740 368 382 520
rect -740 -200 -274 -66
rect -740 -380 -597 -200
rect -417 -380 -274 -200
rect -740 -532 -274 -380
rect 292 -150 382 368
rect 1118 378 1518 526
rect 1728 524 2784 526
rect 1118 344 1158 378
rect 1192 344 1230 378
rect 1264 344 1302 378
rect 1336 344 1374 378
rect 1408 344 1446 378
rect 1480 344 1518 378
rect 1118 332 1518 344
rect 2092 370 2488 524
rect 2092 336 2128 370
rect 2162 336 2200 370
rect 2234 336 2272 370
rect 2306 336 2344 370
rect 2378 336 2416 370
rect 2450 336 2488 370
rect 1220 264 1420 332
rect 2092 322 2488 336
rect 886 220 1180 236
rect 886 186 1138 220
rect 1172 186 1180 220
rect 1220 230 1266 264
rect 1300 230 1338 264
rect 1372 230 1420 264
rect 2188 256 2390 322
rect 1220 216 1420 230
rect 1812 212 2158 230
rect 2188 222 2236 256
rect 2270 222 2308 256
rect 2342 222 2390 256
rect 2188 214 2390 222
rect 2720 226 2784 524
rect 3484 262 3576 658
rect 5558 546 8418 736
rect 5558 518 5962 546
rect 5558 484 5594 518
rect 5628 484 5666 518
rect 5700 484 5738 518
rect 5772 484 5810 518
rect 5844 484 5882 518
rect 5916 484 5962 518
rect 5558 466 5962 484
rect 8004 532 8418 546
rect 9060 618 9144 2308
rect 9396 2206 11592 2310
rect 11856 2298 14386 2310
rect 9396 2172 9428 2206
rect 9462 2172 9500 2206
rect 9534 2172 9572 2206
rect 9606 2172 9644 2206
rect 9678 2172 9716 2206
rect 9750 2172 9788 2206
rect 9822 2172 9860 2206
rect 9894 2172 9932 2206
rect 9966 2172 10004 2206
rect 10038 2172 10076 2206
rect 10110 2172 10148 2206
rect 10182 2172 10220 2206
rect 10254 2172 10292 2206
rect 10326 2172 10364 2206
rect 10398 2172 10436 2206
rect 10470 2172 10508 2206
rect 10542 2172 10580 2206
rect 10614 2172 10652 2206
rect 10686 2172 10724 2206
rect 10758 2172 10796 2206
rect 10830 2172 10868 2206
rect 10902 2172 10940 2206
rect 10974 2172 11012 2206
rect 11046 2172 11084 2206
rect 11118 2172 11156 2206
rect 11190 2172 11228 2206
rect 11262 2172 11300 2206
rect 11334 2172 11372 2206
rect 11406 2172 11444 2206
rect 11478 2172 11516 2206
rect 11550 2172 11592 2206
rect 9396 2158 11592 2172
rect 11962 2204 14172 2298
rect 11962 2170 12002 2204
rect 12036 2170 12074 2204
rect 12108 2170 12146 2204
rect 12180 2170 12218 2204
rect 12252 2170 12290 2204
rect 12324 2170 12362 2204
rect 12396 2170 12434 2204
rect 12468 2170 12506 2204
rect 12540 2170 12578 2204
rect 12612 2170 12650 2204
rect 12684 2170 12722 2204
rect 12756 2170 12794 2204
rect 12828 2170 12866 2204
rect 12900 2170 12938 2204
rect 12972 2170 13010 2204
rect 13044 2170 13082 2204
rect 13116 2170 13154 2204
rect 13188 2170 13226 2204
rect 13260 2170 13298 2204
rect 13332 2170 13370 2204
rect 13404 2170 13442 2204
rect 13476 2170 13514 2204
rect 13548 2170 13586 2204
rect 13620 2170 13658 2204
rect 13692 2170 13730 2204
rect 13764 2170 13802 2204
rect 13836 2170 13874 2204
rect 13908 2170 13946 2204
rect 13980 2170 14018 2204
rect 14052 2170 14090 2204
rect 14124 2170 14172 2204
rect 9488 2140 11494 2158
rect 11962 2146 14172 2170
rect 9488 2092 11450 2140
rect 9488 2058 9501 2092
rect 12056 2090 14062 2146
rect 9488 2046 11450 2058
rect 12056 2056 12075 2090
rect 14051 2056 14062 2090
rect 12056 2048 14062 2056
rect 9342 2040 9430 2044
rect 9228 1867 9430 2040
rect 12056 2038 14056 2048
rect 9228 1815 9289 1867
rect 9341 1815 9430 1867
rect 9228 1803 9430 1815
rect 9228 1751 9289 1803
rect 9341 1751 9430 1803
rect 9228 1684 9430 1751
rect 14096 2028 14206 2052
rect 14096 1700 14110 2028
rect 14018 1660 14110 1700
rect 14144 1660 14206 2028
rect 14018 1646 14206 1660
rect 9574 1634 11308 1646
rect 12330 1632 14206 1646
rect 9574 1538 11308 1600
rect 14051 1598 14206 1632
rect 9574 1432 11436 1538
rect 12330 1536 14206 1598
rect 12330 1522 14172 1536
rect 12330 1464 14068 1522
rect 9574 1406 11492 1432
rect 9486 1294 11492 1406
rect 12060 1294 14068 1464
rect 9486 1134 14120 1294
rect 9486 1018 10128 1134
rect 10244 1018 14120 1134
rect 9486 968 14120 1018
rect 9492 966 14120 968
rect 11172 878 14120 966
rect 12186 636 12298 878
rect 12430 646 12542 878
rect 12692 646 12804 878
rect 13192 838 14120 878
rect 10674 618 11130 620
rect 9060 546 11130 618
rect 9060 542 10926 546
rect 8004 498 8046 532
rect 8080 498 8118 532
rect 8152 498 8190 532
rect 8224 498 8262 532
rect 8296 498 8334 532
rect 8368 498 8418 532
rect 8004 482 8418 498
rect 5652 404 5856 466
rect 5652 370 5702 404
rect 5736 370 5774 404
rect 5808 370 5856 404
rect 5652 354 5856 370
rect 6072 356 6498 430
rect 8104 418 8310 482
rect 11218 458 11330 558
rect 11450 458 11562 556
rect 13190 554 13248 616
rect 11674 458 11786 542
rect 11080 456 13250 458
rect 8104 384 8154 418
rect 8188 384 8226 418
rect 8260 384 8310 418
rect 11078 444 13250 456
rect 11078 410 11101 444
rect 11135 410 11173 444
rect 11207 410 11245 444
rect 11279 410 11317 444
rect 11351 410 11389 444
rect 11423 410 11461 444
rect 11495 410 11533 444
rect 11567 410 11605 444
rect 11639 410 11677 444
rect 11711 410 11749 444
rect 11783 410 11821 444
rect 11855 410 11893 444
rect 11927 410 11965 444
rect 11999 410 12037 444
rect 12071 410 12109 444
rect 12143 410 12181 444
rect 12215 410 12253 444
rect 12287 410 12325 444
rect 12359 410 12397 444
rect 12431 410 12469 444
rect 12503 410 12541 444
rect 12575 410 12613 444
rect 12647 410 12685 444
rect 12719 410 12757 444
rect 12791 410 12829 444
rect 12863 410 12901 444
rect 12935 410 12973 444
rect 13007 410 13045 444
rect 13079 410 13117 444
rect 13151 410 13189 444
rect 13223 410 13250 444
rect 8104 380 8310 384
rect 8112 374 8304 380
rect 8544 376 10392 396
rect 8388 372 10392 376
rect 11078 374 13250 410
rect 5566 290 5618 354
rect 5894 340 6224 356
rect 5894 306 5902 340
rect 5936 306 6224 340
rect 5894 304 6224 306
rect 6276 304 6498 356
rect 8018 304 8072 370
rect 8346 365 10392 372
rect 8346 354 10189 365
rect 8346 320 8354 354
rect 8388 320 10189 354
rect 8346 313 10189 320
rect 10241 313 10392 365
rect 5654 276 5858 292
rect 5894 284 6498 304
rect 8346 300 10392 313
rect 3484 250 3572 262
rect 886 170 1180 186
rect 1222 176 1414 188
rect 886 -46 972 170
rect 1222 142 1266 176
rect 1300 142 1338 176
rect 1372 142 1414 176
rect 886 -144 974 -46
rect 558 -150 974 -144
rect 292 -218 974 -150
rect 1222 -130 1414 142
rect 1812 178 2108 212
rect 2142 178 2158 212
rect 2720 206 3454 226
rect 3484 216 3511 250
rect 3545 216 3572 250
rect 5654 242 5702 276
rect 5736 242 5774 276
rect 5808 242 5858 276
rect 6072 246 6498 284
rect 8106 290 8310 300
rect 8544 290 10392 300
rect 8106 256 8154 290
rect 8188 256 8226 290
rect 8260 256 8310 290
rect 3484 206 3572 216
rect 1812 154 2158 178
rect 2188 168 2392 182
rect 1812 -130 1882 154
rect 1222 -162 1882 -130
rect 2188 134 2236 168
rect 2270 134 2308 168
rect 2342 134 2392 168
rect 2720 172 3414 206
rect 3448 172 3454 206
rect 2720 156 3454 172
rect 3482 162 3572 174
rect 2188 -140 2392 134
rect 3482 128 3511 162
rect 3545 128 3572 162
rect 3600 158 3658 218
rect 3482 64 3572 128
rect 5654 126 5858 242
rect 5652 94 5858 126
rect 3392 48 3660 64
rect 3392 14 3439 48
rect 3473 14 3511 48
rect 3545 14 3583 48
rect 3617 14 3660 48
rect 292 -436 382 -218
rect 294 -448 382 -436
rect 294 -464 319 -448
rect -26 -480 266 -472
rect -26 -532 -3 -480
rect 49 -493 266 -480
rect 296 -482 319 -464
rect 353 -482 382 -448
rect 886 -464 974 -218
rect 1268 -204 1882 -162
rect 296 -490 382 -482
rect 49 -525 222 -493
rect 256 -525 266 -493
rect 410 -493 466 -478
rect 49 -532 266 -525
rect -26 -546 266 -532
rect 296 -536 382 -524
rect 294 -570 319 -536
rect 353 -570 382 -536
rect 410 -525 416 -493
rect 450 -525 466 -493
rect 410 -540 466 -525
rect 886 -534 1238 -464
rect 1268 -480 1400 -204
rect 1812 -466 1882 -204
rect 2250 -202 2384 -140
rect 3392 -160 3660 14
rect 5652 -150 5856 94
rect 5652 -152 6916 -150
rect 3920 -160 4000 -158
rect 3136 -170 4008 -160
rect 2250 -276 2752 -202
rect 3132 -250 4008 -170
rect 2250 -436 2384 -276
rect 294 -580 382 -570
rect 288 -636 382 -580
rect 1268 -632 1402 -516
rect 1432 -532 1486 -470
rect 1812 -480 2220 -466
rect 1812 -514 2178 -480
rect 2212 -514 2220 -480
rect 2250 -470 2262 -436
rect 2296 -470 2334 -436
rect 2368 -440 2384 -436
rect 2368 -470 2382 -440
rect 2652 -456 2750 -276
rect 3132 -430 3218 -250
rect 3920 -422 4008 -250
rect 2652 -464 3096 -456
rect 2250 -482 2382 -470
rect 1812 -528 2220 -514
rect 2250 -514 2380 -510
rect 2250 -524 2382 -514
rect 2250 -558 2262 -524
rect 2296 -558 2334 -524
rect 2368 -558 2382 -524
rect 2414 -528 2464 -466
rect 2652 -516 2676 -464
rect 2728 -516 3096 -464
rect 3132 -472 3216 -430
rect 3442 -450 3518 -422
rect 3442 -454 3886 -450
rect 3138 -476 3216 -472
rect 2652 -524 3096 -516
rect 2652 -526 2750 -524
rect 2250 -626 2382 -558
rect 3126 -614 3216 -506
rect 3244 -520 3300 -458
rect 3442 -506 3455 -454
rect 3507 -506 3886 -454
rect 3920 -456 3945 -422
rect 3979 -456 4008 -422
rect 4698 -170 6916 -152
rect 4698 -222 5197 -170
rect 5249 -174 6916 -170
rect 5249 -222 6313 -174
rect 4698 -226 6313 -222
rect 6365 -226 6916 -174
rect 4698 -398 6916 -226
rect 4698 -414 5700 -398
rect 4698 -448 4713 -414
rect 4747 -448 4785 -414
rect 4819 -448 4857 -414
rect 4891 -448 4929 -414
rect 4963 -448 5001 -414
rect 5035 -448 5073 -414
rect 5107 -448 5145 -414
rect 5179 -448 5217 -414
rect 5251 -448 5289 -414
rect 5323 -448 5361 -414
rect 5395 -448 5433 -414
rect 5467 -448 5505 -414
rect 5539 -448 5577 -414
rect 5611 -448 5649 -414
rect 5683 -448 5700 -414
rect 3920 -466 4008 -456
rect 3924 -502 4004 -498
rect 3442 -516 3886 -506
rect 3920 -510 4004 -502
rect 3920 -544 3945 -510
rect 3979 -544 4004 -510
rect 4036 -514 4092 -452
rect 4698 -458 5700 -448
rect 5914 -414 6916 -398
rect 8106 -372 8310 256
rect 11080 150 13250 374
rect 11020 -108 13422 150
rect 11020 -142 11049 -108
rect 11083 -142 11121 -108
rect 11155 -142 11193 -108
rect 11227 -142 11265 -108
rect 11299 -142 11337 -108
rect 11371 -142 11409 -108
rect 11443 -142 11481 -108
rect 11515 -142 11553 -108
rect 11587 -142 11625 -108
rect 11659 -142 11697 -108
rect 11731 -142 11769 -108
rect 11803 -142 11841 -108
rect 11875 -142 11913 -108
rect 11947 -142 11985 -108
rect 12019 -142 12057 -108
rect 12091 -142 12129 -108
rect 12163 -142 12201 -108
rect 12235 -142 12273 -108
rect 12307 -142 12345 -108
rect 12379 -142 12417 -108
rect 12451 -142 12489 -108
rect 12523 -142 12561 -108
rect 12595 -142 12633 -108
rect 12667 -142 12705 -108
rect 12739 -142 12777 -108
rect 12811 -142 12849 -108
rect 12883 -142 12921 -108
rect 12955 -142 12993 -108
rect 13027 -142 13065 -108
rect 13099 -142 13137 -108
rect 13171 -142 13209 -108
rect 13243 -142 13281 -108
rect 13315 -142 13353 -108
rect 13387 -142 13422 -108
rect 11020 -148 13422 -142
rect 10820 -154 10992 -152
rect 10598 -193 10992 -154
rect 11020 -158 13396 -148
rect 10598 -227 10946 -193
rect 10980 -227 10992 -193
rect 10598 -265 10992 -227
rect 10598 -299 10946 -265
rect 10980 -299 10992 -265
rect 10598 -336 10992 -299
rect 8106 -400 8346 -372
rect 9030 -400 10042 -388
rect 5914 -448 5931 -414
rect 5965 -448 6003 -414
rect 6037 -448 6075 -414
rect 6109 -448 6147 -414
rect 6181 -448 6219 -414
rect 6253 -448 6291 -414
rect 6325 -448 6363 -414
rect 6397 -448 6435 -414
rect 6469 -448 6507 -414
rect 6541 -448 6579 -414
rect 6613 -448 6651 -414
rect 6685 -448 6723 -414
rect 6757 -448 6795 -414
rect 6829 -448 6867 -414
rect 6901 -448 6916 -414
rect 5914 -456 6916 -448
rect 7724 -412 10042 -400
rect 7724 -446 7831 -412
rect 7865 -446 7903 -412
rect 7937 -446 7975 -412
rect 8009 -446 8047 -412
rect 8081 -446 8119 -412
rect 8153 -446 8191 -412
rect 8225 -446 8263 -412
rect 8297 -446 8335 -412
rect 8369 -446 8407 -412
rect 8441 -446 8479 -412
rect 8513 -446 8551 -412
rect 8585 -446 8623 -412
rect 8657 -446 8695 -412
rect 8729 -446 8767 -412
rect 8801 -446 9049 -412
rect 9083 -446 9121 -412
rect 9155 -446 9193 -412
rect 9227 -446 9265 -412
rect 9299 -446 9337 -412
rect 9371 -446 9409 -412
rect 9443 -446 9481 -412
rect 9515 -446 9553 -412
rect 9587 -446 9625 -412
rect 9659 -446 9697 -412
rect 9731 -446 9769 -412
rect 9803 -446 9841 -412
rect 9875 -446 9913 -412
rect 9947 -446 9985 -412
rect 10019 -446 10042 -412
rect 7724 -458 10042 -446
rect 6946 -462 10042 -458
rect 10598 -452 10653 -336
rect 10769 -337 10992 -336
rect 10769 -371 10946 -337
rect 10980 -371 10992 -337
rect 10769 -409 10992 -371
rect 10769 -443 10946 -409
rect 10980 -443 10992 -409
rect 10769 -452 10992 -443
rect 5732 -493 5886 -462
rect 3920 -608 4004 -544
rect 5732 -527 5742 -493
rect 5776 -527 5838 -493
rect 5872 -527 5886 -493
rect 5732 -556 5886 -527
rect 6946 -491 7786 -462
rect 6946 -493 7744 -491
rect 6946 -527 6954 -493
rect 6988 -525 7744 -493
rect 7778 -525 7786 -491
rect 6988 -527 7786 -525
rect 4698 -572 5698 -562
rect 4698 -606 4713 -572
rect 4747 -606 4785 -572
rect 4819 -606 4857 -572
rect 4891 -606 4929 -572
rect 4963 -606 5001 -572
rect 5035 -606 5073 -572
rect 5107 -606 5145 -572
rect 5179 -606 5217 -572
rect 5251 -606 5289 -572
rect 5323 -606 5361 -572
rect 5395 -606 5433 -572
rect 5467 -606 5505 -572
rect 5539 -606 5577 -572
rect 5611 -606 5649 -572
rect 5683 -606 5698 -572
rect 200 -650 466 -636
rect 200 -684 247 -650
rect 281 -684 319 -650
rect 353 -684 391 -650
rect 425 -684 466 -650
rect -743 -840 -150 -838
rect 200 -840 466 -684
rect 1172 -642 1490 -632
rect 1172 -676 1210 -642
rect 1244 -676 1282 -642
rect 1316 -676 1354 -642
rect 1388 -676 1426 -642
rect 1460 -676 1490 -642
rect 1172 -836 1490 -676
rect 2154 -638 2470 -626
rect 2154 -672 2190 -638
rect 2224 -672 2262 -638
rect 2296 -672 2334 -638
rect 2368 -672 2406 -638
rect 2440 -672 2470 -638
rect 2154 -834 2470 -672
rect 3038 -632 3308 -614
rect 3038 -666 3083 -632
rect 3117 -666 3155 -632
rect 3189 -666 3227 -632
rect 3261 -666 3308 -632
rect 1790 -836 2648 -834
rect 3038 -836 3308 -666
rect 3832 -624 4096 -608
rect 3832 -658 3873 -624
rect 3907 -658 3945 -624
rect 3979 -658 4017 -624
rect 4051 -658 4096 -624
rect 3832 -836 4096 -658
rect 4698 -668 5698 -606
rect 5918 -572 6918 -558
rect 6946 -562 7786 -527
rect 8844 -491 9006 -462
rect 8844 -525 8854 -491
rect 8888 -525 8962 -491
rect 8996 -525 9006 -491
rect 8844 -556 9006 -525
rect 10598 -481 10992 -452
rect 10598 -515 10946 -481
rect 10980 -515 10992 -481
rect 10598 -554 10992 -515
rect 11022 -560 13412 -550
rect 5918 -606 5931 -572
rect 5965 -606 6003 -572
rect 6037 -606 6075 -572
rect 6109 -606 6147 -572
rect 6181 -606 6219 -572
rect 6253 -606 6291 -572
rect 6325 -606 6363 -572
rect 6397 -606 6435 -572
rect 6469 -606 6507 -572
rect 6541 -606 6579 -572
rect 6613 -606 6651 -572
rect 6685 -606 6723 -572
rect 6757 -606 6795 -572
rect 6829 -606 6867 -572
rect 6901 -606 6918 -572
rect 4606 -676 5760 -668
rect 5918 -676 6918 -606
rect 7816 -570 8816 -560
rect 7816 -604 7831 -570
rect 7865 -604 7903 -570
rect 7937 -604 7975 -570
rect 8009 -604 8047 -570
rect 8081 -604 8119 -570
rect 8153 -604 8191 -570
rect 8225 -604 8263 -570
rect 8297 -604 8335 -570
rect 8369 -604 8407 -570
rect 8441 -604 8479 -570
rect 8513 -604 8551 -570
rect 8585 -604 8623 -570
rect 8657 -604 8695 -570
rect 8729 -604 8767 -570
rect 8801 -604 8816 -570
rect 7816 -674 8816 -604
rect 9034 -570 10034 -560
rect 9034 -604 9049 -570
rect 9083 -604 9121 -570
rect 9155 -604 9193 -570
rect 9227 -604 9265 -570
rect 9299 -604 9337 -570
rect 9371 -604 9409 -570
rect 9443 -604 9481 -570
rect 9515 -604 9553 -570
rect 9587 -604 9625 -570
rect 9659 -604 9697 -570
rect 9731 -604 9769 -570
rect 9803 -604 9841 -570
rect 9875 -604 9913 -570
rect 9947 -604 9985 -570
rect 10019 -604 10034 -570
rect 9034 -674 10034 -604
rect 11020 -566 13420 -560
rect 11020 -600 11049 -566
rect 11083 -600 11121 -566
rect 11155 -600 11193 -566
rect 11227 -600 11265 -566
rect 11299 -600 11337 -566
rect 11371 -600 11409 -566
rect 11443 -600 11481 -566
rect 11515 -600 11553 -566
rect 11587 -600 11625 -566
rect 11659 -600 11697 -566
rect 11731 -600 11769 -566
rect 11803 -600 11841 -566
rect 11875 -600 11913 -566
rect 11947 -600 11985 -566
rect 12019 -600 12057 -566
rect 12091 -600 12129 -566
rect 12163 -600 12201 -566
rect 12235 -600 12273 -566
rect 12307 -600 12345 -566
rect 12379 -600 12417 -566
rect 12451 -600 12489 -566
rect 12523 -600 12561 -566
rect 12595 -600 12633 -566
rect 12667 -600 12705 -566
rect 12739 -600 12777 -566
rect 12811 -600 12849 -566
rect 12883 -600 12921 -566
rect 12955 -600 12993 -566
rect 13027 -600 13065 -566
rect 13099 -600 13137 -566
rect 13171 -600 13209 -566
rect 13243 -600 13281 -566
rect 13315 -600 13353 -566
rect 13387 -600 13420 -566
rect 11020 -660 13420 -600
rect 7726 -676 10118 -674
rect 4606 -686 7010 -676
rect 4606 -720 4638 -686
rect 4672 -720 4710 -686
rect 4744 -720 4782 -686
rect 4816 -720 4854 -686
rect 4888 -720 4926 -686
rect 4960 -720 4998 -686
rect 5032 -720 5070 -686
rect 5104 -720 5142 -686
rect 5176 -720 5214 -686
rect 5248 -720 5286 -686
rect 5320 -720 5358 -686
rect 5392 -720 5430 -686
rect 5464 -720 5502 -686
rect 5536 -720 5574 -686
rect 5608 -720 5646 -686
rect 5680 -720 5718 -686
rect 5752 -720 5790 -686
rect 5824 -720 5862 -686
rect 5896 -720 5934 -686
rect 5968 -720 6006 -686
rect 6040 -720 6078 -686
rect 6112 -720 6150 -686
rect 6184 -720 6222 -686
rect 6256 -720 6294 -686
rect 6328 -720 6366 -686
rect 6400 -720 6438 -686
rect 6472 -720 6510 -686
rect 6544 -720 6582 -686
rect 6616 -720 6654 -686
rect 6688 -720 6726 -686
rect 6760 -720 6798 -686
rect 6832 -720 6870 -686
rect 6904 -720 6942 -686
rect 6976 -720 7010 -686
rect 4606 -834 7010 -720
rect 7726 -684 10126 -676
rect 7726 -718 7756 -684
rect 7790 -718 7828 -684
rect 7862 -718 7900 -684
rect 7934 -718 7972 -684
rect 8006 -718 8044 -684
rect 8078 -718 8116 -684
rect 8150 -718 8188 -684
rect 8222 -718 8260 -684
rect 8294 -718 8332 -684
rect 8366 -718 8404 -684
rect 8438 -718 8476 -684
rect 8510 -718 8548 -684
rect 8582 -718 8620 -684
rect 8654 -718 8692 -684
rect 8726 -718 8764 -684
rect 8798 -718 8836 -684
rect 8870 -718 8908 -684
rect 8942 -718 8980 -684
rect 9014 -718 9052 -684
rect 9086 -718 9124 -684
rect 9158 -718 9196 -684
rect 9230 -718 9268 -684
rect 9302 -718 9340 -684
rect 9374 -718 9412 -684
rect 9446 -718 9484 -684
rect 9518 -718 9556 -684
rect 9590 -718 9628 -684
rect 9662 -718 9700 -684
rect 9734 -718 9772 -684
rect 9806 -718 9844 -684
rect 9878 -718 9916 -684
rect 9950 -718 9988 -684
rect 10022 -718 10060 -684
rect 10094 -718 10126 -684
rect 7726 -832 10126 -718
rect 10934 -680 13510 -660
rect 10934 -714 10941 -680
rect 10975 -714 11013 -680
rect 11047 -714 11085 -680
rect 11119 -714 11157 -680
rect 11191 -714 11229 -680
rect 11263 -714 11301 -680
rect 11335 -714 11373 -680
rect 11407 -714 11445 -680
rect 11479 -714 11517 -680
rect 11551 -714 11589 -680
rect 11623 -714 11661 -680
rect 11695 -714 11733 -680
rect 11767 -714 11805 -680
rect 11839 -714 11877 -680
rect 11911 -714 11949 -680
rect 11983 -714 12021 -680
rect 12055 -714 12093 -680
rect 12127 -714 12165 -680
rect 12199 -714 12237 -680
rect 12271 -714 12309 -680
rect 12343 -714 12381 -680
rect 12415 -714 12453 -680
rect 12487 -714 12525 -680
rect 12559 -714 12597 -680
rect 12631 -714 12669 -680
rect 12703 -714 12741 -680
rect 12775 -714 12813 -680
rect 12847 -714 12885 -680
rect 12919 -714 12957 -680
rect 12991 -714 13029 -680
rect 13063 -714 13101 -680
rect 13135 -714 13173 -680
rect 13207 -714 13245 -680
rect 13279 -714 13317 -680
rect 13351 -714 13389 -680
rect 13423 -714 13461 -680
rect 13495 -714 13510 -680
rect 10934 -824 13510 -714
rect 10626 -832 13652 -824
rect 7726 -834 13652 -832
rect 4606 -836 13652 -834
rect 766 -840 13652 -836
rect -743 -871 13652 -840
rect -743 -877 11599 -871
rect -743 -883 4647 -877
rect -743 -884 4393 -883
rect -743 -886 2702 -884
rect -743 -888 185 -886
rect -743 -922 -123 -888
rect -89 -922 27 -888
rect 61 -920 185 -888
rect 219 -887 2702 -886
rect 219 -888 716 -887
rect 219 -920 333 -888
rect 61 -922 333 -920
rect 367 -922 483 -888
rect 517 -922 629 -888
rect 663 -921 716 -888
rect 750 -891 984 -887
rect 750 -921 846 -891
rect 663 -922 846 -921
rect -743 -925 846 -922
rect 880 -921 984 -891
rect 1018 -889 1556 -887
rect 1018 -921 1126 -889
rect 880 -923 1126 -921
rect 1160 -893 1414 -889
rect 1160 -923 1268 -893
rect 880 -925 1268 -923
rect -743 -927 1268 -925
rect 1302 -923 1414 -893
rect 1448 -921 1556 -889
rect 1590 -921 1728 -887
rect 1762 -889 2702 -887
rect 1762 -891 2050 -889
rect 1762 -921 1896 -891
rect 1448 -923 1896 -921
rect 1302 -925 1896 -923
rect 1930 -923 2050 -891
rect 2084 -923 2198 -889
rect 2232 -923 2340 -889
rect 2374 -923 2510 -889
rect 2544 -918 2702 -889
rect 2736 -918 2870 -884
rect 2904 -918 3042 -884
rect 3076 -918 3220 -884
rect 3254 -886 4072 -884
rect 3254 -918 3392 -886
rect 2544 -920 3392 -918
rect 3426 -890 3742 -886
rect 3426 -920 3558 -890
rect 2544 -923 3558 -920
rect 1930 -924 3558 -923
rect 3592 -920 3742 -890
rect 3776 -920 3912 -886
rect 3946 -918 4072 -886
rect 4106 -918 4252 -884
rect 4286 -917 4393 -884
rect 4427 -917 4517 -883
rect 4551 -911 4647 -883
rect 4681 -911 4785 -877
rect 4819 -911 4921 -877
rect 4955 -911 5063 -877
rect 5097 -883 5551 -877
rect 5097 -911 5221 -883
rect 4551 -917 5221 -911
rect 5255 -917 5389 -883
rect 5423 -911 5551 -883
rect 5585 -879 6001 -877
rect 5585 -883 5845 -879
rect 5585 -911 5691 -883
rect 5423 -917 5691 -911
rect 5725 -913 5845 -883
rect 5879 -911 6001 -879
rect 6035 -879 10803 -877
rect 6035 -883 6293 -879
rect 6035 -911 6151 -883
rect 5879 -913 6151 -911
rect 5725 -917 6151 -913
rect 6185 -913 6293 -883
rect 6327 -913 6441 -879
rect 6475 -881 10803 -879
rect 6475 -883 10619 -881
rect 6475 -913 6585 -883
rect 6185 -917 6585 -913
rect 6619 -917 6719 -883
rect 6753 -885 7541 -883
rect 6753 -889 7239 -885
rect 6753 -917 6849 -889
rect 4286 -918 6849 -917
rect 3946 -920 6849 -918
rect 3592 -923 6849 -920
rect 6883 -923 6967 -889
rect 7001 -923 7101 -889
rect 7135 -919 7239 -889
rect 7273 -919 7385 -885
rect 7419 -917 7541 -885
rect 7575 -917 7711 -883
rect 7745 -887 8007 -883
rect 7745 -917 7869 -887
rect 7419 -919 7869 -917
rect 7135 -921 7869 -919
rect 7903 -917 8007 -887
rect 8041 -885 9273 -883
rect 8041 -917 8151 -885
rect 7903 -919 8151 -917
rect 8185 -887 9273 -885
rect 8185 -919 8307 -887
rect 7903 -921 8307 -919
rect 8341 -921 8443 -887
rect 8477 -921 8585 -887
rect 8619 -893 8937 -887
rect 8619 -921 8733 -893
rect 7135 -923 8733 -921
rect 3592 -924 8733 -923
rect 1930 -925 8733 -924
rect 1302 -927 8733 -925
rect 8767 -921 8937 -893
rect 8971 -893 9273 -887
rect 8971 -921 9109 -893
rect 8767 -927 9109 -921
rect 9143 -917 9273 -893
rect 9307 -917 9471 -883
rect 9505 -885 9943 -883
rect 9505 -887 9777 -885
rect 9505 -917 9639 -887
rect 9143 -921 9639 -917
rect 9673 -919 9777 -887
rect 9811 -917 9943 -885
rect 9977 -885 10619 -883
rect 9977 -917 10137 -885
rect 9811 -919 10137 -917
rect 10171 -887 10619 -885
rect 10171 -889 10467 -887
rect 10171 -919 10299 -889
rect 9673 -921 10299 -919
rect 9143 -923 10299 -921
rect 10333 -921 10467 -889
rect 10501 -915 10619 -887
rect 10653 -911 10803 -881
rect 10837 -911 11013 -877
rect 11047 -911 11209 -877
rect 11243 -911 11399 -877
rect 11433 -905 11599 -877
rect 11633 -877 13652 -871
rect 11633 -881 11959 -877
rect 11633 -905 11783 -881
rect 11433 -911 11783 -905
rect 10653 -915 11783 -911
rect 11817 -911 11959 -881
rect 11993 -881 12963 -877
rect 11993 -887 12343 -881
rect 11993 -911 12129 -887
rect 11817 -915 12129 -911
rect 10501 -921 12129 -915
rect 12163 -915 12343 -887
rect 12377 -915 12539 -881
rect 12573 -891 12963 -881
rect 12573 -915 12723 -891
rect 12163 -921 12723 -915
rect 10333 -923 12723 -921
rect 9143 -925 12723 -923
rect 12757 -911 12963 -891
rect 12997 -881 13445 -877
rect 12997 -911 13187 -881
rect 12757 -915 13187 -911
rect 13221 -911 13445 -881
rect 13479 -911 13652 -877
rect 13221 -915 13652 -911
rect 12757 -925 13652 -915
rect 9143 -927 13652 -925
rect -743 -974 13652 -927
rect -743 -1046 -150 -974
rect 2598 -976 13652 -974
rect 2598 -978 9278 -976
rect 2598 -980 6084 -978
rect 10626 -984 13652 -976
rect -743 -1226 -600 -1046
rect -420 -1226 -150 -1046
rect -743 -1378 -150 -1226
rect 2475 -1249 2941 -1115
rect 2475 -1429 2618 -1249
rect 2798 -1429 2941 -1249
rect 2475 -1581 2941 -1429
<< via1 >>
rect 2661 2728 2841 2908
rect -597 1535 -417 1715
rect -597 520 -417 700
rect -597 -380 -417 -200
rect 9289 1815 9341 1867
rect 9289 1751 9341 1803
rect 10128 1018 10244 1134
rect 6224 304 6276 356
rect 10189 313 10241 365
rect -3 -532 49 -480
rect 2676 -516 2728 -464
rect 3455 -506 3507 -454
rect 5197 -222 5249 -170
rect 6313 -226 6365 -174
rect 10653 -452 10769 -336
rect -600 -1226 -420 -1046
rect 2618 -1429 2798 -1249
<< metal2 >>
rect 2518 2925 2984 3042
rect 2518 2709 2643 2925
rect 2859 2709 2984 2925
rect 2518 2576 2984 2709
rect -740 1867 9400 2038
rect -740 1815 9289 1867
rect 9341 1815 9400 1867
rect -740 1803 9400 1815
rect -740 1751 9289 1803
rect 9341 1751 9400 1803
rect -740 1732 9400 1751
rect -740 1516 -615 1732
rect -399 1632 9400 1732
rect -399 1516 -274 1632
rect -740 1383 -274 1516
rect -740 717 -274 834
rect -740 501 -615 717
rect -399 501 -274 717
rect -740 368 -274 501
rect 6368 430 6656 1632
rect 10076 1134 10330 1190
rect 10076 1018 10128 1134
rect 10244 1018 10330 1134
rect 10076 978 10330 1018
rect 10076 842 10332 978
rect 6072 356 6656 430
rect 6072 304 6224 356
rect 6276 304 6656 356
rect 6072 246 6656 304
rect 10084 365 10332 842
rect 10084 313 10189 365
rect 10241 313 10332 365
rect 10084 250 10332 313
rect 6368 242 6656 246
rect -740 -154 72 -66
rect 2060 -154 3522 -152
rect 6890 -154 10750 -152
rect -740 -170 10790 -154
rect -740 -183 5197 -170
rect -740 -399 -615 -183
rect -399 -222 5197 -183
rect 5249 -174 10790 -170
rect 5249 -222 6313 -174
rect -399 -226 6313 -222
rect 6365 -226 10790 -174
rect -399 -242 10790 -226
rect -399 -244 3522 -242
rect -399 -399 72 -244
rect -740 -480 72 -399
rect -740 -532 -3 -480
rect 49 -532 72 -480
rect -740 -542 72 -532
rect 2643 -464 2763 -449
rect 2643 -516 2676 -464
rect 2728 -516 2763 -464
rect -743 -1029 -277 -912
rect -743 -1245 -618 -1029
rect -402 -1245 -277 -1029
rect 2643 -1115 2763 -516
rect 3436 -454 3522 -244
rect 6890 -244 10790 -242
rect 6890 -246 10110 -244
rect 3436 -506 3455 -454
rect 3507 -506 3522 -454
rect 10636 -336 10790 -244
rect 10636 -452 10653 -336
rect 10769 -452 10790 -336
rect 10636 -476 10790 -452
rect 3436 -518 3522 -506
rect -743 -1378 -277 -1245
rect 2475 -1232 2941 -1115
rect 2475 -1448 2600 -1232
rect 2816 -1448 2941 -1232
rect 2475 -1581 2941 -1448
<< via2 >>
rect 2643 2908 2859 2925
rect 2643 2728 2661 2908
rect 2661 2728 2841 2908
rect 2841 2728 2859 2908
rect 2643 2709 2859 2728
rect -615 1715 -399 1732
rect -615 1535 -597 1715
rect -597 1535 -417 1715
rect -417 1535 -399 1715
rect -615 1516 -399 1535
rect -615 700 -399 717
rect -615 520 -597 700
rect -597 520 -417 700
rect -417 520 -399 700
rect -615 501 -399 520
rect -615 -200 -399 -183
rect -615 -380 -597 -200
rect -597 -380 -417 -200
rect -417 -380 -399 -200
rect -615 -399 -399 -380
rect -618 -1046 -402 -1029
rect -618 -1226 -600 -1046
rect -600 -1226 -420 -1046
rect -420 -1226 -402 -1046
rect -618 -1245 -402 -1226
rect 2600 -1249 2816 -1232
rect 2600 -1429 2618 -1249
rect 2618 -1429 2798 -1249
rect 2798 -1429 2816 -1249
rect 2600 -1448 2816 -1429
<< metal3 >>
rect 2518 2964 2984 3042
rect 2518 2660 2598 2964
rect 2902 2660 2984 2964
rect 2518 2576 2984 2660
rect -740 1771 -274 1849
rect -740 1467 -660 1771
rect -356 1467 -274 1771
rect -740 1383 -274 1467
rect -740 756 -274 834
rect -740 452 -660 756
rect -356 452 -274 756
rect -740 368 -274 452
rect -740 -144 -274 -66
rect -740 -448 -660 -144
rect -356 -448 -274 -144
rect -740 -532 -274 -448
rect -743 -990 -277 -912
rect -743 -1294 -663 -990
rect -359 -1294 -277 -990
rect -743 -1378 -277 -1294
rect 2475 -1193 2941 -1115
rect 2475 -1497 2555 -1193
rect 2859 -1497 2941 -1193
rect 2475 -1581 2941 -1497
<< via3 >>
rect 2598 2925 2902 2964
rect 2598 2709 2643 2925
rect 2643 2709 2859 2925
rect 2859 2709 2902 2925
rect 2598 2660 2902 2709
rect -660 1732 -356 1771
rect -660 1516 -615 1732
rect -615 1516 -399 1732
rect -399 1516 -356 1732
rect -660 1467 -356 1516
rect -660 717 -356 756
rect -660 501 -615 717
rect -615 501 -399 717
rect -399 501 -356 717
rect -660 452 -356 501
rect -660 -183 -356 -144
rect -660 -399 -615 -183
rect -615 -399 -399 -183
rect -399 -399 -356 -183
rect -660 -448 -356 -399
rect -663 -1029 -359 -990
rect -663 -1245 -618 -1029
rect -618 -1245 -402 -1029
rect -402 -1245 -359 -1029
rect -663 -1294 -359 -1245
rect 2555 -1232 2859 -1193
rect 2555 -1448 2600 -1232
rect 2600 -1448 2816 -1232
rect 2816 -1448 2859 -1232
rect 2555 -1497 2859 -1448
<< metal4 >>
rect 2518 2964 2984 3042
rect 2518 2660 2598 2964
rect 2902 2660 2984 2964
rect 2518 2576 2984 2660
rect -740 1771 -274 1849
rect -740 1467 -660 1771
rect -356 1467 -274 1771
rect -740 1383 -274 1467
rect -740 756 -274 834
rect -740 452 -660 756
rect -356 452 -274 756
rect -740 368 -274 452
rect -740 -144 -274 -66
rect -740 -448 -660 -144
rect -356 -448 -274 -144
rect -740 -532 -274 -448
rect -743 -990 -277 -912
rect -743 -1294 -663 -990
rect -359 -1294 -277 -990
rect -743 -1378 -277 -1294
rect 2475 -1193 2941 -1115
rect 2475 -1497 2555 -1193
rect 2859 -1497 2941 -1193
rect 2475 -1581 2941 -1497
<< via4 >>
rect 2632 2694 2868 2930
rect -626 1501 -390 1737
rect -626 486 -390 722
rect -626 -414 -390 -178
rect -629 -1260 -393 -1024
rect 2589 -1463 2825 -1227
<< metal5 >>
rect 2518 2930 2984 3042
rect 2518 2694 2632 2930
rect 2868 2694 2984 2930
rect 2518 2576 2984 2694
rect -740 1737 -274 1849
rect -740 1501 -626 1737
rect -390 1501 -274 1737
rect -740 1383 -274 1501
rect -740 722 -274 834
rect -740 486 -626 722
rect -390 486 -274 722
rect -740 368 -274 486
rect -740 -178 -274 -66
rect -740 -414 -626 -178
rect -390 -414 -274 -178
rect -740 -532 -274 -414
rect -743 -1024 -277 -912
rect -743 -1260 -629 -1024
rect -393 -1260 -277 -1024
rect -743 -1378 -277 -1260
rect 2475 -1227 2941 -1115
rect 2475 -1463 2589 -1227
rect 2825 -1463 2941 -1227
rect 2475 -1581 2941 -1463
use sky130_fd_pr__nfet_01v8_lvt_XXD9Y4  sky130_fd_pr__nfet_01v8_lvt_XXD9Y4_0
timestamp 1611881054
transform 0 1 336 -1 0 -509
box -175 -216 175 216
use sky130_fd_pr__nfet_01v8_5K7Q63  sky130_fd_pr__nfet_01v8_5K7Q63_1
timestamp 1611881054
transform 0 1 1336 -1 0 -501
box -175 -238 175 238
use sky130_fd_pr__nfet_01v8_5K7Q63  sky130_fd_pr__nfet_01v8_5K7Q63_0
timestamp 1611881054
transform 0 1 2314 -1 0 -497
box -175 -238 175 238
use sky130_fd_pr__pfet_01v8_BFRLXZ  sky130_fd_pr__pfet_01v8_BFRLXZ_1
timestamp 1611881054
transform 0 1 1319 -1 0 203
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_BFRLXZ  sky130_fd_pr__pfet_01v8_BFRLXZ_0
timestamp 1611881054
transform 0 1 2289 -1 0 195
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_XAABVK  sky130_fd_pr__nfet_01v8_XAABVK_1
timestamp 1611881054
transform 0 1 5807 -1 0 -510
box -210 -1283 210 1283
use sky130_fd_pr__pfet_01v8_lvt_YTP334  sky130_fd_pr__pfet_01v8_lvt_YTP334_1
timestamp 1611881054
transform 0 1 5755 -1 0 323
box -231 -319 231 319
use sky130_fd_pr__nfet_01v8_6MNZ3F  sky130_fd_pr__nfet_01v8_6MNZ3F_2
timestamp 1611881054
transform 0 1 3962 -1 0 -483
box -175 -216 175 216
use sky130_fd_pr__nfet_01v8_6MNZ3F  sky130_fd_pr__nfet_01v8_6MNZ3F_1
timestamp 1611881054
transform 0 1 3528 -1 0 189
box -175 -216 175 216
use sky130_fd_pr__nfet_01v8_6MNZ3F  sky130_fd_pr__nfet_01v8_6MNZ3F_0
timestamp 1611881054
transform 0 1 3172 -1 0 -489
box -175 -216 175 216
use sky130_fd_pr__pfet_01v8_lvt_EWYCPT  sky130_fd_pr__pfet_01v8_lvt_EWYCPT_1
timestamp 1611881054
transform 0 1 3839 -1 0 1241
box -696 -969 696 969
use sky130_fd_pr__nfet_01v8_XAABVK  sky130_fd_pr__nfet_01v8_XAABVK_0
timestamp 1611881054
transform 0 1 8925 -1 0 -508
box -210 -1283 210 1283
use sky130_fd_pr__pfet_01v8_lvt_YTP334  sky130_fd_pr__pfet_01v8_lvt_YTP334_0
timestamp 1611881054
transform 0 1 8207 -1 0 337
box -231 -319 231 319
use sky130_fd_pr__nfet_01v8_lvt_VCXMU2  sky130_fd_pr__nfet_01v8_lvt_VCXMU2_0
timestamp 1611881054
transform 0 1 12218 -1 0 -354
box -360 -1374 360 1374
use sky130_fd_pr__nfet_01v8_3BUYA5  sky130_fd_pr__nfet_01v8_3BUYA5_0
timestamp 1611881054
transform 0 1 12162 -1 0 585
box -175 -1174 175 1174
use sky130_fd_pr__pfet_01v8_lvt_EWYCPT  sky130_fd_pr__pfet_01v8_lvt_EWYCPT_0
timestamp 1611881054
transform 0 1 6941 -1 0 1523
box -696 -969 696 969
use sky130_fd_pr__pfet_01v8_lvt_4N9J2Y  sky130_fd_pr__pfet_01v8_lvt_4N9J2Y_1
timestamp 1611881054
transform 0 1 10465 -1 0 1847
box -396 -1219 396 1219
use sky130_fd_pr__pfet_01v8_lvt_4N9J2Y  sky130_fd_pr__pfet_01v8_lvt_4N9J2Y_0
timestamp 1611881054
transform 0 1 13063 -1 0 1845
box -396 -1219 396 1219
<< labels >>
rlabel metal2 s 0 -530 48 -486 4 vbn
port 1 nsew
rlabel metal1 s 302 -224 366 -156 4 Inv1IN
port 2 nsew
rlabel metal1 s 304 -932 368 -864 4 Gnd
port 3 nsew
rlabel metal1 s 1284 -204 1372 -146 4 Inv2IN
port 4 nsew
rlabel metal1 s 2272 -214 2370 -116 4 Vinit
port 5 nsew
rlabel metal1 s 3504 -124 3562 -60 4 AmpBias2
port 6 nsew
rlabel metal1 s 6084 296 6130 348 4 Vcntrl
port 7 nsew
rlabel metal1 s 8576 304 8634 364 4 DiifAmpPos
port 8 nsew
<< end >>
