magic
tech sky130A
magscale 1 2
timestamp 1607669338
<< error_p >>
rect 19 126 77 132
rect 19 92 31 126
rect 19 86 77 92
rect -77 -92 -19 -86
rect -77 -126 -65 -92
rect -77 -132 -19 -126
<< pwell >>
rect -263 -264 263 264
<< nmos >>
rect -63 -54 -33 54
rect 33 -54 63 54
<< ndiff >>
rect -125 42 -63 54
rect -125 -42 -113 42
rect -79 -42 -63 42
rect -125 -54 -63 -42
rect -33 42 33 54
rect -33 -42 -17 42
rect 17 -42 33 42
rect -33 -54 33 -42
rect 63 42 125 54
rect 63 -42 79 42
rect 113 -42 125 42
rect 63 -54 125 -42
<< ndiffc >>
rect -113 -42 -79 42
rect -17 -42 17 42
rect 79 -42 113 42
<< psubdiff >>
rect -227 194 -131 228
rect 131 194 227 228
rect -227 132 -193 194
rect 193 132 227 194
rect -227 -194 -193 -132
rect 193 -194 227 -132
rect -227 -228 -131 -194
rect 131 -228 227 -194
<< psubdiffcont >>
rect -131 194 131 228
rect -227 -132 -193 132
rect 193 -132 227 132
rect -131 -228 131 -194
<< poly >>
rect 15 126 81 142
rect 15 92 31 126
rect 65 92 81 126
rect -63 54 -33 80
rect 15 76 81 92
rect 33 54 63 76
rect -63 -76 -33 -54
rect -81 -92 -15 -76
rect 33 -80 63 -54
rect -81 -126 -65 -92
rect -31 -126 -15 -92
rect -81 -142 -15 -126
<< polycont >>
rect 31 92 65 126
rect -65 -126 -31 -92
<< locali >>
rect -227 194 -131 228
rect 131 194 227 228
rect -227 132 -193 194
rect 193 132 227 194
rect 15 92 31 126
rect 65 92 81 126
rect -113 42 -79 58
rect -113 -58 -79 -42
rect -17 42 17 58
rect -17 -58 17 -42
rect 79 42 113 58
rect 79 -58 113 -42
rect -81 -126 -65 -92
rect -31 -126 -15 -92
rect -227 -194 -193 -132
rect 193 -194 227 -132
rect -227 -228 -131 -194
rect 131 -228 227 -194
<< viali >>
rect 31 92 65 126
rect -113 -42 -79 42
rect -17 -42 17 42
rect 79 -42 113 42
rect -65 -126 -31 -92
<< metal1 >>
rect 19 126 77 132
rect 19 92 31 126
rect 65 92 77 126
rect 19 86 77 92
rect -119 42 -73 54
rect -119 -42 -113 42
rect -79 -42 -73 42
rect -119 -54 -73 -42
rect -23 42 23 54
rect -23 -42 -17 42
rect 17 -42 23 42
rect -23 -54 23 -42
rect 73 42 119 54
rect 73 -42 79 42
rect 113 -42 119 42
rect 73 -54 119 -42
rect -77 -92 -19 -86
rect -77 -126 -65 -92
rect -31 -126 -19 -92
rect -77 -132 -19 -126
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -210 -211 210 211
string parameters w 0.54 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
