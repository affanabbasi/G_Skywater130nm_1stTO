magic
tech sky130A
magscale 1 2
timestamp 1608071797
<< error_p >>
rect -1558 746 -1190 747
rect -1100 746 -732 747
rect -642 746 -274 747
rect -184 746 184 747
rect 274 746 642 747
rect 732 746 1100 747
rect 1190 746 1558 747
rect -1574 -700 -1174 -699
rect -1116 -700 -716 -699
rect -658 -700 -258 -699
rect -200 -700 200 -699
rect 258 -700 658 -699
rect 716 -700 1116 -699
rect 1174 -700 1574 -699
<< nwell >>
rect -1770 -918 1770 918
<< pmos >>
rect -1574 -700 -1174 700
rect -1116 -700 -716 700
rect -658 -700 -258 700
rect -200 -700 200 700
rect 258 -700 658 700
rect 716 -700 1116 700
rect 1174 -700 1574 700
<< pdiff >>
rect -1632 688 -1574 700
rect -1632 -688 -1620 688
rect -1586 -688 -1574 688
rect -1632 -700 -1574 -688
rect -1174 688 -1116 700
rect -1174 -688 -1162 688
rect -1128 -688 -1116 688
rect -1174 -700 -1116 -688
rect -716 688 -658 700
rect -716 -688 -704 688
rect -670 -688 -658 688
rect -716 -700 -658 -688
rect -258 688 -200 700
rect -258 -688 -246 688
rect -212 -688 -200 688
rect -258 -700 -200 -688
rect 200 688 258 700
rect 200 -688 212 688
rect 246 -688 258 688
rect 200 -700 258 -688
rect 658 688 716 700
rect 658 -688 670 688
rect 704 -688 716 688
rect 658 -700 716 -688
rect 1116 688 1174 700
rect 1116 -688 1128 688
rect 1162 -688 1174 688
rect 1116 -700 1174 -688
rect 1574 688 1632 700
rect 1574 -688 1586 688
rect 1620 -688 1632 688
rect 1574 -700 1632 -688
<< pdiffc >>
rect -1620 -688 -1586 688
rect -1162 -688 -1128 688
rect -704 -688 -670 688
rect -246 -688 -212 688
rect 212 -688 246 688
rect 670 -688 704 688
rect 1128 -688 1162 688
rect 1586 -688 1620 688
<< nsubdiff >>
rect -1734 848 -1638 882
rect 1638 848 1734 882
rect -1734 786 -1700 848
rect 1700 786 1734 848
rect -1734 -848 -1700 -786
rect 1700 -848 1734 -786
rect -1734 -882 -1638 -848
rect 1638 -882 1734 -848
<< nsubdiffcont >>
rect -1638 848 1638 882
rect -1734 -786 -1700 786
rect 1700 -786 1734 786
rect -1638 -882 1638 -848
<< poly >>
rect -1574 780 -1174 796
rect -1574 746 -1558 780
rect -1190 746 -1174 780
rect -1574 700 -1174 746
rect -1116 780 -716 796
rect -1116 746 -1100 780
rect -732 746 -716 780
rect -1116 700 -716 746
rect -658 780 -258 796
rect -658 746 -642 780
rect -274 746 -258 780
rect -658 700 -258 746
rect -200 780 200 796
rect -200 746 -184 780
rect 184 746 200 780
rect -200 700 200 746
rect 258 780 658 796
rect 258 746 274 780
rect 642 746 658 780
rect 258 700 658 746
rect 716 780 1116 796
rect 716 746 732 780
rect 1100 746 1116 780
rect 716 700 1116 746
rect 1174 780 1574 796
rect 1174 746 1190 780
rect 1558 746 1574 780
rect 1174 700 1574 746
rect -1574 -746 -1174 -700
rect -1574 -780 -1558 -746
rect -1190 -780 -1174 -746
rect -1574 -796 -1174 -780
rect -1116 -746 -716 -700
rect -1116 -780 -1100 -746
rect -732 -780 -716 -746
rect -1116 -796 -716 -780
rect -658 -746 -258 -700
rect -658 -780 -642 -746
rect -274 -780 -258 -746
rect -658 -796 -258 -780
rect -200 -746 200 -700
rect -200 -780 -184 -746
rect 184 -780 200 -746
rect -200 -796 200 -780
rect 258 -746 658 -700
rect 258 -780 274 -746
rect 642 -780 658 -746
rect 258 -796 658 -780
rect 716 -746 1116 -700
rect 716 -780 732 -746
rect 1100 -780 1116 -746
rect 716 -796 1116 -780
rect 1174 -746 1574 -700
rect 1174 -780 1190 -746
rect 1558 -780 1574 -746
rect 1174 -796 1574 -780
<< polycont >>
rect -1558 746 -1190 780
rect -1100 746 -732 780
rect -642 746 -274 780
rect -184 746 184 780
rect 274 746 642 780
rect 732 746 1100 780
rect 1190 746 1558 780
rect -1558 -780 -1190 -746
rect -1100 -780 -732 -746
rect -642 -780 -274 -746
rect -184 -780 184 -746
rect 274 -780 642 -746
rect 732 -780 1100 -746
rect 1190 -780 1558 -746
<< locali >>
rect -1734 848 -1638 882
rect 1638 848 1734 882
rect -1734 786 -1700 848
rect 1700 786 1734 848
rect -1574 746 -1558 780
rect -1190 746 -1174 780
rect -1116 746 -1100 780
rect -732 746 -716 780
rect -658 746 -642 780
rect -274 746 -258 780
rect -200 746 -184 780
rect 184 746 200 780
rect 258 746 274 780
rect 642 746 658 780
rect 716 746 732 780
rect 1100 746 1116 780
rect 1174 746 1190 780
rect 1558 746 1574 780
rect -1620 688 -1586 704
rect -1620 -704 -1586 -688
rect -1162 688 -1128 704
rect -1162 -704 -1128 -688
rect -704 688 -670 704
rect -704 -704 -670 -688
rect -246 688 -212 704
rect -246 -704 -212 -688
rect 212 688 246 704
rect 212 -704 246 -688
rect 670 688 704 704
rect 670 -704 704 -688
rect 1128 688 1162 704
rect 1128 -704 1162 -688
rect 1586 688 1620 704
rect 1586 -704 1620 -688
rect -1574 -780 -1558 -746
rect -1190 -780 -1174 -746
rect -1116 -780 -1100 -746
rect -732 -780 -716 -746
rect -658 -780 -642 -746
rect -274 -780 -258 -746
rect -200 -780 -184 -746
rect 184 -780 200 -746
rect 258 -780 274 -746
rect 642 -780 658 -746
rect 716 -780 732 -746
rect 1100 -780 1116 -746
rect 1174 -780 1190 -746
rect 1558 -780 1574 -746
rect -1734 -848 -1700 -786
rect 1700 -848 1734 -786
rect -1734 -882 -1638 -848
rect 1638 -882 1734 -848
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1716 -866 1716 866
string parameters w 7 l 2 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
