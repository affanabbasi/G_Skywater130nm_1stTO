magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< error_p >>
rect -29 136 29 142
rect -29 102 -17 136
rect -29 96 29 102
rect -29 -102 29 -96
rect -29 -136 -17 -102
rect -29 -142 29 -136
<< pwell >>
rect -175 204 175 238
rect -175 -204 -141 204
rect 141 -204 175 204
rect -175 -238 175 -204
<< nmos >>
rect -15 -64 15 64
<< ndiff >>
rect -73 51 -15 64
rect -73 17 -61 51
rect -27 17 -15 51
rect -73 -17 -15 17
rect -73 -51 -61 -17
rect -27 -51 -15 -17
rect -73 -64 -15 -51
rect 15 51 73 64
rect 15 17 27 51
rect 61 17 73 51
rect 15 -17 73 17
rect 15 -51 27 -17
rect 61 -51 73 -17
rect 15 -64 73 -51
<< ndiffc >>
rect -61 17 -27 51
rect -61 -51 -27 -17
rect 27 17 61 51
rect 27 -51 61 -17
<< psubdiff >>
rect -175 204 -51 238
rect -17 204 17 238
rect 51 204 175 238
rect -175 119 -141 204
rect 141 119 175 204
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -204 -141 -119
rect 141 -204 175 -119
rect -175 -238 -51 -204
rect -17 -238 17 -204
rect 51 -238 175 -204
<< psubdiffcont >>
rect -51 204 -17 238
rect 17 204 51 238
rect -175 85 -141 119
rect 141 85 175 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect 141 17 175 51
rect 141 -51 175 -17
rect -175 -119 -141 -85
rect 141 -119 175 -85
rect -51 -238 -17 -204
rect 17 -238 51 -204
<< poly >>
rect -33 136 33 152
rect -33 102 -17 136
rect 17 102 33 136
rect -33 86 33 102
rect -15 64 15 86
rect -15 -86 15 -64
rect -33 -102 33 -86
rect -33 -136 -17 -102
rect 17 -136 33 -102
rect -33 -152 33 -136
<< polycont >>
rect -17 102 17 136
rect -17 -136 17 -102
<< locali >>
rect -175 204 -51 238
rect -17 204 17 238
rect 51 204 175 238
rect -175 119 -141 204
rect -33 102 -17 136
rect 17 102 33 136
rect 141 119 175 204
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -61 51 -27 68
rect -61 -68 -27 -51
rect 27 51 61 68
rect 27 -68 61 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -204 -141 -119
rect -33 -136 -17 -102
rect 17 -136 33 -102
rect 141 -204 175 -119
rect -175 -238 -51 -204
rect -17 -238 17 -204
rect 51 -238 175 -204
<< viali >>
rect -17 102 17 136
rect -61 -17 -27 17
rect 27 -17 61 17
rect -17 -136 17 -102
<< metal1 >>
rect -29 136 29 142
rect -29 102 -17 136
rect 17 102 29 136
rect -29 96 29 102
rect -67 17 -21 64
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -64 -21 -17
rect 21 17 67 64
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -64 67 -17
rect -29 -102 29 -96
rect -29 -136 -17 -102
rect 17 -136 29 -102
rect -29 -142 29 -136
<< properties >>
string FIXED_BBOX -158 -221 158 221
<< end >>
