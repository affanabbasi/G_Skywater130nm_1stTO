magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -165 986 165 1020
rect -165 -986 -131 986
rect 131 -986 165 986
rect -165 -1020 165 -986
<< psubdiff >>
rect -165 986 -51 1020
rect -17 986 17 1020
rect 51 986 165 1020
rect -165 901 -131 986
rect 131 901 165 986
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect -165 -986 -131 -901
rect 131 -986 165 -901
rect -165 -1020 -51 -986
rect -17 -1020 17 -986
rect 51 -1020 165 -986
<< psubdiffcont >>
rect -51 986 -17 1020
rect 17 986 51 1020
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect -51 -1020 -17 -986
rect 17 -1020 51 -986
<< xpolycontact >>
rect -35 458 35 890
rect -35 -890 35 -458
<< xpolyres >>
rect -35 -458 35 458
<< locali >>
rect -165 986 -51 1020
rect -17 986 17 1020
rect 51 986 165 1020
rect -165 901 -131 986
rect 131 901 165 986
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect -165 -986 -131 -901
rect 131 -986 165 -901
rect -165 -1020 -51 -986
rect -17 -1020 17 -986
rect 51 -1020 165 -986
<< viali >>
rect -17 836 17 870
rect -17 764 17 798
rect -17 692 17 726
rect -17 620 17 654
rect -17 548 17 582
rect -17 476 17 510
rect -17 -511 17 -477
rect -17 -583 17 -549
rect -17 -655 17 -621
rect -17 -727 17 -693
rect -17 -799 17 -765
rect -17 -871 17 -837
<< metal1 >>
rect -25 870 25 884
rect -25 836 -17 870
rect 17 836 25 870
rect -25 798 25 836
rect -25 764 -17 798
rect 17 764 25 798
rect -25 726 25 764
rect -25 692 -17 726
rect 17 692 25 726
rect -25 654 25 692
rect -25 620 -17 654
rect 17 620 25 654
rect -25 582 25 620
rect -25 548 -17 582
rect 17 548 25 582
rect -25 510 25 548
rect -25 476 -17 510
rect 17 476 25 510
rect -25 463 25 476
rect -25 -477 25 -463
rect -25 -511 -17 -477
rect 17 -511 25 -477
rect -25 -549 25 -511
rect -25 -583 -17 -549
rect 17 -583 25 -549
rect -25 -621 25 -583
rect -25 -655 -17 -621
rect 17 -655 25 -621
rect -25 -693 25 -655
rect -25 -727 -17 -693
rect 17 -727 25 -693
rect -25 -765 25 -727
rect -25 -799 -17 -765
rect 17 -799 25 -765
rect -25 -837 25 -799
rect -25 -871 -17 -837
rect 17 -871 25 -837
rect -25 -884 25 -871
<< properties >>
string FIXED_BBOX -148 -1003 148 1003
<< end >>
