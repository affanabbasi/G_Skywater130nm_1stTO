magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< locali >>
rect 4606 448 4641 449
rect 4640 414 4641 448
rect 13236 448 13271 449
rect 13270 414 13271 448
rect 21862 448 21897 449
rect 21896 414 21897 448
rect 30493 448 30530 449
rect 30493 414 30494 448
rect 30528 414 30530 448
<< viali >>
rect 4606 414 4640 448
rect 13236 414 13270 448
rect 21862 414 21896 448
rect 30494 414 30528 448
<< metal1 >>
rect 3562 5717 6706 5740
rect 3562 5665 3572 5717
rect 3624 5665 3636 5717
rect 3688 5665 3700 5717
rect 3752 5665 3764 5717
rect 3816 5665 3828 5717
rect 3880 5665 3892 5717
rect 3944 5665 3956 5717
rect 4008 5665 4020 5717
rect 4072 5665 4084 5717
rect 4136 5665 4148 5717
rect 4200 5665 4212 5717
rect 4264 5665 4276 5717
rect 4328 5665 4340 5717
rect 4392 5665 4404 5717
rect 4456 5665 4468 5717
rect 4520 5665 4532 5717
rect 4584 5665 4596 5717
rect 4648 5665 4660 5717
rect 4712 5665 4724 5717
rect 4776 5665 4788 5717
rect 4840 5665 4852 5717
rect 4904 5665 4916 5717
rect 4968 5665 4980 5717
rect 5032 5665 5044 5717
rect 5096 5665 5108 5717
rect 5160 5665 5172 5717
rect 5224 5665 5236 5717
rect 5288 5665 5300 5717
rect 5352 5665 5364 5717
rect 5416 5665 5428 5717
rect 5480 5665 5492 5717
rect 5544 5665 5556 5717
rect 5608 5665 5620 5717
rect 5672 5665 5684 5717
rect 5736 5665 5748 5717
rect 5800 5665 5812 5717
rect 5864 5665 5876 5717
rect 5928 5665 5940 5717
rect 5992 5665 6004 5717
rect 6056 5665 6068 5717
rect 6120 5665 6132 5717
rect 6184 5665 6196 5717
rect 6248 5665 6260 5717
rect 6312 5665 6324 5717
rect 6376 5665 6388 5717
rect 6440 5665 6452 5717
rect 6504 5665 6516 5717
rect 6568 5665 6580 5717
rect 6632 5665 6644 5717
rect 6696 5665 6706 5717
rect 3562 5642 6706 5665
rect 12187 5717 15331 5740
rect 12187 5665 12197 5717
rect 12249 5665 12261 5717
rect 12313 5665 12325 5717
rect 12377 5665 12389 5717
rect 12441 5665 12453 5717
rect 12505 5665 12517 5717
rect 12569 5665 12581 5717
rect 12633 5665 12645 5717
rect 12697 5665 12709 5717
rect 12761 5665 12773 5717
rect 12825 5665 12837 5717
rect 12889 5665 12901 5717
rect 12953 5665 12965 5717
rect 13017 5665 13029 5717
rect 13081 5665 13093 5717
rect 13145 5665 13157 5717
rect 13209 5665 13221 5717
rect 13273 5665 13285 5717
rect 13337 5665 13349 5717
rect 13401 5665 13413 5717
rect 13465 5665 13477 5717
rect 13529 5665 13541 5717
rect 13593 5665 13605 5717
rect 13657 5665 13669 5717
rect 13721 5665 13733 5717
rect 13785 5665 13797 5717
rect 13849 5665 13861 5717
rect 13913 5665 13925 5717
rect 13977 5665 13989 5717
rect 14041 5665 14053 5717
rect 14105 5665 14117 5717
rect 14169 5665 14181 5717
rect 14233 5665 14245 5717
rect 14297 5665 14309 5717
rect 14361 5665 14373 5717
rect 14425 5665 14437 5717
rect 14489 5665 14501 5717
rect 14553 5665 14565 5717
rect 14617 5665 14629 5717
rect 14681 5665 14693 5717
rect 14745 5665 14757 5717
rect 14809 5665 14821 5717
rect 14873 5665 14885 5717
rect 14937 5665 14949 5717
rect 15001 5665 15013 5717
rect 15065 5665 15077 5717
rect 15129 5665 15141 5717
rect 15193 5665 15205 5717
rect 15257 5665 15269 5717
rect 15321 5665 15331 5717
rect 12187 5642 15331 5665
rect 20812 5717 23956 5740
rect 20812 5665 20822 5717
rect 20874 5665 20886 5717
rect 20938 5665 20950 5717
rect 21002 5665 21014 5717
rect 21066 5665 21078 5717
rect 21130 5665 21142 5717
rect 21194 5665 21206 5717
rect 21258 5665 21270 5717
rect 21322 5665 21334 5717
rect 21386 5665 21398 5717
rect 21450 5665 21462 5717
rect 21514 5665 21526 5717
rect 21578 5665 21590 5717
rect 21642 5665 21654 5717
rect 21706 5665 21718 5717
rect 21770 5665 21782 5717
rect 21834 5665 21846 5717
rect 21898 5665 21910 5717
rect 21962 5665 21974 5717
rect 22026 5665 22038 5717
rect 22090 5665 22102 5717
rect 22154 5665 22166 5717
rect 22218 5665 22230 5717
rect 22282 5665 22294 5717
rect 22346 5665 22358 5717
rect 22410 5665 22422 5717
rect 22474 5665 22486 5717
rect 22538 5665 22550 5717
rect 22602 5665 22614 5717
rect 22666 5665 22678 5717
rect 22730 5665 22742 5717
rect 22794 5665 22806 5717
rect 22858 5665 22870 5717
rect 22922 5665 22934 5717
rect 22986 5665 22998 5717
rect 23050 5665 23062 5717
rect 23114 5665 23126 5717
rect 23178 5665 23190 5717
rect 23242 5665 23254 5717
rect 23306 5665 23318 5717
rect 23370 5665 23382 5717
rect 23434 5665 23446 5717
rect 23498 5665 23510 5717
rect 23562 5665 23574 5717
rect 23626 5665 23638 5717
rect 23690 5665 23702 5717
rect 23754 5665 23766 5717
rect 23818 5665 23830 5717
rect 23882 5665 23894 5717
rect 23946 5665 23956 5717
rect 20812 5642 23956 5665
rect 29436 5717 32580 5740
rect 29436 5665 29446 5717
rect 29498 5665 29510 5717
rect 29562 5665 29574 5717
rect 29626 5665 29638 5717
rect 29690 5665 29702 5717
rect 29754 5665 29766 5717
rect 29818 5665 29830 5717
rect 29882 5665 29894 5717
rect 29946 5665 29958 5717
rect 30010 5665 30022 5717
rect 30074 5665 30086 5717
rect 30138 5665 30150 5717
rect 30202 5665 30214 5717
rect 30266 5665 30278 5717
rect 30330 5665 30342 5717
rect 30394 5665 30406 5717
rect 30458 5665 30470 5717
rect 30522 5665 30534 5717
rect 30586 5665 30598 5717
rect 30650 5665 30662 5717
rect 30714 5665 30726 5717
rect 30778 5665 30790 5717
rect 30842 5665 30854 5717
rect 30906 5665 30918 5717
rect 30970 5665 30982 5717
rect 31034 5665 31046 5717
rect 31098 5665 31110 5717
rect 31162 5665 31174 5717
rect 31226 5665 31238 5717
rect 31290 5665 31302 5717
rect 31354 5665 31366 5717
rect 31418 5665 31430 5717
rect 31482 5665 31494 5717
rect 31546 5665 31558 5717
rect 31610 5665 31622 5717
rect 31674 5665 31686 5717
rect 31738 5665 31750 5717
rect 31802 5665 31814 5717
rect 31866 5665 31878 5717
rect 31930 5665 31942 5717
rect 31994 5665 32006 5717
rect 32058 5665 32070 5717
rect 32122 5665 32134 5717
rect 32186 5665 32198 5717
rect 32250 5665 32262 5717
rect 32314 5665 32326 5717
rect 32378 5665 32390 5717
rect 32442 5665 32454 5717
rect 32506 5665 32518 5717
rect 32570 5665 32580 5717
rect 29436 5642 32580 5665
rect 37846 5717 40990 5740
rect 37846 5665 37856 5717
rect 37908 5665 37920 5717
rect 37972 5665 37984 5717
rect 38036 5665 38048 5717
rect 38100 5665 38112 5717
rect 38164 5665 38176 5717
rect 38228 5665 38240 5717
rect 38292 5665 38304 5717
rect 38356 5665 38368 5717
rect 38420 5665 38432 5717
rect 38484 5665 38496 5717
rect 38548 5665 38560 5717
rect 38612 5665 38624 5717
rect 38676 5665 38688 5717
rect 38740 5665 38752 5717
rect 38804 5665 38816 5717
rect 38868 5665 38880 5717
rect 38932 5665 38944 5717
rect 38996 5665 39008 5717
rect 39060 5665 39072 5717
rect 39124 5665 39136 5717
rect 39188 5665 39200 5717
rect 39252 5665 39264 5717
rect 39316 5665 39328 5717
rect 39380 5665 39392 5717
rect 39444 5665 39456 5717
rect 39508 5665 39520 5717
rect 39572 5665 39584 5717
rect 39636 5665 39648 5717
rect 39700 5665 39712 5717
rect 39764 5665 39776 5717
rect 39828 5665 39840 5717
rect 39892 5665 39904 5717
rect 39956 5665 39968 5717
rect 40020 5665 40032 5717
rect 40084 5665 40096 5717
rect 40148 5665 40160 5717
rect 40212 5665 40224 5717
rect 40276 5665 40288 5717
rect 40340 5665 40352 5717
rect 40404 5665 40416 5717
rect 40468 5665 40480 5717
rect 40532 5665 40544 5717
rect 40596 5665 40608 5717
rect 40660 5665 40672 5717
rect 40724 5665 40736 5717
rect 40788 5665 40800 5717
rect 40852 5665 40864 5717
rect 40916 5665 40928 5717
rect 40980 5665 40990 5717
rect 37846 5642 40990 5665
rect 5604 5172 5984 5201
rect 5604 4992 5640 5172
rect 5948 4992 5984 5172
rect 5604 4964 5984 4992
rect 5663 4000 5922 4964
rect 6409 4697 6668 5642
rect 14053 5111 14433 5140
rect 14053 4931 14089 5111
rect 14397 4931 14433 5111
rect 14053 4903 14433 4931
rect 6348 4668 6728 4697
rect 6348 4488 6384 4668
rect 6692 4488 6728 4668
rect 6348 4460 6728 4488
rect 14117 4000 14376 4903
rect 14906 4774 15165 5642
rect 22852 5262 23232 5291
rect 22852 5082 22888 5262
rect 23196 5082 23232 5262
rect 22852 5054 23232 5082
rect 14843 4745 15223 4774
rect 14843 4565 14879 4745
rect 15187 4565 15223 4745
rect 14843 4537 15223 4565
rect 22901 4000 23160 5054
rect 23611 4546 23870 5642
rect 31511 5246 31891 5275
rect 31511 5066 31547 5246
rect 31855 5066 31891 5246
rect 31511 5038 31891 5066
rect 23523 4517 23903 4546
rect 23523 4337 23559 4517
rect 23867 4337 23903 4517
rect 23523 4309 23903 4337
rect 31566 4000 31825 5038
rect 32289 4546 32548 5642
rect 32223 4517 32603 4546
rect 32223 4337 32259 4517
rect 32567 4337 32603 4517
rect 32223 4309 32603 4337
rect 3558 3977 6702 4000
rect 3558 3925 3568 3977
rect 3620 3925 3632 3977
rect 3684 3925 3696 3977
rect 3748 3925 3760 3977
rect 3812 3925 3824 3977
rect 3876 3925 3888 3977
rect 3940 3925 3952 3977
rect 4004 3925 4016 3977
rect 4068 3925 4080 3977
rect 4132 3925 4144 3977
rect 4196 3925 4208 3977
rect 4260 3925 4272 3977
rect 4324 3925 4336 3977
rect 4388 3925 4400 3977
rect 4452 3925 4464 3977
rect 4516 3925 4528 3977
rect 4580 3925 4592 3977
rect 4644 3925 4656 3977
rect 4708 3925 4720 3977
rect 4772 3925 4784 3977
rect 4836 3925 4848 3977
rect 4900 3925 4912 3977
rect 4964 3925 4976 3977
rect 5028 3925 5040 3977
rect 5092 3925 5104 3977
rect 5156 3925 5168 3977
rect 5220 3925 5232 3977
rect 5284 3925 5296 3977
rect 5348 3925 5360 3977
rect 5412 3925 5424 3977
rect 5476 3925 5488 3977
rect 5540 3925 5552 3977
rect 5604 3925 5616 3977
rect 5668 3925 5680 3977
rect 5732 3925 5744 3977
rect 5796 3925 5808 3977
rect 5860 3925 5872 3977
rect 5924 3925 5936 3977
rect 5988 3925 6000 3977
rect 6052 3925 6064 3977
rect 6116 3925 6128 3977
rect 6180 3925 6192 3977
rect 6244 3925 6256 3977
rect 6308 3925 6320 3977
rect 6372 3925 6384 3977
rect 6436 3925 6448 3977
rect 6500 3925 6512 3977
rect 6564 3925 6576 3977
rect 6628 3925 6640 3977
rect 6692 3925 6702 3977
rect 3558 3902 6702 3925
rect 12183 3977 15327 4000
rect 12183 3925 12193 3977
rect 12245 3925 12257 3977
rect 12309 3925 12321 3977
rect 12373 3925 12385 3977
rect 12437 3925 12449 3977
rect 12501 3925 12513 3977
rect 12565 3925 12577 3977
rect 12629 3925 12641 3977
rect 12693 3925 12705 3977
rect 12757 3925 12769 3977
rect 12821 3925 12833 3977
rect 12885 3925 12897 3977
rect 12949 3925 12961 3977
rect 13013 3925 13025 3977
rect 13077 3925 13089 3977
rect 13141 3925 13153 3977
rect 13205 3925 13217 3977
rect 13269 3925 13281 3977
rect 13333 3925 13345 3977
rect 13397 3925 13409 3977
rect 13461 3925 13473 3977
rect 13525 3925 13537 3977
rect 13589 3925 13601 3977
rect 13653 3925 13665 3977
rect 13717 3925 13729 3977
rect 13781 3925 13793 3977
rect 13845 3925 13857 3977
rect 13909 3925 13921 3977
rect 13973 3925 13985 3977
rect 14037 3925 14049 3977
rect 14101 3925 14113 3977
rect 14165 3925 14177 3977
rect 14229 3925 14241 3977
rect 14293 3925 14305 3977
rect 14357 3925 14369 3977
rect 14421 3925 14433 3977
rect 14485 3925 14497 3977
rect 14549 3925 14561 3977
rect 14613 3925 14625 3977
rect 14677 3925 14689 3977
rect 14741 3925 14753 3977
rect 14805 3925 14817 3977
rect 14869 3925 14881 3977
rect 14933 3925 14945 3977
rect 14997 3925 15009 3977
rect 15061 3925 15073 3977
rect 15125 3925 15137 3977
rect 15189 3925 15201 3977
rect 15253 3925 15265 3977
rect 15317 3925 15327 3977
rect 12183 3902 15327 3925
rect 20808 3977 23952 4000
rect 20808 3925 20818 3977
rect 20870 3925 20882 3977
rect 20934 3925 20946 3977
rect 20998 3925 21010 3977
rect 21062 3925 21074 3977
rect 21126 3925 21138 3977
rect 21190 3925 21202 3977
rect 21254 3925 21266 3977
rect 21318 3925 21330 3977
rect 21382 3925 21394 3977
rect 21446 3925 21458 3977
rect 21510 3925 21522 3977
rect 21574 3925 21586 3977
rect 21638 3925 21650 3977
rect 21702 3925 21714 3977
rect 21766 3925 21778 3977
rect 21830 3925 21842 3977
rect 21894 3925 21906 3977
rect 21958 3925 21970 3977
rect 22022 3925 22034 3977
rect 22086 3925 22098 3977
rect 22150 3925 22162 3977
rect 22214 3925 22226 3977
rect 22278 3925 22290 3977
rect 22342 3925 22354 3977
rect 22406 3925 22418 3977
rect 22470 3925 22482 3977
rect 22534 3925 22546 3977
rect 22598 3925 22610 3977
rect 22662 3925 22674 3977
rect 22726 3925 22738 3977
rect 22790 3925 22802 3977
rect 22854 3925 22866 3977
rect 22918 3925 22930 3977
rect 22982 3925 22994 3977
rect 23046 3925 23058 3977
rect 23110 3925 23122 3977
rect 23174 3925 23186 3977
rect 23238 3925 23250 3977
rect 23302 3925 23314 3977
rect 23366 3925 23378 3977
rect 23430 3925 23442 3977
rect 23494 3925 23506 3977
rect 23558 3925 23570 3977
rect 23622 3925 23634 3977
rect 23686 3925 23698 3977
rect 23750 3925 23762 3977
rect 23814 3925 23826 3977
rect 23878 3925 23890 3977
rect 23942 3925 23952 3977
rect 20808 3902 23952 3925
rect 29433 3977 32577 4000
rect 29433 3925 29443 3977
rect 29495 3925 29507 3977
rect 29559 3925 29571 3977
rect 29623 3925 29635 3977
rect 29687 3925 29699 3977
rect 29751 3925 29763 3977
rect 29815 3925 29827 3977
rect 29879 3925 29891 3977
rect 29943 3925 29955 3977
rect 30007 3925 30019 3977
rect 30071 3925 30083 3977
rect 30135 3925 30147 3977
rect 30199 3925 30211 3977
rect 30263 3925 30275 3977
rect 30327 3925 30339 3977
rect 30391 3925 30403 3977
rect 30455 3925 30467 3977
rect 30519 3925 30531 3977
rect 30583 3925 30595 3977
rect 30647 3925 30659 3977
rect 30711 3925 30723 3977
rect 30775 3925 30787 3977
rect 30839 3925 30851 3977
rect 30903 3925 30915 3977
rect 30967 3925 30979 3977
rect 31031 3925 31043 3977
rect 31095 3925 31107 3977
rect 31159 3925 31171 3977
rect 31223 3925 31235 3977
rect 31287 3925 31299 3977
rect 31351 3925 31363 3977
rect 31415 3925 31427 3977
rect 31479 3925 31491 3977
rect 31543 3925 31555 3977
rect 31607 3925 31619 3977
rect 31671 3925 31683 3977
rect 31735 3925 31747 3977
rect 31799 3925 31811 3977
rect 31863 3925 31875 3977
rect 31927 3925 31939 3977
rect 31991 3925 32003 3977
rect 32055 3925 32067 3977
rect 32119 3925 32131 3977
rect 32183 3925 32195 3977
rect 32247 3925 32259 3977
rect 32311 3925 32323 3977
rect 32375 3925 32387 3977
rect 32439 3925 32451 3977
rect 32503 3925 32515 3977
rect 32567 3925 32577 3977
rect 29433 3902 32577 3925
rect 37846 3977 40990 4000
rect 37846 3925 37856 3977
rect 37908 3925 37920 3977
rect 37972 3925 37984 3977
rect 38036 3925 38048 3977
rect 38100 3925 38112 3977
rect 38164 3925 38176 3977
rect 38228 3925 38240 3977
rect 38292 3925 38304 3977
rect 38356 3925 38368 3977
rect 38420 3925 38432 3977
rect 38484 3925 38496 3977
rect 38548 3925 38560 3977
rect 38612 3925 38624 3977
rect 38676 3925 38688 3977
rect 38740 3925 38752 3977
rect 38804 3925 38816 3977
rect 38868 3925 38880 3977
rect 38932 3925 38944 3977
rect 38996 3925 39008 3977
rect 39060 3925 39072 3977
rect 39124 3925 39136 3977
rect 39188 3925 39200 3977
rect 39252 3925 39264 3977
rect 39316 3925 39328 3977
rect 39380 3925 39392 3977
rect 39444 3925 39456 3977
rect 39508 3925 39520 3977
rect 39572 3925 39584 3977
rect 39636 3925 39648 3977
rect 39700 3925 39712 3977
rect 39764 3925 39776 3977
rect 39828 3925 39840 3977
rect 39892 3925 39904 3977
rect 39956 3925 39968 3977
rect 40020 3925 40032 3977
rect 40084 3925 40096 3977
rect 40148 3925 40160 3977
rect 40212 3925 40224 3977
rect 40276 3925 40288 3977
rect 40340 3925 40352 3977
rect 40404 3925 40416 3977
rect 40468 3925 40480 3977
rect 40532 3925 40544 3977
rect 40596 3925 40608 3977
rect 40660 3925 40672 3977
rect 40724 3925 40736 3977
rect 40788 3925 40800 3977
rect 40852 3925 40864 3977
rect 40916 3925 40928 3977
rect 40980 3925 40990 3977
rect 37846 3902 40990 3925
rect 4594 452 4653 455
rect 4594 448 9042 452
rect 4594 414 4606 448
rect 4640 414 9042 448
rect 4594 384 9042 414
rect 13224 448 13311 482
rect 21850 452 21909 455
rect 30481 452 30542 455
rect 21840 448 25883 452
rect 13224 414 13236 448
rect 13270 414 17260 448
rect 13224 385 17260 414
rect 13224 384 13271 385
rect 13643 380 17260 385
rect 21840 414 21862 448
rect 21896 414 25883 448
rect 21840 384 25883 414
rect 30481 448 34293 452
rect 30481 414 30494 448
rect 30528 414 34293 448
rect 30481 384 34293 414
<< via1 >>
rect 3572 5665 3624 5717
rect 3636 5665 3688 5717
rect 3700 5665 3752 5717
rect 3764 5665 3816 5717
rect 3828 5665 3880 5717
rect 3892 5665 3944 5717
rect 3956 5665 4008 5717
rect 4020 5665 4072 5717
rect 4084 5665 4136 5717
rect 4148 5665 4200 5717
rect 4212 5665 4264 5717
rect 4276 5665 4328 5717
rect 4340 5665 4392 5717
rect 4404 5665 4456 5717
rect 4468 5665 4520 5717
rect 4532 5665 4584 5717
rect 4596 5665 4648 5717
rect 4660 5665 4712 5717
rect 4724 5665 4776 5717
rect 4788 5665 4840 5717
rect 4852 5665 4904 5717
rect 4916 5665 4968 5717
rect 4980 5665 5032 5717
rect 5044 5665 5096 5717
rect 5108 5665 5160 5717
rect 5172 5665 5224 5717
rect 5236 5665 5288 5717
rect 5300 5665 5352 5717
rect 5364 5665 5416 5717
rect 5428 5665 5480 5717
rect 5492 5665 5544 5717
rect 5556 5665 5608 5717
rect 5620 5665 5672 5717
rect 5684 5665 5736 5717
rect 5748 5665 5800 5717
rect 5812 5665 5864 5717
rect 5876 5665 5928 5717
rect 5940 5665 5992 5717
rect 6004 5665 6056 5717
rect 6068 5665 6120 5717
rect 6132 5665 6184 5717
rect 6196 5665 6248 5717
rect 6260 5665 6312 5717
rect 6324 5665 6376 5717
rect 6388 5665 6440 5717
rect 6452 5665 6504 5717
rect 6516 5665 6568 5717
rect 6580 5665 6632 5717
rect 6644 5665 6696 5717
rect 12197 5665 12249 5717
rect 12261 5665 12313 5717
rect 12325 5665 12377 5717
rect 12389 5665 12441 5717
rect 12453 5665 12505 5717
rect 12517 5665 12569 5717
rect 12581 5665 12633 5717
rect 12645 5665 12697 5717
rect 12709 5665 12761 5717
rect 12773 5665 12825 5717
rect 12837 5665 12889 5717
rect 12901 5665 12953 5717
rect 12965 5665 13017 5717
rect 13029 5665 13081 5717
rect 13093 5665 13145 5717
rect 13157 5665 13209 5717
rect 13221 5665 13273 5717
rect 13285 5665 13337 5717
rect 13349 5665 13401 5717
rect 13413 5665 13465 5717
rect 13477 5665 13529 5717
rect 13541 5665 13593 5717
rect 13605 5665 13657 5717
rect 13669 5665 13721 5717
rect 13733 5665 13785 5717
rect 13797 5665 13849 5717
rect 13861 5665 13913 5717
rect 13925 5665 13977 5717
rect 13989 5665 14041 5717
rect 14053 5665 14105 5717
rect 14117 5665 14169 5717
rect 14181 5665 14233 5717
rect 14245 5665 14297 5717
rect 14309 5665 14361 5717
rect 14373 5665 14425 5717
rect 14437 5665 14489 5717
rect 14501 5665 14553 5717
rect 14565 5665 14617 5717
rect 14629 5665 14681 5717
rect 14693 5665 14745 5717
rect 14757 5665 14809 5717
rect 14821 5665 14873 5717
rect 14885 5665 14937 5717
rect 14949 5665 15001 5717
rect 15013 5665 15065 5717
rect 15077 5665 15129 5717
rect 15141 5665 15193 5717
rect 15205 5665 15257 5717
rect 15269 5665 15321 5717
rect 20822 5665 20874 5717
rect 20886 5665 20938 5717
rect 20950 5665 21002 5717
rect 21014 5665 21066 5717
rect 21078 5665 21130 5717
rect 21142 5665 21194 5717
rect 21206 5665 21258 5717
rect 21270 5665 21322 5717
rect 21334 5665 21386 5717
rect 21398 5665 21450 5717
rect 21462 5665 21514 5717
rect 21526 5665 21578 5717
rect 21590 5665 21642 5717
rect 21654 5665 21706 5717
rect 21718 5665 21770 5717
rect 21782 5665 21834 5717
rect 21846 5665 21898 5717
rect 21910 5665 21962 5717
rect 21974 5665 22026 5717
rect 22038 5665 22090 5717
rect 22102 5665 22154 5717
rect 22166 5665 22218 5717
rect 22230 5665 22282 5717
rect 22294 5665 22346 5717
rect 22358 5665 22410 5717
rect 22422 5665 22474 5717
rect 22486 5665 22538 5717
rect 22550 5665 22602 5717
rect 22614 5665 22666 5717
rect 22678 5665 22730 5717
rect 22742 5665 22794 5717
rect 22806 5665 22858 5717
rect 22870 5665 22922 5717
rect 22934 5665 22986 5717
rect 22998 5665 23050 5717
rect 23062 5665 23114 5717
rect 23126 5665 23178 5717
rect 23190 5665 23242 5717
rect 23254 5665 23306 5717
rect 23318 5665 23370 5717
rect 23382 5665 23434 5717
rect 23446 5665 23498 5717
rect 23510 5665 23562 5717
rect 23574 5665 23626 5717
rect 23638 5665 23690 5717
rect 23702 5665 23754 5717
rect 23766 5665 23818 5717
rect 23830 5665 23882 5717
rect 23894 5665 23946 5717
rect 29446 5665 29498 5717
rect 29510 5665 29562 5717
rect 29574 5665 29626 5717
rect 29638 5665 29690 5717
rect 29702 5665 29754 5717
rect 29766 5665 29818 5717
rect 29830 5665 29882 5717
rect 29894 5665 29946 5717
rect 29958 5665 30010 5717
rect 30022 5665 30074 5717
rect 30086 5665 30138 5717
rect 30150 5665 30202 5717
rect 30214 5665 30266 5717
rect 30278 5665 30330 5717
rect 30342 5665 30394 5717
rect 30406 5665 30458 5717
rect 30470 5665 30522 5717
rect 30534 5665 30586 5717
rect 30598 5665 30650 5717
rect 30662 5665 30714 5717
rect 30726 5665 30778 5717
rect 30790 5665 30842 5717
rect 30854 5665 30906 5717
rect 30918 5665 30970 5717
rect 30982 5665 31034 5717
rect 31046 5665 31098 5717
rect 31110 5665 31162 5717
rect 31174 5665 31226 5717
rect 31238 5665 31290 5717
rect 31302 5665 31354 5717
rect 31366 5665 31418 5717
rect 31430 5665 31482 5717
rect 31494 5665 31546 5717
rect 31558 5665 31610 5717
rect 31622 5665 31674 5717
rect 31686 5665 31738 5717
rect 31750 5665 31802 5717
rect 31814 5665 31866 5717
rect 31878 5665 31930 5717
rect 31942 5665 31994 5717
rect 32006 5665 32058 5717
rect 32070 5665 32122 5717
rect 32134 5665 32186 5717
rect 32198 5665 32250 5717
rect 32262 5665 32314 5717
rect 32326 5665 32378 5717
rect 32390 5665 32442 5717
rect 32454 5665 32506 5717
rect 32518 5665 32570 5717
rect 37856 5665 37908 5717
rect 37920 5665 37972 5717
rect 37984 5665 38036 5717
rect 38048 5665 38100 5717
rect 38112 5665 38164 5717
rect 38176 5665 38228 5717
rect 38240 5665 38292 5717
rect 38304 5665 38356 5717
rect 38368 5665 38420 5717
rect 38432 5665 38484 5717
rect 38496 5665 38548 5717
rect 38560 5665 38612 5717
rect 38624 5665 38676 5717
rect 38688 5665 38740 5717
rect 38752 5665 38804 5717
rect 38816 5665 38868 5717
rect 38880 5665 38932 5717
rect 38944 5665 38996 5717
rect 39008 5665 39060 5717
rect 39072 5665 39124 5717
rect 39136 5665 39188 5717
rect 39200 5665 39252 5717
rect 39264 5665 39316 5717
rect 39328 5665 39380 5717
rect 39392 5665 39444 5717
rect 39456 5665 39508 5717
rect 39520 5665 39572 5717
rect 39584 5665 39636 5717
rect 39648 5665 39700 5717
rect 39712 5665 39764 5717
rect 39776 5665 39828 5717
rect 39840 5665 39892 5717
rect 39904 5665 39956 5717
rect 39968 5665 40020 5717
rect 40032 5665 40084 5717
rect 40096 5665 40148 5717
rect 40160 5665 40212 5717
rect 40224 5665 40276 5717
rect 40288 5665 40340 5717
rect 40352 5665 40404 5717
rect 40416 5665 40468 5717
rect 40480 5665 40532 5717
rect 40544 5665 40596 5717
rect 40608 5665 40660 5717
rect 40672 5665 40724 5717
rect 40736 5665 40788 5717
rect 40800 5665 40852 5717
rect 40864 5665 40916 5717
rect 40928 5665 40980 5717
rect 5640 4992 5948 5172
rect 14089 4931 14397 5111
rect 6384 4488 6692 4668
rect 22888 5082 23196 5262
rect 14879 4565 15187 4745
rect 31547 5066 31855 5246
rect 23559 4337 23867 4517
rect 32259 4337 32567 4517
rect 3568 3925 3620 3977
rect 3632 3925 3684 3977
rect 3696 3925 3748 3977
rect 3760 3925 3812 3977
rect 3824 3925 3876 3977
rect 3888 3925 3940 3977
rect 3952 3925 4004 3977
rect 4016 3925 4068 3977
rect 4080 3925 4132 3977
rect 4144 3925 4196 3977
rect 4208 3925 4260 3977
rect 4272 3925 4324 3977
rect 4336 3925 4388 3977
rect 4400 3925 4452 3977
rect 4464 3925 4516 3977
rect 4528 3925 4580 3977
rect 4592 3925 4644 3977
rect 4656 3925 4708 3977
rect 4720 3925 4772 3977
rect 4784 3925 4836 3977
rect 4848 3925 4900 3977
rect 4912 3925 4964 3977
rect 4976 3925 5028 3977
rect 5040 3925 5092 3977
rect 5104 3925 5156 3977
rect 5168 3925 5220 3977
rect 5232 3925 5284 3977
rect 5296 3925 5348 3977
rect 5360 3925 5412 3977
rect 5424 3925 5476 3977
rect 5488 3925 5540 3977
rect 5552 3925 5604 3977
rect 5616 3925 5668 3977
rect 5680 3925 5732 3977
rect 5744 3925 5796 3977
rect 5808 3925 5860 3977
rect 5872 3925 5924 3977
rect 5936 3925 5988 3977
rect 6000 3925 6052 3977
rect 6064 3925 6116 3977
rect 6128 3925 6180 3977
rect 6192 3925 6244 3977
rect 6256 3925 6308 3977
rect 6320 3925 6372 3977
rect 6384 3925 6436 3977
rect 6448 3925 6500 3977
rect 6512 3925 6564 3977
rect 6576 3925 6628 3977
rect 6640 3925 6692 3977
rect 12193 3925 12245 3977
rect 12257 3925 12309 3977
rect 12321 3925 12373 3977
rect 12385 3925 12437 3977
rect 12449 3925 12501 3977
rect 12513 3925 12565 3977
rect 12577 3925 12629 3977
rect 12641 3925 12693 3977
rect 12705 3925 12757 3977
rect 12769 3925 12821 3977
rect 12833 3925 12885 3977
rect 12897 3925 12949 3977
rect 12961 3925 13013 3977
rect 13025 3925 13077 3977
rect 13089 3925 13141 3977
rect 13153 3925 13205 3977
rect 13217 3925 13269 3977
rect 13281 3925 13333 3977
rect 13345 3925 13397 3977
rect 13409 3925 13461 3977
rect 13473 3925 13525 3977
rect 13537 3925 13589 3977
rect 13601 3925 13653 3977
rect 13665 3925 13717 3977
rect 13729 3925 13781 3977
rect 13793 3925 13845 3977
rect 13857 3925 13909 3977
rect 13921 3925 13973 3977
rect 13985 3925 14037 3977
rect 14049 3925 14101 3977
rect 14113 3925 14165 3977
rect 14177 3925 14229 3977
rect 14241 3925 14293 3977
rect 14305 3925 14357 3977
rect 14369 3925 14421 3977
rect 14433 3925 14485 3977
rect 14497 3925 14549 3977
rect 14561 3925 14613 3977
rect 14625 3925 14677 3977
rect 14689 3925 14741 3977
rect 14753 3925 14805 3977
rect 14817 3925 14869 3977
rect 14881 3925 14933 3977
rect 14945 3925 14997 3977
rect 15009 3925 15061 3977
rect 15073 3925 15125 3977
rect 15137 3925 15189 3977
rect 15201 3925 15253 3977
rect 15265 3925 15317 3977
rect 20818 3925 20870 3977
rect 20882 3925 20934 3977
rect 20946 3925 20998 3977
rect 21010 3925 21062 3977
rect 21074 3925 21126 3977
rect 21138 3925 21190 3977
rect 21202 3925 21254 3977
rect 21266 3925 21318 3977
rect 21330 3925 21382 3977
rect 21394 3925 21446 3977
rect 21458 3925 21510 3977
rect 21522 3925 21574 3977
rect 21586 3925 21638 3977
rect 21650 3925 21702 3977
rect 21714 3925 21766 3977
rect 21778 3925 21830 3977
rect 21842 3925 21894 3977
rect 21906 3925 21958 3977
rect 21970 3925 22022 3977
rect 22034 3925 22086 3977
rect 22098 3925 22150 3977
rect 22162 3925 22214 3977
rect 22226 3925 22278 3977
rect 22290 3925 22342 3977
rect 22354 3925 22406 3977
rect 22418 3925 22470 3977
rect 22482 3925 22534 3977
rect 22546 3925 22598 3977
rect 22610 3925 22662 3977
rect 22674 3925 22726 3977
rect 22738 3925 22790 3977
rect 22802 3925 22854 3977
rect 22866 3925 22918 3977
rect 22930 3925 22982 3977
rect 22994 3925 23046 3977
rect 23058 3925 23110 3977
rect 23122 3925 23174 3977
rect 23186 3925 23238 3977
rect 23250 3925 23302 3977
rect 23314 3925 23366 3977
rect 23378 3925 23430 3977
rect 23442 3925 23494 3977
rect 23506 3925 23558 3977
rect 23570 3925 23622 3977
rect 23634 3925 23686 3977
rect 23698 3925 23750 3977
rect 23762 3925 23814 3977
rect 23826 3925 23878 3977
rect 23890 3925 23942 3977
rect 29443 3925 29495 3977
rect 29507 3925 29559 3977
rect 29571 3925 29623 3977
rect 29635 3925 29687 3977
rect 29699 3925 29751 3977
rect 29763 3925 29815 3977
rect 29827 3925 29879 3977
rect 29891 3925 29943 3977
rect 29955 3925 30007 3977
rect 30019 3925 30071 3977
rect 30083 3925 30135 3977
rect 30147 3925 30199 3977
rect 30211 3925 30263 3977
rect 30275 3925 30327 3977
rect 30339 3925 30391 3977
rect 30403 3925 30455 3977
rect 30467 3925 30519 3977
rect 30531 3925 30583 3977
rect 30595 3925 30647 3977
rect 30659 3925 30711 3977
rect 30723 3925 30775 3977
rect 30787 3925 30839 3977
rect 30851 3925 30903 3977
rect 30915 3925 30967 3977
rect 30979 3925 31031 3977
rect 31043 3925 31095 3977
rect 31107 3925 31159 3977
rect 31171 3925 31223 3977
rect 31235 3925 31287 3977
rect 31299 3925 31351 3977
rect 31363 3925 31415 3977
rect 31427 3925 31479 3977
rect 31491 3925 31543 3977
rect 31555 3925 31607 3977
rect 31619 3925 31671 3977
rect 31683 3925 31735 3977
rect 31747 3925 31799 3977
rect 31811 3925 31863 3977
rect 31875 3925 31927 3977
rect 31939 3925 31991 3977
rect 32003 3925 32055 3977
rect 32067 3925 32119 3977
rect 32131 3925 32183 3977
rect 32195 3925 32247 3977
rect 32259 3925 32311 3977
rect 32323 3925 32375 3977
rect 32387 3925 32439 3977
rect 32451 3925 32503 3977
rect 32515 3925 32567 3977
rect 37856 3925 37908 3977
rect 37920 3925 37972 3977
rect 37984 3925 38036 3977
rect 38048 3925 38100 3977
rect 38112 3925 38164 3977
rect 38176 3925 38228 3977
rect 38240 3925 38292 3977
rect 38304 3925 38356 3977
rect 38368 3925 38420 3977
rect 38432 3925 38484 3977
rect 38496 3925 38548 3977
rect 38560 3925 38612 3977
rect 38624 3925 38676 3977
rect 38688 3925 38740 3977
rect 38752 3925 38804 3977
rect 38816 3925 38868 3977
rect 38880 3925 38932 3977
rect 38944 3925 38996 3977
rect 39008 3925 39060 3977
rect 39072 3925 39124 3977
rect 39136 3925 39188 3977
rect 39200 3925 39252 3977
rect 39264 3925 39316 3977
rect 39328 3925 39380 3977
rect 39392 3925 39444 3977
rect 39456 3925 39508 3977
rect 39520 3925 39572 3977
rect 39584 3925 39636 3977
rect 39648 3925 39700 3977
rect 39712 3925 39764 3977
rect 39776 3925 39828 3977
rect 39840 3925 39892 3977
rect 39904 3925 39956 3977
rect 39968 3925 40020 3977
rect 40032 3925 40084 3977
rect 40096 3925 40148 3977
rect 40160 3925 40212 3977
rect 40224 3925 40276 3977
rect 40288 3925 40340 3977
rect 40352 3925 40404 3977
rect 40416 3925 40468 3977
rect 40480 3925 40532 3977
rect 40544 3925 40596 3977
rect 40608 3925 40660 3977
rect 40672 3925 40724 3977
rect 40736 3925 40788 3977
rect 40800 3925 40852 3977
rect 40864 3925 40916 3977
rect 40928 3925 40980 3977
<< metal2 >>
rect 190 10210 39486 10301
rect 39793 5924 40443 5945
rect -2189 5618 -1676 5796
rect 39793 5750 39810 5924
rect 3572 5717 6696 5750
rect 3624 5665 3636 5717
rect 3688 5665 3700 5717
rect 3752 5665 3764 5717
rect 3816 5665 3828 5717
rect 3880 5665 3892 5717
rect 3944 5665 3956 5717
rect 4008 5665 4020 5717
rect 4072 5665 4084 5717
rect 4136 5665 4148 5717
rect 4200 5665 4212 5717
rect 4264 5665 4276 5717
rect 4328 5665 4340 5717
rect 4392 5665 4404 5717
rect 4456 5665 4468 5717
rect 4520 5665 4532 5717
rect 4584 5665 4596 5717
rect 4648 5665 4660 5717
rect 4712 5665 4724 5717
rect 4776 5665 4788 5717
rect 4840 5665 4852 5717
rect 4904 5665 4916 5717
rect 4968 5665 4980 5717
rect 5032 5665 5044 5717
rect 5096 5665 5108 5717
rect 5160 5665 5172 5717
rect 5224 5665 5236 5717
rect 5288 5665 5300 5717
rect 5352 5665 5364 5717
rect 5416 5665 5428 5717
rect 5480 5665 5492 5717
rect 5544 5665 5556 5717
rect 5608 5665 5620 5717
rect 5672 5665 5684 5717
rect 5736 5665 5748 5717
rect 5800 5665 5812 5717
rect 5864 5665 5876 5717
rect 5928 5665 5940 5717
rect 5992 5665 6004 5717
rect 6056 5665 6068 5717
rect 6120 5665 6132 5717
rect 6184 5665 6196 5717
rect 6248 5665 6260 5717
rect 6312 5665 6324 5717
rect 6376 5665 6388 5717
rect 6440 5665 6452 5717
rect 6504 5665 6516 5717
rect 6568 5665 6580 5717
rect 6632 5665 6644 5717
rect 3572 5632 6696 5665
rect 12197 5717 15321 5750
rect 12249 5665 12261 5717
rect 12313 5665 12325 5717
rect 12377 5665 12389 5717
rect 12441 5665 12453 5717
rect 12505 5665 12517 5717
rect 12569 5665 12581 5717
rect 12633 5665 12645 5717
rect 12697 5665 12709 5717
rect 12761 5665 12773 5717
rect 12825 5665 12837 5717
rect 12889 5665 12901 5717
rect 12953 5665 12965 5717
rect 13017 5665 13029 5717
rect 13081 5665 13093 5717
rect 13145 5665 13157 5717
rect 13209 5665 13221 5717
rect 13273 5665 13285 5717
rect 13337 5665 13349 5717
rect 13401 5665 13413 5717
rect 13465 5665 13477 5717
rect 13529 5665 13541 5717
rect 13593 5665 13605 5717
rect 13657 5665 13669 5717
rect 13721 5665 13733 5717
rect 13785 5665 13797 5717
rect 13849 5665 13861 5717
rect 13913 5665 13925 5717
rect 13977 5665 13989 5717
rect 14041 5665 14053 5717
rect 14105 5665 14117 5717
rect 14169 5665 14181 5717
rect 14233 5665 14245 5717
rect 14297 5665 14309 5717
rect 14361 5665 14373 5717
rect 14425 5665 14437 5717
rect 14489 5665 14501 5717
rect 14553 5665 14565 5717
rect 14617 5665 14629 5717
rect 14681 5665 14693 5717
rect 14745 5665 14757 5717
rect 14809 5665 14821 5717
rect 14873 5665 14885 5717
rect 14937 5665 14949 5717
rect 15001 5665 15013 5717
rect 15065 5665 15077 5717
rect 15129 5665 15141 5717
rect 15193 5665 15205 5717
rect 15257 5665 15269 5717
rect 12197 5632 15321 5665
rect 20822 5717 23946 5750
rect 20874 5665 20886 5717
rect 20938 5665 20950 5717
rect 21002 5665 21014 5717
rect 21066 5665 21078 5717
rect 21130 5665 21142 5717
rect 21194 5665 21206 5717
rect 21258 5665 21270 5717
rect 21322 5665 21334 5717
rect 21386 5665 21398 5717
rect 21450 5665 21462 5717
rect 21514 5665 21526 5717
rect 21578 5665 21590 5717
rect 21642 5665 21654 5717
rect 21706 5665 21718 5717
rect 21770 5665 21782 5717
rect 21834 5665 21846 5717
rect 21898 5665 21910 5717
rect 21962 5665 21974 5717
rect 22026 5665 22038 5717
rect 22090 5665 22102 5717
rect 22154 5665 22166 5717
rect 22218 5665 22230 5717
rect 22282 5665 22294 5717
rect 22346 5665 22358 5717
rect 22410 5665 22422 5717
rect 22474 5665 22486 5717
rect 22538 5665 22550 5717
rect 22602 5665 22614 5717
rect 22666 5665 22678 5717
rect 22730 5665 22742 5717
rect 22794 5665 22806 5717
rect 22858 5665 22870 5717
rect 22922 5665 22934 5717
rect 22986 5665 22998 5717
rect 23050 5665 23062 5717
rect 23114 5665 23126 5717
rect 23178 5665 23190 5717
rect 23242 5665 23254 5717
rect 23306 5665 23318 5717
rect 23370 5665 23382 5717
rect 23434 5665 23446 5717
rect 23498 5665 23510 5717
rect 23562 5665 23574 5717
rect 23626 5665 23638 5717
rect 23690 5665 23702 5717
rect 23754 5665 23766 5717
rect 23818 5665 23830 5717
rect 23882 5665 23894 5717
rect 20822 5632 23946 5665
rect 29446 5717 32570 5750
rect 29498 5665 29510 5717
rect 29562 5665 29574 5717
rect 29626 5665 29638 5717
rect 29690 5665 29702 5717
rect 29754 5665 29766 5717
rect 29818 5665 29830 5717
rect 29882 5665 29894 5717
rect 29946 5665 29958 5717
rect 30010 5665 30022 5717
rect 30074 5665 30086 5717
rect 30138 5665 30150 5717
rect 30202 5665 30214 5717
rect 30266 5665 30278 5717
rect 30330 5665 30342 5717
rect 30394 5665 30406 5717
rect 30458 5665 30470 5717
rect 30522 5665 30534 5717
rect 30586 5665 30598 5717
rect 30650 5665 30662 5717
rect 30714 5665 30726 5717
rect 30778 5665 30790 5717
rect 30842 5665 30854 5717
rect 30906 5665 30918 5717
rect 30970 5665 30982 5717
rect 31034 5665 31046 5717
rect 31098 5665 31110 5717
rect 31162 5665 31174 5717
rect 31226 5665 31238 5717
rect 31290 5665 31302 5717
rect 31354 5665 31366 5717
rect 31418 5665 31430 5717
rect 31482 5665 31494 5717
rect 31546 5665 31558 5717
rect 31610 5665 31622 5717
rect 31674 5665 31686 5717
rect 31738 5665 31750 5717
rect 31802 5665 31814 5717
rect 31866 5665 31878 5717
rect 31930 5665 31942 5717
rect 31994 5665 32006 5717
rect 32058 5665 32070 5717
rect 32122 5665 32134 5717
rect 32186 5665 32198 5717
rect 32250 5665 32262 5717
rect 32314 5665 32326 5717
rect 32378 5665 32390 5717
rect 32442 5665 32454 5717
rect 32506 5665 32518 5717
rect 29446 5632 32570 5665
rect 37856 5717 39810 5750
rect 40426 5750 40443 5924
rect 40426 5717 40980 5750
rect 37908 5665 37920 5717
rect 37972 5665 37984 5717
rect 38036 5665 38048 5717
rect 38100 5665 38112 5717
rect 38164 5665 38176 5717
rect 38228 5665 38240 5717
rect 38292 5665 38304 5717
rect 38356 5665 38368 5717
rect 38420 5665 38432 5717
rect 38484 5665 38496 5717
rect 38548 5665 38560 5717
rect 38612 5665 38624 5717
rect 38676 5665 38688 5717
rect 38740 5665 38752 5717
rect 38804 5665 38816 5717
rect 38868 5665 38880 5717
rect 38932 5665 38944 5717
rect 38996 5665 39008 5717
rect 39060 5665 39072 5717
rect 39124 5665 39136 5717
rect 39188 5665 39200 5717
rect 39252 5665 39264 5717
rect 39316 5665 39328 5717
rect 39380 5665 39392 5717
rect 39444 5665 39456 5717
rect 39508 5665 39520 5717
rect 39572 5665 39584 5717
rect 39636 5665 39648 5717
rect 39700 5665 39712 5717
rect 39764 5665 39776 5717
rect 40468 5665 40480 5717
rect 40532 5665 40544 5717
rect 40596 5665 40608 5717
rect 40660 5665 40672 5717
rect 40724 5665 40736 5717
rect 40788 5665 40800 5717
rect 40852 5665 40864 5717
rect 40916 5665 40928 5717
rect 37856 5632 39810 5665
rect -2259 5597 -1609 5618
rect -2259 5141 -2242 5597
rect -1626 5188 -1609 5597
rect 39793 5468 39810 5632
rect 40426 5632 40980 5665
rect 40426 5468 40443 5632
rect 39793 5447 40443 5468
rect 22862 5262 23222 5301
rect -1626 5141 1093 5188
rect -2259 5120 1093 5141
rect -2189 5114 1093 5120
rect 5614 5172 5974 5211
rect -2189 5054 1568 5114
rect -2189 4946 1093 5054
rect 5614 4992 5640 5172
rect 5948 5114 5974 5172
rect 14063 5114 14423 5150
rect 5948 5054 10193 5114
rect 14063 5111 18822 5114
rect 5948 4992 5974 5054
rect 5614 4954 5974 4992
rect -2189 4918 -1676 4946
rect 14063 4931 14089 5111
rect 14397 5054 18822 5111
rect 22862 5082 22888 5262
rect 23196 5114 23222 5262
rect 31521 5246 31881 5285
rect 23196 5082 27443 5114
rect 22862 5054 27443 5082
rect 31521 5066 31547 5246
rect 31855 5114 31881 5246
rect 31855 5066 35856 5114
rect 31521 5054 35856 5066
rect 14397 4931 14423 5054
rect 22862 5044 23222 5054
rect 31521 5028 31881 5054
rect 14063 4893 14423 4931
rect 14853 4745 15213 4784
rect -857 4644 -344 4675
rect 6358 4668 6718 4707
rect -857 4562 1093 4644
rect -857 4502 1564 4562
rect -857 4398 1093 4502
rect 6358 4488 6384 4668
rect 6692 4562 6718 4668
rect 14853 4565 14879 4745
rect 15187 4565 15213 4745
rect 14853 4562 15213 4565
rect 6692 4502 10189 4562
rect 14853 4502 18802 4562
rect 23522 4517 27439 4562
rect 23522 4502 23559 4517
rect 6692 4488 6718 4502
rect 6358 4450 6718 4488
rect -857 4197 -344 4398
rect 23533 4337 23559 4502
rect 23867 4502 27439 4517
rect 32233 4517 35852 4562
rect 23867 4337 23893 4502
rect 23533 4299 23893 4337
rect 32233 4337 32259 4517
rect 32567 4502 35852 4517
rect 32567 4337 32593 4502
rect 32233 4299 32593 4337
rect -923 4176 -273 4197
rect -923 3720 -906 4176
rect -290 3720 -273 4176
rect 40737 4176 41387 4197
rect 40737 4010 40754 4176
rect 3568 3977 6692 4010
rect 3620 3925 3632 3977
rect 3684 3925 3696 3977
rect 3748 3925 3760 3977
rect 3812 3925 3824 3977
rect 3876 3925 3888 3977
rect 3940 3925 3952 3977
rect 4004 3925 4016 3977
rect 4068 3925 4080 3977
rect 4132 3925 4144 3977
rect 4196 3925 4208 3977
rect 4260 3925 4272 3977
rect 4324 3925 4336 3977
rect 4388 3925 4400 3977
rect 4452 3925 4464 3977
rect 4516 3925 4528 3977
rect 4580 3925 4592 3977
rect 4644 3925 4656 3977
rect 4708 3925 4720 3977
rect 4772 3925 4784 3977
rect 4836 3925 4848 3977
rect 4900 3925 4912 3977
rect 4964 3925 4976 3977
rect 5028 3925 5040 3977
rect 5092 3925 5104 3977
rect 5156 3925 5168 3977
rect 5220 3925 5232 3977
rect 5284 3925 5296 3977
rect 5348 3925 5360 3977
rect 5412 3925 5424 3977
rect 5476 3925 5488 3977
rect 5540 3925 5552 3977
rect 5604 3925 5616 3977
rect 5668 3925 5680 3977
rect 5732 3925 5744 3977
rect 5796 3925 5808 3977
rect 5860 3925 5872 3977
rect 5924 3925 5936 3977
rect 5988 3925 6000 3977
rect 6052 3925 6064 3977
rect 6116 3925 6128 3977
rect 6180 3925 6192 3977
rect 6244 3925 6256 3977
rect 6308 3925 6320 3977
rect 6372 3925 6384 3977
rect 6436 3925 6448 3977
rect 6500 3925 6512 3977
rect 6564 3925 6576 3977
rect 6628 3925 6640 3977
rect 3568 3892 6692 3925
rect 12193 3977 15317 4010
rect 12245 3925 12257 3977
rect 12309 3925 12321 3977
rect 12373 3925 12385 3977
rect 12437 3925 12449 3977
rect 12501 3925 12513 3977
rect 12565 3925 12577 3977
rect 12629 3925 12641 3977
rect 12693 3925 12705 3977
rect 12757 3925 12769 3977
rect 12821 3925 12833 3977
rect 12885 3925 12897 3977
rect 12949 3925 12961 3977
rect 13013 3925 13025 3977
rect 13077 3925 13089 3977
rect 13141 3925 13153 3977
rect 13205 3925 13217 3977
rect 13269 3925 13281 3977
rect 13333 3925 13345 3977
rect 13397 3925 13409 3977
rect 13461 3925 13473 3977
rect 13525 3925 13537 3977
rect 13589 3925 13601 3977
rect 13653 3925 13665 3977
rect 13717 3925 13729 3977
rect 13781 3925 13793 3977
rect 13845 3925 13857 3977
rect 13909 3925 13921 3977
rect 13973 3925 13985 3977
rect 14037 3925 14049 3977
rect 14101 3925 14113 3977
rect 14165 3925 14177 3977
rect 14229 3925 14241 3977
rect 14293 3925 14305 3977
rect 14357 3925 14369 3977
rect 14421 3925 14433 3977
rect 14485 3925 14497 3977
rect 14549 3925 14561 3977
rect 14613 3925 14625 3977
rect 14677 3925 14689 3977
rect 14741 3925 14753 3977
rect 14805 3925 14817 3977
rect 14869 3925 14881 3977
rect 14933 3925 14945 3977
rect 14997 3925 15009 3977
rect 15061 3925 15073 3977
rect 15125 3925 15137 3977
rect 15189 3925 15201 3977
rect 15253 3925 15265 3977
rect 12193 3892 15317 3925
rect 20818 3977 23942 4010
rect 20870 3925 20882 3977
rect 20934 3925 20946 3977
rect 20998 3925 21010 3977
rect 21062 3925 21074 3977
rect 21126 3925 21138 3977
rect 21190 3925 21202 3977
rect 21254 3925 21266 3977
rect 21318 3925 21330 3977
rect 21382 3925 21394 3977
rect 21446 3925 21458 3977
rect 21510 3925 21522 3977
rect 21574 3925 21586 3977
rect 21638 3925 21650 3977
rect 21702 3925 21714 3977
rect 21766 3925 21778 3977
rect 21830 3925 21842 3977
rect 21894 3925 21906 3977
rect 21958 3925 21970 3977
rect 22022 3925 22034 3977
rect 22086 3925 22098 3977
rect 22150 3925 22162 3977
rect 22214 3925 22226 3977
rect 22278 3925 22290 3977
rect 22342 3925 22354 3977
rect 22406 3925 22418 3977
rect 22470 3925 22482 3977
rect 22534 3925 22546 3977
rect 22598 3925 22610 3977
rect 22662 3925 22674 3977
rect 22726 3925 22738 3977
rect 22790 3925 22802 3977
rect 22854 3925 22866 3977
rect 22918 3925 22930 3977
rect 22982 3925 22994 3977
rect 23046 3925 23058 3977
rect 23110 3925 23122 3977
rect 23174 3925 23186 3977
rect 23238 3925 23250 3977
rect 23302 3925 23314 3977
rect 23366 3925 23378 3977
rect 23430 3925 23442 3977
rect 23494 3925 23506 3977
rect 23558 3925 23570 3977
rect 23622 3925 23634 3977
rect 23686 3925 23698 3977
rect 23750 3925 23762 3977
rect 23814 3925 23826 3977
rect 23878 3925 23890 3977
rect 20818 3892 23942 3925
rect 29443 3977 32567 4010
rect 29495 3925 29507 3977
rect 29559 3925 29571 3977
rect 29623 3925 29635 3977
rect 29687 3925 29699 3977
rect 29751 3925 29763 3977
rect 29815 3925 29827 3977
rect 29879 3925 29891 3977
rect 29943 3925 29955 3977
rect 30007 3925 30019 3977
rect 30071 3925 30083 3977
rect 30135 3925 30147 3977
rect 30199 3925 30211 3977
rect 30263 3925 30275 3977
rect 30327 3925 30339 3977
rect 30391 3925 30403 3977
rect 30455 3925 30467 3977
rect 30519 3925 30531 3977
rect 30583 3925 30595 3977
rect 30647 3925 30659 3977
rect 30711 3925 30723 3977
rect 30775 3925 30787 3977
rect 30839 3925 30851 3977
rect 30903 3925 30915 3977
rect 30967 3925 30979 3977
rect 31031 3925 31043 3977
rect 31095 3925 31107 3977
rect 31159 3925 31171 3977
rect 31223 3925 31235 3977
rect 31287 3925 31299 3977
rect 31351 3925 31363 3977
rect 31415 3925 31427 3977
rect 31479 3925 31491 3977
rect 31543 3925 31555 3977
rect 31607 3925 31619 3977
rect 31671 3925 31683 3977
rect 31735 3925 31747 3977
rect 31799 3925 31811 3977
rect 31863 3925 31875 3977
rect 31927 3925 31939 3977
rect 31991 3925 32003 3977
rect 32055 3925 32067 3977
rect 32119 3925 32131 3977
rect 32183 3925 32195 3977
rect 32247 3925 32259 3977
rect 32311 3925 32323 3977
rect 32375 3925 32387 3977
rect 32439 3925 32451 3977
rect 32503 3925 32515 3977
rect 29443 3892 32567 3925
rect 37856 3977 40754 4010
rect 37908 3925 37920 3977
rect 37972 3925 37984 3977
rect 38036 3925 38048 3977
rect 38100 3925 38112 3977
rect 38164 3925 38176 3977
rect 38228 3925 38240 3977
rect 38292 3925 38304 3977
rect 38356 3925 38368 3977
rect 38420 3925 38432 3977
rect 38484 3925 38496 3977
rect 38548 3925 38560 3977
rect 38612 3925 38624 3977
rect 38676 3925 38688 3977
rect 38740 3925 38752 3977
rect 38804 3925 38816 3977
rect 38868 3925 38880 3977
rect 38932 3925 38944 3977
rect 38996 3925 39008 3977
rect 39060 3925 39072 3977
rect 39124 3925 39136 3977
rect 39188 3925 39200 3977
rect 39252 3925 39264 3977
rect 39316 3925 39328 3977
rect 39380 3925 39392 3977
rect 39444 3925 39456 3977
rect 39508 3925 39520 3977
rect 39572 3925 39584 3977
rect 39636 3925 39648 3977
rect 39700 3925 39712 3977
rect 39764 3925 39776 3977
rect 39828 3925 39840 3977
rect 39892 3925 39904 3977
rect 39956 3925 39968 3977
rect 40020 3925 40032 3977
rect 40084 3925 40096 3977
rect 40148 3925 40160 3977
rect 40212 3925 40224 3977
rect 40276 3925 40288 3977
rect 40340 3925 40352 3977
rect 40404 3925 40416 3977
rect 40468 3925 40480 3977
rect 40532 3925 40544 3977
rect 40596 3925 40608 3977
rect 40660 3925 40672 3977
rect 40724 3925 40736 3977
rect 37856 3892 40754 3925
rect -923 3699 -273 3720
rect 40737 3720 40754 3892
rect 41370 3720 41387 4176
rect 40737 3699 41387 3720
rect 702 -13 39167 191
<< via2 >>
rect 39810 5717 40426 5924
rect 39810 5665 39828 5717
rect 39828 5665 39840 5717
rect 39840 5665 39892 5717
rect 39892 5665 39904 5717
rect 39904 5665 39956 5717
rect 39956 5665 39968 5717
rect 39968 5665 40020 5717
rect 40020 5665 40032 5717
rect 40032 5665 40084 5717
rect 40084 5665 40096 5717
rect 40096 5665 40148 5717
rect 40148 5665 40160 5717
rect 40160 5665 40212 5717
rect 40212 5665 40224 5717
rect 40224 5665 40276 5717
rect 40276 5665 40288 5717
rect 40288 5665 40340 5717
rect 40340 5665 40352 5717
rect 40352 5665 40404 5717
rect 40404 5665 40416 5717
rect 40416 5665 40426 5717
rect -2242 5141 -1626 5597
rect 39810 5468 40426 5665
rect -906 3720 -290 4176
rect 40754 3977 41370 4176
rect 40754 3925 40788 3977
rect 40788 3925 40800 3977
rect 40800 3925 40852 3977
rect 40852 3925 40864 3977
rect 40864 3925 40916 3977
rect 40916 3925 40928 3977
rect 40928 3925 40980 3977
rect 40980 3925 41370 3977
rect 40754 3720 41370 3925
<< metal3 >>
rect -2269 11844 41397 12427
rect -2269 5597 -1598 11844
rect -2269 5141 -2242 5597
rect -1626 5141 -1598 5597
rect -2269 5120 -1598 5141
rect -933 10751 40451 11216
rect -933 10633 40452 10751
rect -933 4176 -263 10633
rect 0 6320 39656 6406
rect 39783 5940 40452 10633
rect 39783 5924 40453 5940
rect 39783 5468 39810 5924
rect 40426 5468 40453 5924
rect 39783 5452 40453 5468
rect 39783 5447 40452 5452
rect -933 3720 -906 4176
rect -290 3720 -263 4176
rect -933 3699 -263 3720
rect 40727 4176 41397 11844
rect 40727 3720 40754 4176
rect 41370 3720 41397 4176
rect 40727 3699 41397 3720
use DelayCell  DelayCell_1
array 0 3 8625 0 0 693
timestamp 1611881054
transform 1 0 1404 0 1 3676
box -1404 -3676 3964 6620
use DelayCell  DelayCell_0
timestamp 1611881054
transform 1 0 35692 0 1 3676
box -1404 -3676 3964 6620
<< end >>
