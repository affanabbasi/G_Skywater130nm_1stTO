magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< ndiff >>
rect 35469 1159 35503 3135
<< locali >>
rect 29170 3223 38624 3226
rect 29170 3219 29200 3223
rect 29165 3189 29200 3219
rect 29234 3189 29272 3223
rect 29306 3189 29344 3223
rect 29378 3189 29416 3223
rect 29450 3189 29488 3223
rect 29522 3189 29560 3223
rect 29594 3189 29632 3223
rect 29666 3189 29704 3223
rect 29738 3189 29776 3223
rect 29810 3189 29848 3223
rect 29882 3189 29920 3223
rect 29954 3189 29992 3223
rect 30026 3189 30064 3223
rect 30098 3189 30136 3223
rect 30170 3189 30208 3223
rect 30242 3189 30280 3223
rect 30314 3189 30352 3223
rect 30386 3189 30424 3223
rect 30458 3189 30496 3223
rect 30530 3189 30568 3223
rect 30602 3189 30640 3223
rect 30674 3189 30712 3223
rect 30746 3189 30784 3223
rect 30818 3189 30856 3223
rect 30890 3189 30928 3223
rect 30962 3189 31000 3223
rect 31034 3189 31072 3223
rect 31106 3189 31144 3223
rect 31178 3189 31216 3223
rect 31250 3189 31288 3223
rect 31322 3189 31360 3223
rect 31394 3189 31432 3223
rect 31466 3189 31504 3223
rect 31538 3189 31576 3223
rect 31610 3189 31648 3223
rect 31682 3189 31720 3223
rect 31754 3189 31792 3223
rect 31826 3189 31864 3223
rect 31898 3189 31936 3223
rect 31970 3189 32008 3223
rect 32042 3189 32080 3223
rect 32114 3189 32152 3223
rect 32186 3189 32224 3223
rect 32258 3189 32296 3223
rect 32330 3189 32368 3223
rect 32402 3189 32440 3223
rect 32474 3189 32512 3223
rect 32546 3189 32584 3223
rect 32618 3189 32656 3223
rect 32690 3189 32728 3223
rect 32762 3189 32800 3223
rect 32834 3189 32872 3223
rect 32906 3189 32944 3223
rect 32978 3189 33016 3223
rect 33050 3189 33088 3223
rect 33122 3189 33160 3223
rect 33194 3189 33232 3223
rect 33266 3189 33304 3223
rect 33338 3189 33376 3223
rect 33410 3189 33448 3223
rect 33482 3189 33520 3223
rect 33554 3189 33592 3223
rect 33626 3189 33664 3223
rect 33698 3189 33736 3223
rect 33770 3189 33808 3223
rect 33842 3189 33880 3223
rect 33914 3189 33952 3223
rect 33986 3189 34024 3223
rect 34058 3189 34096 3223
rect 34130 3189 34168 3223
rect 34202 3189 34240 3223
rect 34274 3189 34312 3223
rect 34346 3189 34384 3223
rect 34418 3189 34456 3223
rect 34490 3189 34528 3223
rect 34562 3189 34600 3223
rect 34634 3189 34672 3223
rect 34706 3189 34744 3223
rect 34778 3189 34816 3223
rect 34850 3189 34888 3223
rect 34922 3189 34960 3223
rect 34994 3189 35032 3223
rect 35066 3189 35104 3223
rect 35138 3189 35176 3223
rect 35210 3189 35248 3223
rect 35282 3189 35320 3223
rect 35354 3189 35392 3223
rect 35426 3189 35464 3223
rect 35498 3189 35536 3223
rect 35570 3189 35608 3223
rect 35642 3189 35680 3223
rect 35714 3189 35752 3223
rect 35786 3189 35824 3223
rect 35858 3189 35896 3223
rect 35930 3189 35968 3223
rect 36002 3189 36040 3223
rect 36074 3189 36112 3223
rect 36146 3189 36184 3223
rect 36218 3189 36256 3223
rect 36290 3189 36328 3223
rect 36362 3189 36400 3223
rect 36434 3189 36472 3223
rect 36506 3189 36544 3223
rect 36578 3189 36616 3223
rect 36650 3189 36688 3223
rect 36722 3189 36760 3223
rect 36794 3189 36832 3223
rect 36866 3189 36904 3223
rect 36938 3189 36976 3223
rect 37010 3189 37048 3223
rect 37082 3189 37120 3223
rect 37154 3189 37192 3223
rect 37226 3189 37264 3223
rect 37298 3189 37336 3223
rect 37370 3189 37408 3223
rect 37442 3189 37480 3223
rect 37514 3189 37552 3223
rect 37586 3189 37624 3223
rect 37658 3189 37696 3223
rect 37730 3189 37768 3223
rect 37802 3189 37840 3223
rect 37874 3189 37912 3223
rect 37946 3189 37984 3223
rect 38018 3189 38056 3223
rect 38090 3189 38128 3223
rect 38162 3189 38200 3223
rect 38234 3189 38272 3223
rect 38306 3189 38344 3223
rect 38378 3189 38416 3223
rect 38450 3189 38488 3223
rect 38522 3189 38560 3223
rect 38594 3219 38624 3223
rect 38594 3189 38639 3219
rect 29165 3185 38639 3189
rect 29037 3100 29071 3135
rect 29037 3028 29071 3066
rect 29037 2956 29071 2994
rect 29037 2884 29071 2922
rect 29037 2812 29071 2850
rect 29037 2740 29071 2778
rect 29037 2668 29071 2706
rect 29037 2596 29071 2634
rect 29037 2524 29071 2562
rect 29037 2452 29071 2490
rect 29037 2380 29071 2418
rect 29037 2308 29071 2346
rect 29037 2236 29071 2274
rect 29037 2164 29071 2202
rect 29037 2092 29071 2130
rect 29037 2020 29071 2058
rect 29037 1948 29071 1986
rect 29037 1876 29071 1914
rect 29037 1804 29071 1842
rect 29037 1732 29071 1770
rect 29037 1660 29071 1698
rect 29037 1588 29071 1626
rect 29037 1516 29071 1554
rect 29037 1444 29071 1482
rect 29037 1372 29071 1410
rect 29037 1300 29071 1338
rect 29037 1228 29071 1266
rect 29037 1159 29071 1194
rect 29133 3100 29167 3135
rect 29133 3028 29167 3066
rect 29133 2956 29167 2994
rect 29133 2884 29167 2922
rect 29133 2812 29167 2850
rect 29133 2740 29167 2778
rect 29133 2668 29167 2706
rect 29133 2596 29167 2634
rect 29133 2524 29167 2562
rect 29133 2452 29167 2490
rect 29133 2380 29167 2418
rect 29133 2308 29167 2346
rect 29133 2236 29167 2274
rect 29133 2164 29167 2202
rect 29133 2092 29167 2130
rect 29133 2020 29167 2058
rect 29133 1948 29167 1986
rect 29133 1876 29167 1914
rect 29133 1804 29167 1842
rect 29133 1732 29167 1770
rect 29133 1660 29167 1698
rect 29133 1588 29167 1626
rect 29133 1516 29167 1554
rect 29133 1444 29167 1482
rect 29133 1372 29167 1410
rect 29133 1300 29167 1338
rect 29133 1228 29167 1266
rect 29133 1159 29167 1194
rect 29229 3100 29263 3135
rect 29229 3028 29263 3066
rect 29229 2956 29263 2994
rect 29229 2884 29263 2922
rect 29229 2812 29263 2850
rect 29229 2740 29263 2778
rect 29229 2668 29263 2706
rect 29229 2596 29263 2634
rect 29229 2524 29263 2562
rect 29229 2452 29263 2490
rect 29229 2380 29263 2418
rect 29229 2308 29263 2346
rect 29229 2236 29263 2274
rect 29229 2164 29263 2202
rect 29229 2092 29263 2130
rect 29229 2020 29263 2058
rect 29229 1948 29263 1986
rect 29229 1876 29263 1914
rect 29229 1804 29263 1842
rect 29229 1732 29263 1770
rect 29229 1660 29263 1698
rect 29229 1588 29263 1626
rect 29229 1516 29263 1554
rect 29229 1444 29263 1482
rect 29229 1372 29263 1410
rect 29229 1300 29263 1338
rect 29229 1228 29263 1266
rect 29229 1159 29263 1194
rect 29325 3100 29359 3135
rect 29325 3028 29359 3066
rect 29325 2956 29359 2994
rect 29325 2884 29359 2922
rect 29325 2812 29359 2850
rect 29325 2740 29359 2778
rect 29325 2668 29359 2706
rect 29325 2596 29359 2634
rect 29325 2524 29359 2562
rect 29325 2452 29359 2490
rect 29325 2380 29359 2418
rect 29325 2308 29359 2346
rect 29325 2236 29359 2274
rect 29325 2164 29359 2202
rect 29325 2092 29359 2130
rect 29325 2020 29359 2058
rect 29325 1948 29359 1986
rect 29325 1876 29359 1914
rect 29325 1804 29359 1842
rect 29325 1732 29359 1770
rect 29325 1660 29359 1698
rect 29325 1588 29359 1626
rect 29325 1516 29359 1554
rect 29325 1444 29359 1482
rect 29325 1372 29359 1410
rect 29325 1300 29359 1338
rect 29325 1228 29359 1266
rect 29325 1159 29359 1194
rect 29421 3100 29455 3135
rect 29421 3028 29455 3066
rect 29421 2956 29455 2994
rect 29421 2884 29455 2922
rect 29421 2812 29455 2850
rect 29421 2740 29455 2778
rect 29421 2668 29455 2706
rect 29421 2596 29455 2634
rect 29421 2524 29455 2562
rect 29421 2452 29455 2490
rect 29421 2380 29455 2418
rect 29421 2308 29455 2346
rect 29421 2236 29455 2274
rect 29421 2164 29455 2202
rect 29421 2092 29455 2130
rect 29421 2020 29455 2058
rect 29421 1948 29455 1986
rect 29421 1876 29455 1914
rect 29421 1804 29455 1842
rect 29421 1732 29455 1770
rect 29421 1660 29455 1698
rect 29421 1588 29455 1626
rect 29421 1516 29455 1554
rect 29421 1444 29455 1482
rect 29421 1372 29455 1410
rect 29421 1300 29455 1338
rect 29421 1228 29455 1266
rect 29421 1159 29455 1194
rect 29517 3100 29551 3135
rect 29517 3028 29551 3066
rect 29517 2956 29551 2994
rect 29517 2884 29551 2922
rect 29517 2812 29551 2850
rect 29517 2740 29551 2778
rect 29517 2668 29551 2706
rect 29517 2596 29551 2634
rect 29517 2524 29551 2562
rect 29517 2452 29551 2490
rect 29517 2380 29551 2418
rect 29517 2308 29551 2346
rect 29517 2236 29551 2274
rect 29517 2164 29551 2202
rect 29517 2092 29551 2130
rect 29517 2020 29551 2058
rect 29517 1948 29551 1986
rect 29517 1876 29551 1914
rect 29517 1804 29551 1842
rect 29517 1732 29551 1770
rect 29517 1660 29551 1698
rect 29517 1588 29551 1626
rect 29517 1516 29551 1554
rect 29517 1444 29551 1482
rect 29517 1372 29551 1410
rect 29517 1300 29551 1338
rect 29517 1228 29551 1266
rect 29517 1159 29551 1194
rect 29613 3100 29647 3135
rect 29613 3028 29647 3066
rect 29613 2956 29647 2994
rect 29613 2884 29647 2922
rect 29613 2812 29647 2850
rect 29613 2740 29647 2778
rect 29613 2668 29647 2706
rect 29613 2596 29647 2634
rect 29613 2524 29647 2562
rect 29613 2452 29647 2490
rect 29613 2380 29647 2418
rect 29613 2308 29647 2346
rect 29613 2236 29647 2274
rect 29613 2164 29647 2202
rect 29613 2092 29647 2130
rect 29613 2020 29647 2058
rect 29613 1948 29647 1986
rect 29613 1876 29647 1914
rect 29613 1804 29647 1842
rect 29613 1732 29647 1770
rect 29613 1660 29647 1698
rect 29613 1588 29647 1626
rect 29613 1516 29647 1554
rect 29613 1444 29647 1482
rect 29613 1372 29647 1410
rect 29613 1300 29647 1338
rect 29613 1228 29647 1266
rect 29613 1159 29647 1194
rect 29709 3100 29743 3135
rect 29709 3028 29743 3066
rect 29709 2956 29743 2994
rect 29709 2884 29743 2922
rect 29709 2812 29743 2850
rect 29709 2740 29743 2778
rect 29709 2668 29743 2706
rect 29709 2596 29743 2634
rect 29709 2524 29743 2562
rect 29709 2452 29743 2490
rect 29709 2380 29743 2418
rect 29709 2308 29743 2346
rect 29709 2236 29743 2274
rect 29709 2164 29743 2202
rect 29709 2092 29743 2130
rect 29709 2020 29743 2058
rect 29709 1948 29743 1986
rect 29709 1876 29743 1914
rect 29709 1804 29743 1842
rect 29709 1732 29743 1770
rect 29709 1660 29743 1698
rect 29709 1588 29743 1626
rect 29709 1516 29743 1554
rect 29709 1444 29743 1482
rect 29709 1372 29743 1410
rect 29709 1300 29743 1338
rect 29709 1228 29743 1266
rect 29709 1159 29743 1194
rect 29805 3100 29839 3135
rect 29805 3028 29839 3066
rect 29805 2956 29839 2994
rect 29805 2884 29839 2922
rect 29805 2812 29839 2850
rect 29805 2740 29839 2778
rect 29805 2668 29839 2706
rect 29805 2596 29839 2634
rect 29805 2524 29839 2562
rect 29805 2452 29839 2490
rect 29805 2380 29839 2418
rect 29805 2308 29839 2346
rect 29805 2236 29839 2274
rect 29805 2164 29839 2202
rect 29805 2092 29839 2130
rect 29805 2020 29839 2058
rect 29805 1948 29839 1986
rect 29805 1876 29839 1914
rect 29805 1804 29839 1842
rect 29805 1732 29839 1770
rect 29805 1660 29839 1698
rect 29805 1588 29839 1626
rect 29805 1516 29839 1554
rect 29805 1444 29839 1482
rect 29805 1372 29839 1410
rect 29805 1300 29839 1338
rect 29805 1228 29839 1266
rect 29805 1159 29839 1194
rect 29901 3100 29935 3135
rect 29901 3028 29935 3066
rect 29901 2956 29935 2994
rect 29901 2884 29935 2922
rect 29901 2812 29935 2850
rect 29901 2740 29935 2778
rect 29901 2668 29935 2706
rect 29901 2596 29935 2634
rect 29901 2524 29935 2562
rect 29901 2452 29935 2490
rect 29901 2380 29935 2418
rect 29901 2308 29935 2346
rect 29901 2236 29935 2274
rect 29901 2164 29935 2202
rect 29901 2092 29935 2130
rect 29901 2020 29935 2058
rect 29901 1948 29935 1986
rect 29901 1876 29935 1914
rect 29901 1804 29935 1842
rect 29901 1732 29935 1770
rect 29901 1660 29935 1698
rect 29901 1588 29935 1626
rect 29901 1516 29935 1554
rect 29901 1444 29935 1482
rect 29901 1372 29935 1410
rect 29901 1300 29935 1338
rect 29901 1228 29935 1266
rect 29901 1159 29935 1194
rect 29997 3100 30031 3135
rect 29997 3028 30031 3066
rect 29997 2956 30031 2994
rect 29997 2884 30031 2922
rect 29997 2812 30031 2850
rect 29997 2740 30031 2778
rect 29997 2668 30031 2706
rect 29997 2596 30031 2634
rect 29997 2524 30031 2562
rect 29997 2452 30031 2490
rect 29997 2380 30031 2418
rect 29997 2308 30031 2346
rect 29997 2236 30031 2274
rect 29997 2164 30031 2202
rect 29997 2092 30031 2130
rect 29997 2020 30031 2058
rect 29997 1948 30031 1986
rect 29997 1876 30031 1914
rect 29997 1804 30031 1842
rect 29997 1732 30031 1770
rect 29997 1660 30031 1698
rect 29997 1588 30031 1626
rect 29997 1516 30031 1554
rect 29997 1444 30031 1482
rect 29997 1372 30031 1410
rect 29997 1300 30031 1338
rect 29997 1228 30031 1266
rect 29997 1159 30031 1194
rect 30093 3100 30127 3135
rect 30093 3028 30127 3066
rect 30093 2956 30127 2994
rect 30093 2884 30127 2922
rect 30093 2812 30127 2850
rect 30093 2740 30127 2778
rect 30093 2668 30127 2706
rect 30093 2596 30127 2634
rect 30093 2524 30127 2562
rect 30093 2452 30127 2490
rect 30093 2380 30127 2418
rect 30093 2308 30127 2346
rect 30093 2236 30127 2274
rect 30093 2164 30127 2202
rect 30093 2092 30127 2130
rect 30093 2020 30127 2058
rect 30093 1948 30127 1986
rect 30093 1876 30127 1914
rect 30093 1804 30127 1842
rect 30093 1732 30127 1770
rect 30093 1660 30127 1698
rect 30093 1588 30127 1626
rect 30093 1516 30127 1554
rect 30093 1444 30127 1482
rect 30093 1372 30127 1410
rect 30093 1300 30127 1338
rect 30093 1228 30127 1266
rect 30093 1159 30127 1194
rect 30189 3100 30223 3135
rect 30189 3028 30223 3066
rect 30189 2956 30223 2994
rect 30189 2884 30223 2922
rect 30189 2812 30223 2850
rect 30189 2740 30223 2778
rect 30189 2668 30223 2706
rect 30189 2596 30223 2634
rect 30189 2524 30223 2562
rect 30189 2452 30223 2490
rect 30189 2380 30223 2418
rect 30189 2308 30223 2346
rect 30189 2236 30223 2274
rect 30189 2164 30223 2202
rect 30189 2092 30223 2130
rect 30189 2020 30223 2058
rect 30189 1948 30223 1986
rect 30189 1876 30223 1914
rect 30189 1804 30223 1842
rect 30189 1732 30223 1770
rect 30189 1660 30223 1698
rect 30189 1588 30223 1626
rect 30189 1516 30223 1554
rect 30189 1444 30223 1482
rect 30189 1372 30223 1410
rect 30189 1300 30223 1338
rect 30189 1228 30223 1266
rect 30189 1159 30223 1194
rect 30285 3100 30319 3135
rect 30285 3028 30319 3066
rect 30285 2956 30319 2994
rect 30285 2884 30319 2922
rect 30285 2812 30319 2850
rect 30285 2740 30319 2778
rect 30285 2668 30319 2706
rect 30285 2596 30319 2634
rect 30285 2524 30319 2562
rect 30285 2452 30319 2490
rect 30285 2380 30319 2418
rect 30285 2308 30319 2346
rect 30285 2236 30319 2274
rect 30285 2164 30319 2202
rect 30285 2092 30319 2130
rect 30285 2020 30319 2058
rect 30285 1948 30319 1986
rect 30285 1876 30319 1914
rect 30285 1804 30319 1842
rect 30285 1732 30319 1770
rect 30285 1660 30319 1698
rect 30285 1588 30319 1626
rect 30285 1516 30319 1554
rect 30285 1444 30319 1482
rect 30285 1372 30319 1410
rect 30285 1300 30319 1338
rect 30285 1228 30319 1266
rect 30285 1159 30319 1194
rect 30381 3100 30415 3135
rect 30381 3028 30415 3066
rect 30381 2956 30415 2994
rect 30381 2884 30415 2922
rect 30381 2812 30415 2850
rect 30381 2740 30415 2778
rect 30381 2668 30415 2706
rect 30381 2596 30415 2634
rect 30381 2524 30415 2562
rect 30381 2452 30415 2490
rect 30381 2380 30415 2418
rect 30381 2308 30415 2346
rect 30381 2236 30415 2274
rect 30381 2164 30415 2202
rect 30381 2092 30415 2130
rect 30381 2020 30415 2058
rect 30381 1948 30415 1986
rect 30381 1876 30415 1914
rect 30381 1804 30415 1842
rect 30381 1732 30415 1770
rect 30381 1660 30415 1698
rect 30381 1588 30415 1626
rect 30381 1516 30415 1554
rect 30381 1444 30415 1482
rect 30381 1372 30415 1410
rect 30381 1300 30415 1338
rect 30381 1228 30415 1266
rect 30381 1159 30415 1194
rect 30477 3100 30511 3135
rect 30477 3028 30511 3066
rect 30477 2956 30511 2994
rect 30477 2884 30511 2922
rect 30477 2812 30511 2850
rect 30477 2740 30511 2778
rect 30477 2668 30511 2706
rect 30477 2596 30511 2634
rect 30477 2524 30511 2562
rect 30477 2452 30511 2490
rect 30477 2380 30511 2418
rect 30477 2308 30511 2346
rect 30477 2236 30511 2274
rect 30477 2164 30511 2202
rect 30477 2092 30511 2130
rect 30477 2020 30511 2058
rect 30477 1948 30511 1986
rect 30477 1876 30511 1914
rect 30477 1804 30511 1842
rect 30477 1732 30511 1770
rect 30477 1660 30511 1698
rect 30477 1588 30511 1626
rect 30477 1516 30511 1554
rect 30477 1444 30511 1482
rect 30477 1372 30511 1410
rect 30477 1300 30511 1338
rect 30477 1228 30511 1266
rect 30477 1159 30511 1194
rect 30573 3100 30607 3135
rect 30573 3028 30607 3066
rect 30573 2956 30607 2994
rect 30573 2884 30607 2922
rect 30573 2812 30607 2850
rect 30573 2740 30607 2778
rect 30573 2668 30607 2706
rect 30573 2596 30607 2634
rect 30573 2524 30607 2562
rect 30573 2452 30607 2490
rect 30573 2380 30607 2418
rect 30573 2308 30607 2346
rect 30573 2236 30607 2274
rect 30573 2164 30607 2202
rect 30573 2092 30607 2130
rect 30573 2020 30607 2058
rect 30573 1948 30607 1986
rect 30573 1876 30607 1914
rect 30573 1804 30607 1842
rect 30573 1732 30607 1770
rect 30573 1660 30607 1698
rect 30573 1588 30607 1626
rect 30573 1516 30607 1554
rect 30573 1444 30607 1482
rect 30573 1372 30607 1410
rect 30573 1300 30607 1338
rect 30573 1228 30607 1266
rect 30573 1159 30607 1194
rect 30669 3100 30703 3135
rect 30669 3028 30703 3066
rect 30669 2956 30703 2994
rect 30669 2884 30703 2922
rect 30669 2812 30703 2850
rect 30669 2740 30703 2778
rect 30669 2668 30703 2706
rect 30669 2596 30703 2634
rect 30669 2524 30703 2562
rect 30669 2452 30703 2490
rect 30669 2380 30703 2418
rect 30669 2308 30703 2346
rect 30669 2236 30703 2274
rect 30669 2164 30703 2202
rect 30669 2092 30703 2130
rect 30669 2020 30703 2058
rect 30669 1948 30703 1986
rect 30669 1876 30703 1914
rect 30669 1804 30703 1842
rect 30669 1732 30703 1770
rect 30669 1660 30703 1698
rect 30669 1588 30703 1626
rect 30669 1516 30703 1554
rect 30669 1444 30703 1482
rect 30669 1372 30703 1410
rect 30669 1300 30703 1338
rect 30669 1228 30703 1266
rect 30669 1159 30703 1194
rect 30765 3100 30799 3135
rect 30765 3028 30799 3066
rect 30765 2956 30799 2994
rect 30765 2884 30799 2922
rect 30765 2812 30799 2850
rect 30765 2740 30799 2778
rect 30765 2668 30799 2706
rect 30765 2596 30799 2634
rect 30765 2524 30799 2562
rect 30765 2452 30799 2490
rect 30765 2380 30799 2418
rect 30765 2308 30799 2346
rect 30765 2236 30799 2274
rect 30765 2164 30799 2202
rect 30765 2092 30799 2130
rect 30765 2020 30799 2058
rect 30765 1948 30799 1986
rect 30765 1876 30799 1914
rect 30765 1804 30799 1842
rect 30765 1732 30799 1770
rect 30765 1660 30799 1698
rect 30765 1588 30799 1626
rect 30765 1516 30799 1554
rect 30765 1444 30799 1482
rect 30765 1372 30799 1410
rect 30765 1300 30799 1338
rect 30765 1228 30799 1266
rect 30765 1159 30799 1194
rect 30861 3100 30895 3135
rect 30861 3028 30895 3066
rect 30861 2956 30895 2994
rect 30861 2884 30895 2922
rect 30861 2812 30895 2850
rect 30861 2740 30895 2778
rect 30861 2668 30895 2706
rect 30861 2596 30895 2634
rect 30861 2524 30895 2562
rect 30861 2452 30895 2490
rect 30861 2380 30895 2418
rect 30861 2308 30895 2346
rect 30861 2236 30895 2274
rect 30861 2164 30895 2202
rect 30861 2092 30895 2130
rect 30861 2020 30895 2058
rect 30861 1948 30895 1986
rect 30861 1876 30895 1914
rect 30861 1804 30895 1842
rect 30861 1732 30895 1770
rect 30861 1660 30895 1698
rect 30861 1588 30895 1626
rect 30861 1516 30895 1554
rect 30861 1444 30895 1482
rect 30861 1372 30895 1410
rect 30861 1300 30895 1338
rect 30861 1228 30895 1266
rect 30861 1159 30895 1194
rect 30957 3100 30991 3135
rect 30957 3028 30991 3066
rect 30957 2956 30991 2994
rect 30957 2884 30991 2922
rect 30957 2812 30991 2850
rect 30957 2740 30991 2778
rect 30957 2668 30991 2706
rect 30957 2596 30991 2634
rect 30957 2524 30991 2562
rect 30957 2452 30991 2490
rect 30957 2380 30991 2418
rect 30957 2308 30991 2346
rect 30957 2236 30991 2274
rect 30957 2164 30991 2202
rect 30957 2092 30991 2130
rect 30957 2020 30991 2058
rect 30957 1948 30991 1986
rect 30957 1876 30991 1914
rect 30957 1804 30991 1842
rect 30957 1732 30991 1770
rect 30957 1660 30991 1698
rect 30957 1588 30991 1626
rect 30957 1516 30991 1554
rect 30957 1444 30991 1482
rect 30957 1372 30991 1410
rect 30957 1300 30991 1338
rect 30957 1228 30991 1266
rect 30957 1159 30991 1194
rect 31053 3100 31087 3135
rect 31053 3028 31087 3066
rect 31053 2956 31087 2994
rect 31053 2884 31087 2922
rect 31053 2812 31087 2850
rect 31053 2740 31087 2778
rect 31053 2668 31087 2706
rect 31053 2596 31087 2634
rect 31053 2524 31087 2562
rect 31053 2452 31087 2490
rect 31053 2380 31087 2418
rect 31053 2308 31087 2346
rect 31053 2236 31087 2274
rect 31053 2164 31087 2202
rect 31053 2092 31087 2130
rect 31053 2020 31087 2058
rect 31053 1948 31087 1986
rect 31053 1876 31087 1914
rect 31053 1804 31087 1842
rect 31053 1732 31087 1770
rect 31053 1660 31087 1698
rect 31053 1588 31087 1626
rect 31053 1516 31087 1554
rect 31053 1444 31087 1482
rect 31053 1372 31087 1410
rect 31053 1300 31087 1338
rect 31053 1228 31087 1266
rect 31053 1159 31087 1194
rect 31149 3100 31183 3135
rect 31149 3028 31183 3066
rect 31149 2956 31183 2994
rect 31149 2884 31183 2922
rect 31149 2812 31183 2850
rect 31149 2740 31183 2778
rect 31149 2668 31183 2706
rect 31149 2596 31183 2634
rect 31149 2524 31183 2562
rect 31149 2452 31183 2490
rect 31149 2380 31183 2418
rect 31149 2308 31183 2346
rect 31149 2236 31183 2274
rect 31149 2164 31183 2202
rect 31149 2092 31183 2130
rect 31149 2020 31183 2058
rect 31149 1948 31183 1986
rect 31149 1876 31183 1914
rect 31149 1804 31183 1842
rect 31149 1732 31183 1770
rect 31149 1660 31183 1698
rect 31149 1588 31183 1626
rect 31149 1516 31183 1554
rect 31149 1444 31183 1482
rect 31149 1372 31183 1410
rect 31149 1300 31183 1338
rect 31149 1228 31183 1266
rect 31149 1159 31183 1194
rect 31245 3100 31279 3135
rect 31245 3028 31279 3066
rect 31245 2956 31279 2994
rect 31245 2884 31279 2922
rect 31245 2812 31279 2850
rect 31245 2740 31279 2778
rect 31245 2668 31279 2706
rect 31245 2596 31279 2634
rect 31245 2524 31279 2562
rect 31245 2452 31279 2490
rect 31245 2380 31279 2418
rect 31245 2308 31279 2346
rect 31245 2236 31279 2274
rect 31245 2164 31279 2202
rect 31245 2092 31279 2130
rect 31245 2020 31279 2058
rect 31245 1948 31279 1986
rect 31245 1876 31279 1914
rect 31245 1804 31279 1842
rect 31245 1732 31279 1770
rect 31245 1660 31279 1698
rect 31245 1588 31279 1626
rect 31245 1516 31279 1554
rect 31245 1444 31279 1482
rect 31245 1372 31279 1410
rect 31245 1300 31279 1338
rect 31245 1228 31279 1266
rect 31245 1159 31279 1194
rect 31341 3100 31375 3135
rect 31341 3028 31375 3066
rect 31341 2956 31375 2994
rect 31341 2884 31375 2922
rect 31341 2812 31375 2850
rect 31341 2740 31375 2778
rect 31341 2668 31375 2706
rect 31341 2596 31375 2634
rect 31341 2524 31375 2562
rect 31341 2452 31375 2490
rect 31341 2380 31375 2418
rect 31341 2308 31375 2346
rect 31341 2236 31375 2274
rect 31341 2164 31375 2202
rect 31341 2092 31375 2130
rect 31341 2020 31375 2058
rect 31341 1948 31375 1986
rect 31341 1876 31375 1914
rect 31341 1804 31375 1842
rect 31341 1732 31375 1770
rect 31341 1660 31375 1698
rect 31341 1588 31375 1626
rect 31341 1516 31375 1554
rect 31341 1444 31375 1482
rect 31341 1372 31375 1410
rect 31341 1300 31375 1338
rect 31341 1228 31375 1266
rect 31341 1159 31375 1194
rect 31437 3100 31471 3135
rect 31437 3028 31471 3066
rect 31437 2956 31471 2994
rect 31437 2884 31471 2922
rect 31437 2812 31471 2850
rect 31437 2740 31471 2778
rect 31437 2668 31471 2706
rect 31437 2596 31471 2634
rect 31437 2524 31471 2562
rect 31437 2452 31471 2490
rect 31437 2380 31471 2418
rect 31437 2308 31471 2346
rect 31437 2236 31471 2274
rect 31437 2164 31471 2202
rect 31437 2092 31471 2130
rect 31437 2020 31471 2058
rect 31437 1948 31471 1986
rect 31437 1876 31471 1914
rect 31437 1804 31471 1842
rect 31437 1732 31471 1770
rect 31437 1660 31471 1698
rect 31437 1588 31471 1626
rect 31437 1516 31471 1554
rect 31437 1444 31471 1482
rect 31437 1372 31471 1410
rect 31437 1300 31471 1338
rect 31437 1228 31471 1266
rect 31437 1159 31471 1194
rect 31533 3100 31567 3135
rect 31533 3028 31567 3066
rect 31533 2956 31567 2994
rect 31533 2884 31567 2922
rect 31533 2812 31567 2850
rect 31533 2740 31567 2778
rect 31533 2668 31567 2706
rect 31533 2596 31567 2634
rect 31533 2524 31567 2562
rect 31533 2452 31567 2490
rect 31533 2380 31567 2418
rect 31533 2308 31567 2346
rect 31533 2236 31567 2274
rect 31533 2164 31567 2202
rect 31533 2092 31567 2130
rect 31533 2020 31567 2058
rect 31533 1948 31567 1986
rect 31533 1876 31567 1914
rect 31533 1804 31567 1842
rect 31533 1732 31567 1770
rect 31533 1660 31567 1698
rect 31533 1588 31567 1626
rect 31533 1516 31567 1554
rect 31533 1444 31567 1482
rect 31533 1372 31567 1410
rect 31533 1300 31567 1338
rect 31533 1228 31567 1266
rect 31533 1159 31567 1194
rect 31629 3100 31663 3135
rect 31629 3028 31663 3066
rect 31629 2956 31663 2994
rect 31629 2884 31663 2922
rect 31629 2812 31663 2850
rect 31629 2740 31663 2778
rect 31629 2668 31663 2706
rect 31629 2596 31663 2634
rect 31629 2524 31663 2562
rect 31629 2452 31663 2490
rect 31629 2380 31663 2418
rect 31629 2308 31663 2346
rect 31629 2236 31663 2274
rect 31629 2164 31663 2202
rect 31629 2092 31663 2130
rect 31629 2020 31663 2058
rect 31629 1948 31663 1986
rect 31629 1876 31663 1914
rect 31629 1804 31663 1842
rect 31629 1732 31663 1770
rect 31629 1660 31663 1698
rect 31629 1588 31663 1626
rect 31629 1516 31663 1554
rect 31629 1444 31663 1482
rect 31629 1372 31663 1410
rect 31629 1300 31663 1338
rect 31629 1228 31663 1266
rect 31629 1159 31663 1194
rect 31725 3100 31759 3135
rect 31725 3028 31759 3066
rect 31725 2956 31759 2994
rect 31725 2884 31759 2922
rect 31725 2812 31759 2850
rect 31725 2740 31759 2778
rect 31725 2668 31759 2706
rect 31725 2596 31759 2634
rect 31725 2524 31759 2562
rect 31725 2452 31759 2490
rect 31725 2380 31759 2418
rect 31725 2308 31759 2346
rect 31725 2236 31759 2274
rect 31725 2164 31759 2202
rect 31725 2092 31759 2130
rect 31725 2020 31759 2058
rect 31725 1948 31759 1986
rect 31725 1876 31759 1914
rect 31725 1804 31759 1842
rect 31725 1732 31759 1770
rect 31725 1660 31759 1698
rect 31725 1588 31759 1626
rect 31725 1516 31759 1554
rect 31725 1444 31759 1482
rect 31725 1372 31759 1410
rect 31725 1300 31759 1338
rect 31725 1228 31759 1266
rect 31725 1159 31759 1194
rect 31821 3100 31855 3135
rect 31821 3028 31855 3066
rect 31821 2956 31855 2994
rect 31821 2884 31855 2922
rect 31821 2812 31855 2850
rect 31821 2740 31855 2778
rect 31821 2668 31855 2706
rect 31821 2596 31855 2634
rect 31821 2524 31855 2562
rect 31821 2452 31855 2490
rect 31821 2380 31855 2418
rect 31821 2308 31855 2346
rect 31821 2236 31855 2274
rect 31821 2164 31855 2202
rect 31821 2092 31855 2130
rect 31821 2020 31855 2058
rect 31821 1948 31855 1986
rect 31821 1876 31855 1914
rect 31821 1804 31855 1842
rect 31821 1732 31855 1770
rect 31821 1660 31855 1698
rect 31821 1588 31855 1626
rect 31821 1516 31855 1554
rect 31821 1444 31855 1482
rect 31821 1372 31855 1410
rect 31821 1300 31855 1338
rect 31821 1228 31855 1266
rect 31821 1159 31855 1194
rect 31917 3100 31951 3135
rect 31917 3028 31951 3066
rect 31917 2956 31951 2994
rect 31917 2884 31951 2922
rect 31917 2812 31951 2850
rect 31917 2740 31951 2778
rect 31917 2668 31951 2706
rect 31917 2596 31951 2634
rect 31917 2524 31951 2562
rect 31917 2452 31951 2490
rect 31917 2380 31951 2418
rect 31917 2308 31951 2346
rect 31917 2236 31951 2274
rect 31917 2164 31951 2202
rect 31917 2092 31951 2130
rect 31917 2020 31951 2058
rect 31917 1948 31951 1986
rect 31917 1876 31951 1914
rect 31917 1804 31951 1842
rect 31917 1732 31951 1770
rect 31917 1660 31951 1698
rect 31917 1588 31951 1626
rect 31917 1516 31951 1554
rect 31917 1444 31951 1482
rect 31917 1372 31951 1410
rect 31917 1300 31951 1338
rect 31917 1228 31951 1266
rect 31917 1159 31951 1194
rect 32013 3100 32047 3135
rect 32013 3028 32047 3066
rect 32013 2956 32047 2994
rect 32013 2884 32047 2922
rect 32013 2812 32047 2850
rect 32013 2740 32047 2778
rect 32013 2668 32047 2706
rect 32013 2596 32047 2634
rect 32013 2524 32047 2562
rect 32013 2452 32047 2490
rect 32013 2380 32047 2418
rect 32013 2308 32047 2346
rect 32013 2236 32047 2274
rect 32013 2164 32047 2202
rect 32013 2092 32047 2130
rect 32013 2020 32047 2058
rect 32013 1948 32047 1986
rect 32013 1876 32047 1914
rect 32013 1804 32047 1842
rect 32013 1732 32047 1770
rect 32013 1660 32047 1698
rect 32013 1588 32047 1626
rect 32013 1516 32047 1554
rect 32013 1444 32047 1482
rect 32013 1372 32047 1410
rect 32013 1300 32047 1338
rect 32013 1228 32047 1266
rect 32013 1159 32047 1194
rect 32109 3100 32143 3135
rect 32109 3028 32143 3066
rect 32109 2956 32143 2994
rect 32109 2884 32143 2922
rect 32109 2812 32143 2850
rect 32109 2740 32143 2778
rect 32109 2668 32143 2706
rect 32109 2596 32143 2634
rect 32109 2524 32143 2562
rect 32109 2452 32143 2490
rect 32109 2380 32143 2418
rect 32109 2308 32143 2346
rect 32109 2236 32143 2274
rect 32109 2164 32143 2202
rect 32109 2092 32143 2130
rect 32109 2020 32143 2058
rect 32109 1948 32143 1986
rect 32109 1876 32143 1914
rect 32109 1804 32143 1842
rect 32109 1732 32143 1770
rect 32109 1660 32143 1698
rect 32109 1588 32143 1626
rect 32109 1516 32143 1554
rect 32109 1444 32143 1482
rect 32109 1372 32143 1410
rect 32109 1300 32143 1338
rect 32109 1228 32143 1266
rect 32109 1159 32143 1194
rect 32205 3100 32239 3135
rect 32205 3028 32239 3066
rect 32205 2956 32239 2994
rect 32205 2884 32239 2922
rect 32205 2812 32239 2850
rect 32205 2740 32239 2778
rect 32205 2668 32239 2706
rect 32205 2596 32239 2634
rect 32205 2524 32239 2562
rect 32205 2452 32239 2490
rect 32205 2380 32239 2418
rect 32205 2308 32239 2346
rect 32205 2236 32239 2274
rect 32205 2164 32239 2202
rect 32205 2092 32239 2130
rect 32205 2020 32239 2058
rect 32205 1948 32239 1986
rect 32205 1876 32239 1914
rect 32205 1804 32239 1842
rect 32205 1732 32239 1770
rect 32205 1660 32239 1698
rect 32205 1588 32239 1626
rect 32205 1516 32239 1554
rect 32205 1444 32239 1482
rect 32205 1372 32239 1410
rect 32205 1300 32239 1338
rect 32205 1228 32239 1266
rect 32205 1159 32239 1194
rect 32301 3100 32335 3135
rect 32301 3028 32335 3066
rect 32301 2956 32335 2994
rect 32301 2884 32335 2922
rect 32301 2812 32335 2850
rect 32301 2740 32335 2778
rect 32301 2668 32335 2706
rect 32301 2596 32335 2634
rect 32301 2524 32335 2562
rect 32301 2452 32335 2490
rect 32301 2380 32335 2418
rect 32301 2308 32335 2346
rect 32301 2236 32335 2274
rect 32301 2164 32335 2202
rect 32301 2092 32335 2130
rect 32301 2020 32335 2058
rect 32301 1948 32335 1986
rect 32301 1876 32335 1914
rect 32301 1804 32335 1842
rect 32301 1732 32335 1770
rect 32301 1660 32335 1698
rect 32301 1588 32335 1626
rect 32301 1516 32335 1554
rect 32301 1444 32335 1482
rect 32301 1372 32335 1410
rect 32301 1300 32335 1338
rect 32301 1228 32335 1266
rect 32301 1159 32335 1194
rect 32397 3100 32431 3135
rect 32397 3028 32431 3066
rect 32397 2956 32431 2994
rect 32397 2884 32431 2922
rect 32397 2812 32431 2850
rect 32397 2740 32431 2778
rect 32397 2668 32431 2706
rect 32397 2596 32431 2634
rect 32397 2524 32431 2562
rect 32397 2452 32431 2490
rect 32397 2380 32431 2418
rect 32397 2308 32431 2346
rect 32397 2236 32431 2274
rect 32397 2164 32431 2202
rect 32397 2092 32431 2130
rect 32397 2020 32431 2058
rect 32397 1948 32431 1986
rect 32397 1876 32431 1914
rect 32397 1804 32431 1842
rect 32397 1732 32431 1770
rect 32397 1660 32431 1698
rect 32397 1588 32431 1626
rect 32397 1516 32431 1554
rect 32397 1444 32431 1482
rect 32397 1372 32431 1410
rect 32397 1300 32431 1338
rect 32397 1228 32431 1266
rect 32397 1159 32431 1194
rect 32493 3100 32527 3135
rect 32493 3028 32527 3066
rect 32493 2956 32527 2994
rect 32493 2884 32527 2922
rect 32493 2812 32527 2850
rect 32493 2740 32527 2778
rect 32493 2668 32527 2706
rect 32493 2596 32527 2634
rect 32493 2524 32527 2562
rect 32493 2452 32527 2490
rect 32493 2380 32527 2418
rect 32493 2308 32527 2346
rect 32493 2236 32527 2274
rect 32493 2164 32527 2202
rect 32493 2092 32527 2130
rect 32493 2020 32527 2058
rect 32493 1948 32527 1986
rect 32493 1876 32527 1914
rect 32493 1804 32527 1842
rect 32493 1732 32527 1770
rect 32493 1660 32527 1698
rect 32493 1588 32527 1626
rect 32493 1516 32527 1554
rect 32493 1444 32527 1482
rect 32493 1372 32527 1410
rect 32493 1300 32527 1338
rect 32493 1228 32527 1266
rect 32493 1159 32527 1194
rect 32589 3100 32623 3135
rect 32589 3028 32623 3066
rect 32589 2956 32623 2994
rect 32589 2884 32623 2922
rect 32589 2812 32623 2850
rect 32589 2740 32623 2778
rect 32589 2668 32623 2706
rect 32589 2596 32623 2634
rect 32589 2524 32623 2562
rect 32589 2452 32623 2490
rect 32589 2380 32623 2418
rect 32589 2308 32623 2346
rect 32589 2236 32623 2274
rect 32589 2164 32623 2202
rect 32589 2092 32623 2130
rect 32589 2020 32623 2058
rect 32589 1948 32623 1986
rect 32589 1876 32623 1914
rect 32589 1804 32623 1842
rect 32589 1732 32623 1770
rect 32589 1660 32623 1698
rect 32589 1588 32623 1626
rect 32589 1516 32623 1554
rect 32589 1444 32623 1482
rect 32589 1372 32623 1410
rect 32589 1300 32623 1338
rect 32589 1228 32623 1266
rect 32589 1159 32623 1194
rect 32685 3100 32719 3135
rect 32685 3028 32719 3066
rect 32685 2956 32719 2994
rect 32685 2884 32719 2922
rect 32685 2812 32719 2850
rect 32685 2740 32719 2778
rect 32685 2668 32719 2706
rect 32685 2596 32719 2634
rect 32685 2524 32719 2562
rect 32685 2452 32719 2490
rect 32685 2380 32719 2418
rect 32685 2308 32719 2346
rect 32685 2236 32719 2274
rect 32685 2164 32719 2202
rect 32685 2092 32719 2130
rect 32685 2020 32719 2058
rect 32685 1948 32719 1986
rect 32685 1876 32719 1914
rect 32685 1804 32719 1842
rect 32685 1732 32719 1770
rect 32685 1660 32719 1698
rect 32685 1588 32719 1626
rect 32685 1516 32719 1554
rect 32685 1444 32719 1482
rect 32685 1372 32719 1410
rect 32685 1300 32719 1338
rect 32685 1228 32719 1266
rect 32685 1159 32719 1194
rect 32781 3100 32815 3135
rect 32781 3028 32815 3066
rect 32781 2956 32815 2994
rect 32781 2884 32815 2922
rect 32781 2812 32815 2850
rect 32781 2740 32815 2778
rect 32781 2668 32815 2706
rect 32781 2596 32815 2634
rect 32781 2524 32815 2562
rect 32781 2452 32815 2490
rect 32781 2380 32815 2418
rect 32781 2308 32815 2346
rect 32781 2236 32815 2274
rect 32781 2164 32815 2202
rect 32781 2092 32815 2130
rect 32781 2020 32815 2058
rect 32781 1948 32815 1986
rect 32781 1876 32815 1914
rect 32781 1804 32815 1842
rect 32781 1732 32815 1770
rect 32781 1660 32815 1698
rect 32781 1588 32815 1626
rect 32781 1516 32815 1554
rect 32781 1444 32815 1482
rect 32781 1372 32815 1410
rect 32781 1300 32815 1338
rect 32781 1228 32815 1266
rect 32781 1159 32815 1194
rect 32877 3100 32911 3135
rect 32877 3028 32911 3066
rect 32877 2956 32911 2994
rect 32877 2884 32911 2922
rect 32877 2812 32911 2850
rect 32877 2740 32911 2778
rect 32877 2668 32911 2706
rect 32877 2596 32911 2634
rect 32877 2524 32911 2562
rect 32877 2452 32911 2490
rect 32877 2380 32911 2418
rect 32877 2308 32911 2346
rect 32877 2236 32911 2274
rect 32877 2164 32911 2202
rect 32877 2092 32911 2130
rect 32877 2020 32911 2058
rect 32877 1948 32911 1986
rect 32877 1876 32911 1914
rect 32877 1804 32911 1842
rect 32877 1732 32911 1770
rect 32877 1660 32911 1698
rect 32877 1588 32911 1626
rect 32877 1516 32911 1554
rect 32877 1444 32911 1482
rect 32877 1372 32911 1410
rect 32877 1300 32911 1338
rect 32877 1228 32911 1266
rect 32877 1159 32911 1194
rect 32973 3100 33007 3135
rect 32973 3028 33007 3066
rect 32973 2956 33007 2994
rect 32973 2884 33007 2922
rect 32973 2812 33007 2850
rect 32973 2740 33007 2778
rect 32973 2668 33007 2706
rect 32973 2596 33007 2634
rect 32973 2524 33007 2562
rect 32973 2452 33007 2490
rect 32973 2380 33007 2418
rect 32973 2308 33007 2346
rect 32973 2236 33007 2274
rect 32973 2164 33007 2202
rect 32973 2092 33007 2130
rect 32973 2020 33007 2058
rect 32973 1948 33007 1986
rect 32973 1876 33007 1914
rect 32973 1804 33007 1842
rect 32973 1732 33007 1770
rect 32973 1660 33007 1698
rect 32973 1588 33007 1626
rect 32973 1516 33007 1554
rect 32973 1444 33007 1482
rect 32973 1372 33007 1410
rect 32973 1300 33007 1338
rect 32973 1228 33007 1266
rect 32973 1159 33007 1194
rect 33069 3100 33103 3135
rect 33069 3028 33103 3066
rect 33069 2956 33103 2994
rect 33069 2884 33103 2922
rect 33069 2812 33103 2850
rect 33069 2740 33103 2778
rect 33069 2668 33103 2706
rect 33069 2596 33103 2634
rect 33069 2524 33103 2562
rect 33069 2452 33103 2490
rect 33069 2380 33103 2418
rect 33069 2308 33103 2346
rect 33069 2236 33103 2274
rect 33069 2164 33103 2202
rect 33069 2092 33103 2130
rect 33069 2020 33103 2058
rect 33069 1948 33103 1986
rect 33069 1876 33103 1914
rect 33069 1804 33103 1842
rect 33069 1732 33103 1770
rect 33069 1660 33103 1698
rect 33069 1588 33103 1626
rect 33069 1516 33103 1554
rect 33069 1444 33103 1482
rect 33069 1372 33103 1410
rect 33069 1300 33103 1338
rect 33069 1228 33103 1266
rect 33069 1159 33103 1194
rect 33165 3100 33199 3135
rect 33165 3028 33199 3066
rect 33165 2956 33199 2994
rect 33165 2884 33199 2922
rect 33165 2812 33199 2850
rect 33165 2740 33199 2778
rect 33165 2668 33199 2706
rect 33165 2596 33199 2634
rect 33165 2524 33199 2562
rect 33165 2452 33199 2490
rect 33165 2380 33199 2418
rect 33165 2308 33199 2346
rect 33165 2236 33199 2274
rect 33165 2164 33199 2202
rect 33165 2092 33199 2130
rect 33165 2020 33199 2058
rect 33165 1948 33199 1986
rect 33165 1876 33199 1914
rect 33165 1804 33199 1842
rect 33165 1732 33199 1770
rect 33165 1660 33199 1698
rect 33165 1588 33199 1626
rect 33165 1516 33199 1554
rect 33165 1444 33199 1482
rect 33165 1372 33199 1410
rect 33165 1300 33199 1338
rect 33165 1228 33199 1266
rect 33165 1159 33199 1194
rect 33261 3100 33295 3135
rect 33261 3028 33295 3066
rect 33261 2956 33295 2994
rect 33261 2884 33295 2922
rect 33261 2812 33295 2850
rect 33261 2740 33295 2778
rect 33261 2668 33295 2706
rect 33261 2596 33295 2634
rect 33261 2524 33295 2562
rect 33261 2452 33295 2490
rect 33261 2380 33295 2418
rect 33261 2308 33295 2346
rect 33261 2236 33295 2274
rect 33261 2164 33295 2202
rect 33261 2092 33295 2130
rect 33261 2020 33295 2058
rect 33261 1948 33295 1986
rect 33261 1876 33295 1914
rect 33261 1804 33295 1842
rect 33261 1732 33295 1770
rect 33261 1660 33295 1698
rect 33261 1588 33295 1626
rect 33261 1516 33295 1554
rect 33261 1444 33295 1482
rect 33261 1372 33295 1410
rect 33261 1300 33295 1338
rect 33261 1228 33295 1266
rect 33261 1159 33295 1194
rect 33357 3100 33391 3135
rect 33357 3028 33391 3066
rect 33357 2956 33391 2994
rect 33357 2884 33391 2922
rect 33357 2812 33391 2850
rect 33357 2740 33391 2778
rect 33357 2668 33391 2706
rect 33357 2596 33391 2634
rect 33357 2524 33391 2562
rect 33357 2452 33391 2490
rect 33357 2380 33391 2418
rect 33357 2308 33391 2346
rect 33357 2236 33391 2274
rect 33357 2164 33391 2202
rect 33357 2092 33391 2130
rect 33357 2020 33391 2058
rect 33357 1948 33391 1986
rect 33357 1876 33391 1914
rect 33357 1804 33391 1842
rect 33357 1732 33391 1770
rect 33357 1660 33391 1698
rect 33357 1588 33391 1626
rect 33357 1516 33391 1554
rect 33357 1444 33391 1482
rect 33357 1372 33391 1410
rect 33357 1300 33391 1338
rect 33357 1228 33391 1266
rect 33357 1159 33391 1194
rect 33453 3100 33487 3135
rect 33453 3028 33487 3066
rect 33453 2956 33487 2994
rect 33453 2884 33487 2922
rect 33453 2812 33487 2850
rect 33453 2740 33487 2778
rect 33453 2668 33487 2706
rect 33453 2596 33487 2634
rect 33453 2524 33487 2562
rect 33453 2452 33487 2490
rect 33453 2380 33487 2418
rect 33453 2308 33487 2346
rect 33453 2236 33487 2274
rect 33453 2164 33487 2202
rect 33453 2092 33487 2130
rect 33453 2020 33487 2058
rect 33453 1948 33487 1986
rect 33453 1876 33487 1914
rect 33453 1804 33487 1842
rect 33453 1732 33487 1770
rect 33453 1660 33487 1698
rect 33453 1588 33487 1626
rect 33453 1516 33487 1554
rect 33453 1444 33487 1482
rect 33453 1372 33487 1410
rect 33453 1300 33487 1338
rect 33453 1228 33487 1266
rect 33453 1159 33487 1194
rect 33549 3100 33583 3135
rect 33549 3028 33583 3066
rect 33549 2956 33583 2994
rect 33549 2884 33583 2922
rect 33549 2812 33583 2850
rect 33549 2740 33583 2778
rect 33549 2668 33583 2706
rect 33549 2596 33583 2634
rect 33549 2524 33583 2562
rect 33549 2452 33583 2490
rect 33549 2380 33583 2418
rect 33549 2308 33583 2346
rect 33549 2236 33583 2274
rect 33549 2164 33583 2202
rect 33549 2092 33583 2130
rect 33549 2020 33583 2058
rect 33549 1948 33583 1986
rect 33549 1876 33583 1914
rect 33549 1804 33583 1842
rect 33549 1732 33583 1770
rect 33549 1660 33583 1698
rect 33549 1588 33583 1626
rect 33549 1516 33583 1554
rect 33549 1444 33583 1482
rect 33549 1372 33583 1410
rect 33549 1300 33583 1338
rect 33549 1228 33583 1266
rect 33549 1159 33583 1194
rect 33645 3100 33679 3135
rect 33645 3028 33679 3066
rect 33645 2956 33679 2994
rect 33645 2884 33679 2922
rect 33645 2812 33679 2850
rect 33645 2740 33679 2778
rect 33645 2668 33679 2706
rect 33645 2596 33679 2634
rect 33645 2524 33679 2562
rect 33645 2452 33679 2490
rect 33645 2380 33679 2418
rect 33645 2308 33679 2346
rect 33645 2236 33679 2274
rect 33645 2164 33679 2202
rect 33645 2092 33679 2130
rect 33645 2020 33679 2058
rect 33645 1948 33679 1986
rect 33645 1876 33679 1914
rect 33645 1804 33679 1842
rect 33645 1732 33679 1770
rect 33645 1660 33679 1698
rect 33645 1588 33679 1626
rect 33645 1516 33679 1554
rect 33645 1444 33679 1482
rect 33645 1372 33679 1410
rect 33645 1300 33679 1338
rect 33645 1228 33679 1266
rect 33645 1159 33679 1194
rect 33741 3100 33775 3135
rect 33741 3028 33775 3066
rect 33741 2956 33775 2994
rect 33741 2884 33775 2922
rect 33741 2812 33775 2850
rect 33741 2740 33775 2778
rect 33741 2668 33775 2706
rect 33741 2596 33775 2634
rect 33741 2524 33775 2562
rect 33741 2452 33775 2490
rect 33741 2380 33775 2418
rect 33741 2308 33775 2346
rect 33741 2236 33775 2274
rect 33741 2164 33775 2202
rect 33741 2092 33775 2130
rect 33741 2020 33775 2058
rect 33741 1948 33775 1986
rect 33741 1876 33775 1914
rect 33741 1804 33775 1842
rect 33741 1732 33775 1770
rect 33741 1660 33775 1698
rect 33741 1588 33775 1626
rect 33741 1516 33775 1554
rect 33741 1444 33775 1482
rect 33741 1372 33775 1410
rect 33741 1300 33775 1338
rect 33741 1228 33775 1266
rect 33741 1159 33775 1194
rect 33837 3100 33871 3135
rect 33837 3028 33871 3066
rect 33837 2956 33871 2994
rect 33837 2884 33871 2922
rect 33837 2812 33871 2850
rect 33837 2740 33871 2778
rect 33837 2668 33871 2706
rect 33837 2596 33871 2634
rect 33837 2524 33871 2562
rect 33837 2452 33871 2490
rect 33837 2380 33871 2418
rect 33837 2308 33871 2346
rect 33837 2236 33871 2274
rect 33837 2164 33871 2202
rect 33837 2092 33871 2130
rect 33837 2020 33871 2058
rect 33837 1948 33871 1986
rect 33837 1876 33871 1914
rect 33837 1804 33871 1842
rect 33837 1732 33871 1770
rect 33837 1660 33871 1698
rect 33837 1588 33871 1626
rect 33837 1516 33871 1554
rect 33837 1444 33871 1482
rect 33837 1372 33871 1410
rect 33837 1300 33871 1338
rect 33837 1228 33871 1266
rect 33837 1159 33871 1194
rect 33933 3100 33967 3135
rect 33933 3028 33967 3066
rect 33933 2956 33967 2994
rect 33933 2884 33967 2922
rect 33933 2812 33967 2850
rect 33933 2740 33967 2778
rect 33933 2668 33967 2706
rect 33933 2596 33967 2634
rect 33933 2524 33967 2562
rect 33933 2452 33967 2490
rect 33933 2380 33967 2418
rect 33933 2308 33967 2346
rect 33933 2236 33967 2274
rect 33933 2164 33967 2202
rect 33933 2092 33967 2130
rect 33933 2020 33967 2058
rect 33933 1948 33967 1986
rect 33933 1876 33967 1914
rect 33933 1804 33967 1842
rect 33933 1732 33967 1770
rect 33933 1660 33967 1698
rect 33933 1588 33967 1626
rect 33933 1516 33967 1554
rect 33933 1444 33967 1482
rect 33933 1372 33967 1410
rect 33933 1300 33967 1338
rect 33933 1228 33967 1266
rect 33933 1159 33967 1194
rect 34029 3100 34063 3135
rect 34029 3028 34063 3066
rect 34029 2956 34063 2994
rect 34029 2884 34063 2922
rect 34029 2812 34063 2850
rect 34029 2740 34063 2778
rect 34029 2668 34063 2706
rect 34029 2596 34063 2634
rect 34029 2524 34063 2562
rect 34029 2452 34063 2490
rect 34029 2380 34063 2418
rect 34029 2308 34063 2346
rect 34029 2236 34063 2274
rect 34029 2164 34063 2202
rect 34029 2092 34063 2130
rect 34029 2020 34063 2058
rect 34029 1948 34063 1986
rect 34029 1876 34063 1914
rect 34029 1804 34063 1842
rect 34029 1732 34063 1770
rect 34029 1660 34063 1698
rect 34029 1588 34063 1626
rect 34029 1516 34063 1554
rect 34029 1444 34063 1482
rect 34029 1372 34063 1410
rect 34029 1300 34063 1338
rect 34029 1228 34063 1266
rect 34029 1159 34063 1194
rect 34125 3100 34159 3135
rect 34125 3028 34159 3066
rect 34125 2956 34159 2994
rect 34125 2884 34159 2922
rect 34125 2812 34159 2850
rect 34125 2740 34159 2778
rect 34125 2668 34159 2706
rect 34125 2596 34159 2634
rect 34125 2524 34159 2562
rect 34125 2452 34159 2490
rect 34125 2380 34159 2418
rect 34125 2308 34159 2346
rect 34125 2236 34159 2274
rect 34125 2164 34159 2202
rect 34125 2092 34159 2130
rect 34125 2020 34159 2058
rect 34125 1948 34159 1986
rect 34125 1876 34159 1914
rect 34125 1804 34159 1842
rect 34125 1732 34159 1770
rect 34125 1660 34159 1698
rect 34125 1588 34159 1626
rect 34125 1516 34159 1554
rect 34125 1444 34159 1482
rect 34125 1372 34159 1410
rect 34125 1300 34159 1338
rect 34125 1228 34159 1266
rect 34125 1159 34159 1194
rect 34221 3100 34255 3135
rect 34221 3028 34255 3066
rect 34221 2956 34255 2994
rect 34221 2884 34255 2922
rect 34221 2812 34255 2850
rect 34221 2740 34255 2778
rect 34221 2668 34255 2706
rect 34221 2596 34255 2634
rect 34221 2524 34255 2562
rect 34221 2452 34255 2490
rect 34221 2380 34255 2418
rect 34221 2308 34255 2346
rect 34221 2236 34255 2274
rect 34221 2164 34255 2202
rect 34221 2092 34255 2130
rect 34221 2020 34255 2058
rect 34221 1948 34255 1986
rect 34221 1876 34255 1914
rect 34221 1804 34255 1842
rect 34221 1732 34255 1770
rect 34221 1660 34255 1698
rect 34221 1588 34255 1626
rect 34221 1516 34255 1554
rect 34221 1444 34255 1482
rect 34221 1372 34255 1410
rect 34221 1300 34255 1338
rect 34221 1228 34255 1266
rect 34221 1159 34255 1194
rect 34317 3100 34351 3135
rect 34317 3028 34351 3066
rect 34317 2956 34351 2994
rect 34317 2884 34351 2922
rect 34317 2812 34351 2850
rect 34317 2740 34351 2778
rect 34317 2668 34351 2706
rect 34317 2596 34351 2634
rect 34317 2524 34351 2562
rect 34317 2452 34351 2490
rect 34317 2380 34351 2418
rect 34317 2308 34351 2346
rect 34317 2236 34351 2274
rect 34317 2164 34351 2202
rect 34317 2092 34351 2130
rect 34317 2020 34351 2058
rect 34317 1948 34351 1986
rect 34317 1876 34351 1914
rect 34317 1804 34351 1842
rect 34317 1732 34351 1770
rect 34317 1660 34351 1698
rect 34317 1588 34351 1626
rect 34317 1516 34351 1554
rect 34317 1444 34351 1482
rect 34317 1372 34351 1410
rect 34317 1300 34351 1338
rect 34317 1228 34351 1266
rect 34317 1159 34351 1194
rect 34413 3100 34447 3135
rect 34413 3028 34447 3066
rect 34413 2956 34447 2994
rect 34413 2884 34447 2922
rect 34413 2812 34447 2850
rect 34413 2740 34447 2778
rect 34413 2668 34447 2706
rect 34413 2596 34447 2634
rect 34413 2524 34447 2562
rect 34413 2452 34447 2490
rect 34413 2380 34447 2418
rect 34413 2308 34447 2346
rect 34413 2236 34447 2274
rect 34413 2164 34447 2202
rect 34413 2092 34447 2130
rect 34413 2020 34447 2058
rect 34413 1948 34447 1986
rect 34413 1876 34447 1914
rect 34413 1804 34447 1842
rect 34413 1732 34447 1770
rect 34413 1660 34447 1698
rect 34413 1588 34447 1626
rect 34413 1516 34447 1554
rect 34413 1444 34447 1482
rect 34413 1372 34447 1410
rect 34413 1300 34447 1338
rect 34413 1228 34447 1266
rect 34413 1159 34447 1194
rect 34509 3100 34543 3135
rect 34509 3028 34543 3066
rect 34509 2956 34543 2994
rect 34509 2884 34543 2922
rect 34509 2812 34543 2850
rect 34509 2740 34543 2778
rect 34509 2668 34543 2706
rect 34509 2596 34543 2634
rect 34509 2524 34543 2562
rect 34509 2452 34543 2490
rect 34509 2380 34543 2418
rect 34509 2308 34543 2346
rect 34509 2236 34543 2274
rect 34509 2164 34543 2202
rect 34509 2092 34543 2130
rect 34509 2020 34543 2058
rect 34509 1948 34543 1986
rect 34509 1876 34543 1914
rect 34509 1804 34543 1842
rect 34509 1732 34543 1770
rect 34509 1660 34543 1698
rect 34509 1588 34543 1626
rect 34509 1516 34543 1554
rect 34509 1444 34543 1482
rect 34509 1372 34543 1410
rect 34509 1300 34543 1338
rect 34509 1228 34543 1266
rect 34509 1159 34543 1194
rect 34605 3100 34639 3135
rect 34605 3028 34639 3066
rect 34605 2956 34639 2994
rect 34605 2884 34639 2922
rect 34605 2812 34639 2850
rect 34605 2740 34639 2778
rect 34605 2668 34639 2706
rect 34605 2596 34639 2634
rect 34605 2524 34639 2562
rect 34605 2452 34639 2490
rect 34605 2380 34639 2418
rect 34605 2308 34639 2346
rect 34605 2236 34639 2274
rect 34605 2164 34639 2202
rect 34605 2092 34639 2130
rect 34605 2020 34639 2058
rect 34605 1948 34639 1986
rect 34605 1876 34639 1914
rect 34605 1804 34639 1842
rect 34605 1732 34639 1770
rect 34605 1660 34639 1698
rect 34605 1588 34639 1626
rect 34605 1516 34639 1554
rect 34605 1444 34639 1482
rect 34605 1372 34639 1410
rect 34605 1300 34639 1338
rect 34605 1228 34639 1266
rect 34605 1159 34639 1194
rect 34701 3100 34735 3135
rect 34701 3028 34735 3066
rect 34701 2956 34735 2994
rect 34701 2884 34735 2922
rect 34701 2812 34735 2850
rect 34701 2740 34735 2778
rect 34701 2668 34735 2706
rect 34701 2596 34735 2634
rect 34701 2524 34735 2562
rect 34701 2452 34735 2490
rect 34701 2380 34735 2418
rect 34701 2308 34735 2346
rect 34701 2236 34735 2274
rect 34701 2164 34735 2202
rect 34701 2092 34735 2130
rect 34701 2020 34735 2058
rect 34701 1948 34735 1986
rect 34701 1876 34735 1914
rect 34701 1804 34735 1842
rect 34701 1732 34735 1770
rect 34701 1660 34735 1698
rect 34701 1588 34735 1626
rect 34701 1516 34735 1554
rect 34701 1444 34735 1482
rect 34701 1372 34735 1410
rect 34701 1300 34735 1338
rect 34701 1228 34735 1266
rect 34701 1159 34735 1194
rect 34797 3100 34831 3135
rect 34797 3028 34831 3066
rect 34797 2956 34831 2994
rect 34797 2884 34831 2922
rect 34797 2812 34831 2850
rect 34797 2740 34831 2778
rect 34797 2668 34831 2706
rect 34797 2596 34831 2634
rect 34797 2524 34831 2562
rect 34797 2452 34831 2490
rect 34797 2380 34831 2418
rect 34797 2308 34831 2346
rect 34797 2236 34831 2274
rect 34797 2164 34831 2202
rect 34797 2092 34831 2130
rect 34797 2020 34831 2058
rect 34797 1948 34831 1986
rect 34797 1876 34831 1914
rect 34797 1804 34831 1842
rect 34797 1732 34831 1770
rect 34797 1660 34831 1698
rect 34797 1588 34831 1626
rect 34797 1516 34831 1554
rect 34797 1444 34831 1482
rect 34797 1372 34831 1410
rect 34797 1300 34831 1338
rect 34797 1228 34831 1266
rect 34797 1159 34831 1194
rect 34893 3100 34927 3135
rect 34893 3028 34927 3066
rect 34893 2956 34927 2994
rect 34893 2884 34927 2922
rect 34893 2812 34927 2850
rect 34893 2740 34927 2778
rect 34893 2668 34927 2706
rect 34893 2596 34927 2634
rect 34893 2524 34927 2562
rect 34893 2452 34927 2490
rect 34893 2380 34927 2418
rect 34893 2308 34927 2346
rect 34893 2236 34927 2274
rect 34893 2164 34927 2202
rect 34893 2092 34927 2130
rect 34893 2020 34927 2058
rect 34893 1948 34927 1986
rect 34893 1876 34927 1914
rect 34893 1804 34927 1842
rect 34893 1732 34927 1770
rect 34893 1660 34927 1698
rect 34893 1588 34927 1626
rect 34893 1516 34927 1554
rect 34893 1444 34927 1482
rect 34893 1372 34927 1410
rect 34893 1300 34927 1338
rect 34893 1228 34927 1266
rect 34893 1159 34927 1194
rect 34989 3100 35023 3135
rect 34989 3028 35023 3066
rect 34989 2956 35023 2994
rect 34989 2884 35023 2922
rect 34989 2812 35023 2850
rect 34989 2740 35023 2778
rect 34989 2668 35023 2706
rect 34989 2596 35023 2634
rect 34989 2524 35023 2562
rect 34989 2452 35023 2490
rect 34989 2380 35023 2418
rect 34989 2308 35023 2346
rect 34989 2236 35023 2274
rect 34989 2164 35023 2202
rect 34989 2092 35023 2130
rect 34989 2020 35023 2058
rect 34989 1948 35023 1986
rect 34989 1876 35023 1914
rect 34989 1804 35023 1842
rect 34989 1732 35023 1770
rect 34989 1660 35023 1698
rect 34989 1588 35023 1626
rect 34989 1516 35023 1554
rect 34989 1444 35023 1482
rect 34989 1372 35023 1410
rect 34989 1300 35023 1338
rect 34989 1228 35023 1266
rect 34989 1159 35023 1194
rect 35085 3100 35119 3135
rect 35085 3028 35119 3066
rect 35085 2956 35119 2994
rect 35085 2884 35119 2922
rect 35085 2812 35119 2850
rect 35085 2740 35119 2778
rect 35085 2668 35119 2706
rect 35085 2596 35119 2634
rect 35085 2524 35119 2562
rect 35085 2452 35119 2490
rect 35085 2380 35119 2418
rect 35085 2308 35119 2346
rect 35085 2236 35119 2274
rect 35085 2164 35119 2202
rect 35085 2092 35119 2130
rect 35085 2020 35119 2058
rect 35085 1948 35119 1986
rect 35085 1876 35119 1914
rect 35085 1804 35119 1842
rect 35085 1732 35119 1770
rect 35085 1660 35119 1698
rect 35085 1588 35119 1626
rect 35085 1516 35119 1554
rect 35085 1444 35119 1482
rect 35085 1372 35119 1410
rect 35085 1300 35119 1338
rect 35085 1228 35119 1266
rect 35085 1159 35119 1194
rect 35181 3100 35215 3135
rect 35181 3028 35215 3066
rect 35181 2956 35215 2994
rect 35181 2884 35215 2922
rect 35181 2812 35215 2850
rect 35181 2740 35215 2778
rect 35181 2668 35215 2706
rect 35181 2596 35215 2634
rect 35181 2524 35215 2562
rect 35181 2452 35215 2490
rect 35181 2380 35215 2418
rect 35181 2308 35215 2346
rect 35181 2236 35215 2274
rect 35181 2164 35215 2202
rect 35181 2092 35215 2130
rect 35181 2020 35215 2058
rect 35181 1948 35215 1986
rect 35181 1876 35215 1914
rect 35181 1804 35215 1842
rect 35181 1732 35215 1770
rect 35181 1660 35215 1698
rect 35181 1588 35215 1626
rect 35181 1516 35215 1554
rect 35181 1444 35215 1482
rect 35181 1372 35215 1410
rect 35181 1300 35215 1338
rect 35181 1228 35215 1266
rect 35181 1159 35215 1194
rect 35277 3100 35311 3135
rect 35277 3028 35311 3066
rect 35277 2956 35311 2994
rect 35277 2884 35311 2922
rect 35277 2812 35311 2850
rect 35277 2740 35311 2778
rect 35277 2668 35311 2706
rect 35277 2596 35311 2634
rect 35277 2524 35311 2562
rect 35277 2452 35311 2490
rect 35277 2380 35311 2418
rect 35277 2308 35311 2346
rect 35277 2236 35311 2274
rect 35277 2164 35311 2202
rect 35277 2092 35311 2130
rect 35277 2020 35311 2058
rect 35277 1948 35311 1986
rect 35277 1876 35311 1914
rect 35277 1804 35311 1842
rect 35277 1732 35311 1770
rect 35277 1660 35311 1698
rect 35277 1588 35311 1626
rect 35277 1516 35311 1554
rect 35277 1444 35311 1482
rect 35277 1372 35311 1410
rect 35277 1300 35311 1338
rect 35277 1228 35311 1266
rect 35277 1159 35311 1194
rect 35373 3100 35407 3135
rect 35373 3028 35407 3066
rect 35373 2956 35407 2994
rect 35373 2884 35407 2922
rect 35373 2812 35407 2850
rect 35373 2740 35407 2778
rect 35373 2668 35407 2706
rect 35373 2596 35407 2634
rect 35373 2524 35407 2562
rect 35373 2452 35407 2490
rect 35373 2380 35407 2418
rect 35373 2308 35407 2346
rect 35373 2236 35407 2274
rect 35373 2164 35407 2202
rect 35373 2092 35407 2130
rect 35373 2020 35407 2058
rect 35373 1948 35407 1986
rect 35373 1876 35407 1914
rect 35373 1804 35407 1842
rect 35373 1732 35407 1770
rect 35373 1660 35407 1698
rect 35373 1588 35407 1626
rect 35373 1516 35407 1554
rect 35373 1444 35407 1482
rect 35373 1372 35407 1410
rect 35373 1300 35407 1338
rect 35373 1228 35407 1266
rect 35373 1159 35407 1194
rect 35469 3100 35503 3135
rect 35469 3028 35503 3066
rect 35469 2956 35503 2994
rect 35469 2884 35503 2922
rect 35469 2812 35503 2850
rect 35469 2740 35503 2778
rect 35469 2668 35503 2706
rect 35469 2596 35503 2634
rect 35469 2524 35503 2562
rect 35469 2452 35503 2490
rect 35469 2380 35503 2418
rect 35469 2308 35503 2346
rect 35469 2236 35503 2274
rect 35469 2164 35503 2202
rect 35469 2092 35503 2130
rect 35469 2020 35503 2058
rect 35469 1948 35503 1986
rect 35469 1876 35503 1914
rect 35469 1804 35503 1842
rect 35469 1732 35503 1770
rect 35469 1660 35503 1698
rect 35469 1588 35503 1626
rect 35469 1516 35503 1554
rect 35469 1444 35503 1482
rect 35469 1372 35503 1410
rect 35469 1300 35503 1338
rect 35469 1228 35503 1266
rect 35469 1159 35503 1194
rect 35565 3100 35599 3135
rect 35565 3028 35599 3066
rect 35565 2956 35599 2994
rect 35565 2884 35599 2922
rect 35565 2812 35599 2850
rect 35565 2740 35599 2778
rect 35565 2668 35599 2706
rect 35565 2596 35599 2634
rect 35565 2524 35599 2562
rect 35565 2452 35599 2490
rect 35565 2380 35599 2418
rect 35565 2308 35599 2346
rect 35565 2236 35599 2274
rect 35565 2164 35599 2202
rect 35565 2092 35599 2130
rect 35565 2020 35599 2058
rect 35565 1948 35599 1986
rect 35565 1876 35599 1914
rect 35565 1804 35599 1842
rect 35565 1732 35599 1770
rect 35565 1660 35599 1698
rect 35565 1588 35599 1626
rect 35565 1516 35599 1554
rect 35565 1444 35599 1482
rect 35565 1372 35599 1410
rect 35565 1300 35599 1338
rect 35565 1228 35599 1266
rect 35565 1159 35599 1194
rect 35661 3100 35695 3135
rect 35661 3028 35695 3066
rect 35661 2956 35695 2994
rect 35661 2884 35695 2922
rect 35661 2812 35695 2850
rect 35661 2740 35695 2778
rect 35661 2668 35695 2706
rect 35661 2596 35695 2634
rect 35661 2524 35695 2562
rect 35661 2452 35695 2490
rect 35661 2380 35695 2418
rect 35661 2308 35695 2346
rect 35661 2236 35695 2274
rect 35661 2164 35695 2202
rect 35661 2092 35695 2130
rect 35661 2020 35695 2058
rect 35661 1948 35695 1986
rect 35661 1876 35695 1914
rect 35661 1804 35695 1842
rect 35661 1732 35695 1770
rect 35661 1660 35695 1698
rect 35661 1588 35695 1626
rect 35661 1516 35695 1554
rect 35661 1444 35695 1482
rect 35661 1372 35695 1410
rect 35661 1300 35695 1338
rect 35661 1228 35695 1266
rect 35661 1159 35695 1194
rect 35757 3100 35791 3135
rect 35757 3028 35791 3066
rect 35757 2956 35791 2994
rect 35757 2884 35791 2922
rect 35757 2812 35791 2850
rect 35757 2740 35791 2778
rect 35757 2668 35791 2706
rect 35757 2596 35791 2634
rect 35757 2524 35791 2562
rect 35757 2452 35791 2490
rect 35757 2380 35791 2418
rect 35757 2308 35791 2346
rect 35757 2236 35791 2274
rect 35757 2164 35791 2202
rect 35757 2092 35791 2130
rect 35757 2020 35791 2058
rect 35757 1948 35791 1986
rect 35757 1876 35791 1914
rect 35757 1804 35791 1842
rect 35757 1732 35791 1770
rect 35757 1660 35791 1698
rect 35757 1588 35791 1626
rect 35757 1516 35791 1554
rect 35757 1444 35791 1482
rect 35757 1372 35791 1410
rect 35757 1300 35791 1338
rect 35757 1228 35791 1266
rect 35757 1159 35791 1194
rect 35853 3100 35887 3135
rect 35853 3028 35887 3066
rect 35853 2956 35887 2994
rect 35853 2884 35887 2922
rect 35853 2812 35887 2850
rect 35853 2740 35887 2778
rect 35853 2668 35887 2706
rect 35853 2596 35887 2634
rect 35853 2524 35887 2562
rect 35853 2452 35887 2490
rect 35853 2380 35887 2418
rect 35853 2308 35887 2346
rect 35853 2236 35887 2274
rect 35853 2164 35887 2202
rect 35853 2092 35887 2130
rect 35853 2020 35887 2058
rect 35853 1948 35887 1986
rect 35853 1876 35887 1914
rect 35853 1804 35887 1842
rect 35853 1732 35887 1770
rect 35853 1660 35887 1698
rect 35853 1588 35887 1626
rect 35853 1516 35887 1554
rect 35853 1444 35887 1482
rect 35853 1372 35887 1410
rect 35853 1300 35887 1338
rect 35853 1228 35887 1266
rect 35853 1159 35887 1194
rect 35949 3100 35983 3135
rect 35949 3028 35983 3066
rect 35949 2956 35983 2994
rect 35949 2884 35983 2922
rect 35949 2812 35983 2850
rect 35949 2740 35983 2778
rect 35949 2668 35983 2706
rect 35949 2596 35983 2634
rect 35949 2524 35983 2562
rect 35949 2452 35983 2490
rect 35949 2380 35983 2418
rect 35949 2308 35983 2346
rect 35949 2236 35983 2274
rect 35949 2164 35983 2202
rect 35949 2092 35983 2130
rect 35949 2020 35983 2058
rect 35949 1948 35983 1986
rect 35949 1876 35983 1914
rect 35949 1804 35983 1842
rect 35949 1732 35983 1770
rect 35949 1660 35983 1698
rect 35949 1588 35983 1626
rect 35949 1516 35983 1554
rect 35949 1444 35983 1482
rect 35949 1372 35983 1410
rect 35949 1300 35983 1338
rect 35949 1228 35983 1266
rect 35949 1159 35983 1194
rect 36045 3100 36079 3135
rect 36045 3028 36079 3066
rect 36045 2956 36079 2994
rect 36045 2884 36079 2922
rect 36045 2812 36079 2850
rect 36045 2740 36079 2778
rect 36045 2668 36079 2706
rect 36045 2596 36079 2634
rect 36045 2524 36079 2562
rect 36045 2452 36079 2490
rect 36045 2380 36079 2418
rect 36045 2308 36079 2346
rect 36045 2236 36079 2274
rect 36045 2164 36079 2202
rect 36045 2092 36079 2130
rect 36045 2020 36079 2058
rect 36045 1948 36079 1986
rect 36045 1876 36079 1914
rect 36045 1804 36079 1842
rect 36045 1732 36079 1770
rect 36045 1660 36079 1698
rect 36045 1588 36079 1626
rect 36045 1516 36079 1554
rect 36045 1444 36079 1482
rect 36045 1372 36079 1410
rect 36045 1300 36079 1338
rect 36045 1228 36079 1266
rect 36045 1159 36079 1194
rect 36141 3100 36175 3135
rect 36141 3028 36175 3066
rect 36141 2956 36175 2994
rect 36141 2884 36175 2922
rect 36141 2812 36175 2850
rect 36141 2740 36175 2778
rect 36141 2668 36175 2706
rect 36141 2596 36175 2634
rect 36141 2524 36175 2562
rect 36141 2452 36175 2490
rect 36141 2380 36175 2418
rect 36141 2308 36175 2346
rect 36141 2236 36175 2274
rect 36141 2164 36175 2202
rect 36141 2092 36175 2130
rect 36141 2020 36175 2058
rect 36141 1948 36175 1986
rect 36141 1876 36175 1914
rect 36141 1804 36175 1842
rect 36141 1732 36175 1770
rect 36141 1660 36175 1698
rect 36141 1588 36175 1626
rect 36141 1516 36175 1554
rect 36141 1444 36175 1482
rect 36141 1372 36175 1410
rect 36141 1300 36175 1338
rect 36141 1228 36175 1266
rect 36141 1159 36175 1194
rect 36237 3100 36271 3135
rect 36237 3028 36271 3066
rect 36237 2956 36271 2994
rect 36237 2884 36271 2922
rect 36237 2812 36271 2850
rect 36237 2740 36271 2778
rect 36237 2668 36271 2706
rect 36237 2596 36271 2634
rect 36237 2524 36271 2562
rect 36237 2452 36271 2490
rect 36237 2380 36271 2418
rect 36237 2308 36271 2346
rect 36237 2236 36271 2274
rect 36237 2164 36271 2202
rect 36237 2092 36271 2130
rect 36237 2020 36271 2058
rect 36237 1948 36271 1986
rect 36237 1876 36271 1914
rect 36237 1804 36271 1842
rect 36237 1732 36271 1770
rect 36237 1660 36271 1698
rect 36237 1588 36271 1626
rect 36237 1516 36271 1554
rect 36237 1444 36271 1482
rect 36237 1372 36271 1410
rect 36237 1300 36271 1338
rect 36237 1228 36271 1266
rect 36237 1159 36271 1194
rect 36333 3100 36367 3135
rect 36333 3028 36367 3066
rect 36333 2956 36367 2994
rect 36333 2884 36367 2922
rect 36333 2812 36367 2850
rect 36333 2740 36367 2778
rect 36333 2668 36367 2706
rect 36333 2596 36367 2634
rect 36333 2524 36367 2562
rect 36333 2452 36367 2490
rect 36333 2380 36367 2418
rect 36333 2308 36367 2346
rect 36333 2236 36367 2274
rect 36333 2164 36367 2202
rect 36333 2092 36367 2130
rect 36333 2020 36367 2058
rect 36333 1948 36367 1986
rect 36333 1876 36367 1914
rect 36333 1804 36367 1842
rect 36333 1732 36367 1770
rect 36333 1660 36367 1698
rect 36333 1588 36367 1626
rect 36333 1516 36367 1554
rect 36333 1444 36367 1482
rect 36333 1372 36367 1410
rect 36333 1300 36367 1338
rect 36333 1228 36367 1266
rect 36333 1159 36367 1194
rect 36429 3100 36463 3135
rect 36429 3028 36463 3066
rect 36429 2956 36463 2994
rect 36429 2884 36463 2922
rect 36429 2812 36463 2850
rect 36429 2740 36463 2778
rect 36429 2668 36463 2706
rect 36429 2596 36463 2634
rect 36429 2524 36463 2562
rect 36429 2452 36463 2490
rect 36429 2380 36463 2418
rect 36429 2308 36463 2346
rect 36429 2236 36463 2274
rect 36429 2164 36463 2202
rect 36429 2092 36463 2130
rect 36429 2020 36463 2058
rect 36429 1948 36463 1986
rect 36429 1876 36463 1914
rect 36429 1804 36463 1842
rect 36429 1732 36463 1770
rect 36429 1660 36463 1698
rect 36429 1588 36463 1626
rect 36429 1516 36463 1554
rect 36429 1444 36463 1482
rect 36429 1372 36463 1410
rect 36429 1300 36463 1338
rect 36429 1228 36463 1266
rect 36429 1159 36463 1194
rect 36525 3100 36559 3135
rect 36525 3028 36559 3066
rect 36525 2956 36559 2994
rect 36525 2884 36559 2922
rect 36525 2812 36559 2850
rect 36525 2740 36559 2778
rect 36525 2668 36559 2706
rect 36525 2596 36559 2634
rect 36525 2524 36559 2562
rect 36525 2452 36559 2490
rect 36525 2380 36559 2418
rect 36525 2308 36559 2346
rect 36525 2236 36559 2274
rect 36525 2164 36559 2202
rect 36525 2092 36559 2130
rect 36525 2020 36559 2058
rect 36525 1948 36559 1986
rect 36525 1876 36559 1914
rect 36525 1804 36559 1842
rect 36525 1732 36559 1770
rect 36525 1660 36559 1698
rect 36525 1588 36559 1626
rect 36525 1516 36559 1554
rect 36525 1444 36559 1482
rect 36525 1372 36559 1410
rect 36525 1300 36559 1338
rect 36525 1228 36559 1266
rect 36525 1159 36559 1194
rect 36621 3100 36655 3135
rect 36621 3028 36655 3066
rect 36621 2956 36655 2994
rect 36621 2884 36655 2922
rect 36621 2812 36655 2850
rect 36621 2740 36655 2778
rect 36621 2668 36655 2706
rect 36621 2596 36655 2634
rect 36621 2524 36655 2562
rect 36621 2452 36655 2490
rect 36621 2380 36655 2418
rect 36621 2308 36655 2346
rect 36621 2236 36655 2274
rect 36621 2164 36655 2202
rect 36621 2092 36655 2130
rect 36621 2020 36655 2058
rect 36621 1948 36655 1986
rect 36621 1876 36655 1914
rect 36621 1804 36655 1842
rect 36621 1732 36655 1770
rect 36621 1660 36655 1698
rect 36621 1588 36655 1626
rect 36621 1516 36655 1554
rect 36621 1444 36655 1482
rect 36621 1372 36655 1410
rect 36621 1300 36655 1338
rect 36621 1228 36655 1266
rect 36621 1159 36655 1194
rect 36717 3100 36751 3135
rect 36717 3028 36751 3066
rect 36717 2956 36751 2994
rect 36717 2884 36751 2922
rect 36717 2812 36751 2850
rect 36717 2740 36751 2778
rect 36717 2668 36751 2706
rect 36717 2596 36751 2634
rect 36717 2524 36751 2562
rect 36717 2452 36751 2490
rect 36717 2380 36751 2418
rect 36717 2308 36751 2346
rect 36717 2236 36751 2274
rect 36717 2164 36751 2202
rect 36717 2092 36751 2130
rect 36717 2020 36751 2058
rect 36717 1948 36751 1986
rect 36717 1876 36751 1914
rect 36717 1804 36751 1842
rect 36717 1732 36751 1770
rect 36717 1660 36751 1698
rect 36717 1588 36751 1626
rect 36717 1516 36751 1554
rect 36717 1444 36751 1482
rect 36717 1372 36751 1410
rect 36717 1300 36751 1338
rect 36717 1228 36751 1266
rect 36717 1159 36751 1194
rect 36813 3100 36847 3135
rect 36813 3028 36847 3066
rect 36813 2956 36847 2994
rect 36813 2884 36847 2922
rect 36813 2812 36847 2850
rect 36813 2740 36847 2778
rect 36813 2668 36847 2706
rect 36813 2596 36847 2634
rect 36813 2524 36847 2562
rect 36813 2452 36847 2490
rect 36813 2380 36847 2418
rect 36813 2308 36847 2346
rect 36813 2236 36847 2274
rect 36813 2164 36847 2202
rect 36813 2092 36847 2130
rect 36813 2020 36847 2058
rect 36813 1948 36847 1986
rect 36813 1876 36847 1914
rect 36813 1804 36847 1842
rect 36813 1732 36847 1770
rect 36813 1660 36847 1698
rect 36813 1588 36847 1626
rect 36813 1516 36847 1554
rect 36813 1444 36847 1482
rect 36813 1372 36847 1410
rect 36813 1300 36847 1338
rect 36813 1228 36847 1266
rect 36813 1159 36847 1194
rect 36909 3100 36943 3135
rect 36909 3028 36943 3066
rect 36909 2956 36943 2994
rect 36909 2884 36943 2922
rect 36909 2812 36943 2850
rect 36909 2740 36943 2778
rect 36909 2668 36943 2706
rect 36909 2596 36943 2634
rect 36909 2524 36943 2562
rect 36909 2452 36943 2490
rect 36909 2380 36943 2418
rect 36909 2308 36943 2346
rect 36909 2236 36943 2274
rect 36909 2164 36943 2202
rect 36909 2092 36943 2130
rect 36909 2020 36943 2058
rect 36909 1948 36943 1986
rect 36909 1876 36943 1914
rect 36909 1804 36943 1842
rect 36909 1732 36943 1770
rect 36909 1660 36943 1698
rect 36909 1588 36943 1626
rect 36909 1516 36943 1554
rect 36909 1444 36943 1482
rect 36909 1372 36943 1410
rect 36909 1300 36943 1338
rect 36909 1228 36943 1266
rect 36909 1159 36943 1194
rect 37005 3100 37039 3135
rect 37005 3028 37039 3066
rect 37005 2956 37039 2994
rect 37005 2884 37039 2922
rect 37005 2812 37039 2850
rect 37005 2740 37039 2778
rect 37005 2668 37039 2706
rect 37005 2596 37039 2634
rect 37005 2524 37039 2562
rect 37005 2452 37039 2490
rect 37005 2380 37039 2418
rect 37005 2308 37039 2346
rect 37005 2236 37039 2274
rect 37005 2164 37039 2202
rect 37005 2092 37039 2130
rect 37005 2020 37039 2058
rect 37005 1948 37039 1986
rect 37005 1876 37039 1914
rect 37005 1804 37039 1842
rect 37005 1732 37039 1770
rect 37005 1660 37039 1698
rect 37005 1588 37039 1626
rect 37005 1516 37039 1554
rect 37005 1444 37039 1482
rect 37005 1372 37039 1410
rect 37005 1300 37039 1338
rect 37005 1228 37039 1266
rect 37005 1159 37039 1194
rect 37101 3100 37135 3135
rect 37101 3028 37135 3066
rect 37101 2956 37135 2994
rect 37101 2884 37135 2922
rect 37101 2812 37135 2850
rect 37101 2740 37135 2778
rect 37101 2668 37135 2706
rect 37101 2596 37135 2634
rect 37101 2524 37135 2562
rect 37101 2452 37135 2490
rect 37101 2380 37135 2418
rect 37101 2308 37135 2346
rect 37101 2236 37135 2274
rect 37101 2164 37135 2202
rect 37101 2092 37135 2130
rect 37101 2020 37135 2058
rect 37101 1948 37135 1986
rect 37101 1876 37135 1914
rect 37101 1804 37135 1842
rect 37101 1732 37135 1770
rect 37101 1660 37135 1698
rect 37101 1588 37135 1626
rect 37101 1516 37135 1554
rect 37101 1444 37135 1482
rect 37101 1372 37135 1410
rect 37101 1300 37135 1338
rect 37101 1228 37135 1266
rect 37101 1159 37135 1194
rect 37197 3100 37231 3135
rect 37197 3028 37231 3066
rect 37197 2956 37231 2994
rect 37197 2884 37231 2922
rect 37197 2812 37231 2850
rect 37197 2740 37231 2778
rect 37197 2668 37231 2706
rect 37197 2596 37231 2634
rect 37197 2524 37231 2562
rect 37197 2452 37231 2490
rect 37197 2380 37231 2418
rect 37197 2308 37231 2346
rect 37197 2236 37231 2274
rect 37197 2164 37231 2202
rect 37197 2092 37231 2130
rect 37197 2020 37231 2058
rect 37197 1948 37231 1986
rect 37197 1876 37231 1914
rect 37197 1804 37231 1842
rect 37197 1732 37231 1770
rect 37197 1660 37231 1698
rect 37197 1588 37231 1626
rect 37197 1516 37231 1554
rect 37197 1444 37231 1482
rect 37197 1372 37231 1410
rect 37197 1300 37231 1338
rect 37197 1228 37231 1266
rect 37197 1159 37231 1194
rect 37293 3100 37327 3135
rect 37293 3028 37327 3066
rect 37293 2956 37327 2994
rect 37293 2884 37327 2922
rect 37293 2812 37327 2850
rect 37293 2740 37327 2778
rect 37293 2668 37327 2706
rect 37293 2596 37327 2634
rect 37293 2524 37327 2562
rect 37293 2452 37327 2490
rect 37293 2380 37327 2418
rect 37293 2308 37327 2346
rect 37293 2236 37327 2274
rect 37293 2164 37327 2202
rect 37293 2092 37327 2130
rect 37293 2020 37327 2058
rect 37293 1948 37327 1986
rect 37293 1876 37327 1914
rect 37293 1804 37327 1842
rect 37293 1732 37327 1770
rect 37293 1660 37327 1698
rect 37293 1588 37327 1626
rect 37293 1516 37327 1554
rect 37293 1444 37327 1482
rect 37293 1372 37327 1410
rect 37293 1300 37327 1338
rect 37293 1228 37327 1266
rect 37293 1159 37327 1194
rect 37389 3100 37423 3135
rect 37389 3028 37423 3066
rect 37389 2956 37423 2994
rect 37389 2884 37423 2922
rect 37389 2812 37423 2850
rect 37389 2740 37423 2778
rect 37389 2668 37423 2706
rect 37389 2596 37423 2634
rect 37389 2524 37423 2562
rect 37389 2452 37423 2490
rect 37389 2380 37423 2418
rect 37389 2308 37423 2346
rect 37389 2236 37423 2274
rect 37389 2164 37423 2202
rect 37389 2092 37423 2130
rect 37389 2020 37423 2058
rect 37389 1948 37423 1986
rect 37389 1876 37423 1914
rect 37389 1804 37423 1842
rect 37389 1732 37423 1770
rect 37389 1660 37423 1698
rect 37389 1588 37423 1626
rect 37389 1516 37423 1554
rect 37389 1444 37423 1482
rect 37389 1372 37423 1410
rect 37389 1300 37423 1338
rect 37389 1228 37423 1266
rect 37389 1159 37423 1194
rect 37485 3100 37519 3135
rect 37485 3028 37519 3066
rect 37485 2956 37519 2994
rect 37485 2884 37519 2922
rect 37485 2812 37519 2850
rect 37485 2740 37519 2778
rect 37485 2668 37519 2706
rect 37485 2596 37519 2634
rect 37485 2524 37519 2562
rect 37485 2452 37519 2490
rect 37485 2380 37519 2418
rect 37485 2308 37519 2346
rect 37485 2236 37519 2274
rect 37485 2164 37519 2202
rect 37485 2092 37519 2130
rect 37485 2020 37519 2058
rect 37485 1948 37519 1986
rect 37485 1876 37519 1914
rect 37485 1804 37519 1842
rect 37485 1732 37519 1770
rect 37485 1660 37519 1698
rect 37485 1588 37519 1626
rect 37485 1516 37519 1554
rect 37485 1444 37519 1482
rect 37485 1372 37519 1410
rect 37485 1300 37519 1338
rect 37485 1228 37519 1266
rect 37485 1159 37519 1194
rect 37581 3100 37615 3135
rect 37581 3028 37615 3066
rect 37581 2956 37615 2994
rect 37581 2884 37615 2922
rect 37581 2812 37615 2850
rect 37581 2740 37615 2778
rect 37581 2668 37615 2706
rect 37581 2596 37615 2634
rect 37581 2524 37615 2562
rect 37581 2452 37615 2490
rect 37581 2380 37615 2418
rect 37581 2308 37615 2346
rect 37581 2236 37615 2274
rect 37581 2164 37615 2202
rect 37581 2092 37615 2130
rect 37581 2020 37615 2058
rect 37581 1948 37615 1986
rect 37581 1876 37615 1914
rect 37581 1804 37615 1842
rect 37581 1732 37615 1770
rect 37581 1660 37615 1698
rect 37581 1588 37615 1626
rect 37581 1516 37615 1554
rect 37581 1444 37615 1482
rect 37581 1372 37615 1410
rect 37581 1300 37615 1338
rect 37581 1228 37615 1266
rect 37581 1159 37615 1194
rect 37677 3100 37711 3135
rect 37677 3028 37711 3066
rect 37677 2956 37711 2994
rect 37677 2884 37711 2922
rect 37677 2812 37711 2850
rect 37677 2740 37711 2778
rect 37677 2668 37711 2706
rect 37677 2596 37711 2634
rect 37677 2524 37711 2562
rect 37677 2452 37711 2490
rect 37677 2380 37711 2418
rect 37677 2308 37711 2346
rect 37677 2236 37711 2274
rect 37677 2164 37711 2202
rect 37677 2092 37711 2130
rect 37677 2020 37711 2058
rect 37677 1948 37711 1986
rect 37677 1876 37711 1914
rect 37677 1804 37711 1842
rect 37677 1732 37711 1770
rect 37677 1660 37711 1698
rect 37677 1588 37711 1626
rect 37677 1516 37711 1554
rect 37677 1444 37711 1482
rect 37677 1372 37711 1410
rect 37677 1300 37711 1338
rect 37677 1228 37711 1266
rect 37677 1159 37711 1194
rect 37773 3100 37807 3135
rect 37773 3028 37807 3066
rect 37773 2956 37807 2994
rect 37773 2884 37807 2922
rect 37773 2812 37807 2850
rect 37773 2740 37807 2778
rect 37773 2668 37807 2706
rect 37773 2596 37807 2634
rect 37773 2524 37807 2562
rect 37773 2452 37807 2490
rect 37773 2380 37807 2418
rect 37773 2308 37807 2346
rect 37773 2236 37807 2274
rect 37773 2164 37807 2202
rect 37773 2092 37807 2130
rect 37773 2020 37807 2058
rect 37773 1948 37807 1986
rect 37773 1876 37807 1914
rect 37773 1804 37807 1842
rect 37773 1732 37807 1770
rect 37773 1660 37807 1698
rect 37773 1588 37807 1626
rect 37773 1516 37807 1554
rect 37773 1444 37807 1482
rect 37773 1372 37807 1410
rect 37773 1300 37807 1338
rect 37773 1228 37807 1266
rect 37773 1159 37807 1194
rect 37869 3100 37903 3135
rect 37869 3028 37903 3066
rect 37869 2956 37903 2994
rect 37869 2884 37903 2922
rect 37869 2812 37903 2850
rect 37869 2740 37903 2778
rect 37869 2668 37903 2706
rect 37869 2596 37903 2634
rect 37869 2524 37903 2562
rect 37869 2452 37903 2490
rect 37869 2380 37903 2418
rect 37869 2308 37903 2346
rect 37869 2236 37903 2274
rect 37869 2164 37903 2202
rect 37869 2092 37903 2130
rect 37869 2020 37903 2058
rect 37869 1948 37903 1986
rect 37869 1876 37903 1914
rect 37869 1804 37903 1842
rect 37869 1732 37903 1770
rect 37869 1660 37903 1698
rect 37869 1588 37903 1626
rect 37869 1516 37903 1554
rect 37869 1444 37903 1482
rect 37869 1372 37903 1410
rect 37869 1300 37903 1338
rect 37869 1228 37903 1266
rect 37869 1159 37903 1194
rect 37965 3100 37999 3135
rect 37965 3028 37999 3066
rect 37965 2956 37999 2994
rect 37965 2884 37999 2922
rect 37965 2812 37999 2850
rect 37965 2740 37999 2778
rect 37965 2668 37999 2706
rect 37965 2596 37999 2634
rect 37965 2524 37999 2562
rect 37965 2452 37999 2490
rect 37965 2380 37999 2418
rect 37965 2308 37999 2346
rect 37965 2236 37999 2274
rect 37965 2164 37999 2202
rect 37965 2092 37999 2130
rect 37965 2020 37999 2058
rect 37965 1948 37999 1986
rect 37965 1876 37999 1914
rect 37965 1804 37999 1842
rect 37965 1732 37999 1770
rect 37965 1660 37999 1698
rect 37965 1588 37999 1626
rect 37965 1516 37999 1554
rect 37965 1444 37999 1482
rect 37965 1372 37999 1410
rect 37965 1300 37999 1338
rect 37965 1228 37999 1266
rect 37965 1159 37999 1194
rect 38061 3100 38095 3135
rect 38061 3028 38095 3066
rect 38061 2956 38095 2994
rect 38061 2884 38095 2922
rect 38061 2812 38095 2850
rect 38061 2740 38095 2778
rect 38061 2668 38095 2706
rect 38061 2596 38095 2634
rect 38061 2524 38095 2562
rect 38061 2452 38095 2490
rect 38061 2380 38095 2418
rect 38061 2308 38095 2346
rect 38061 2236 38095 2274
rect 38061 2164 38095 2202
rect 38061 2092 38095 2130
rect 38061 2020 38095 2058
rect 38061 1948 38095 1986
rect 38061 1876 38095 1914
rect 38061 1804 38095 1842
rect 38061 1732 38095 1770
rect 38061 1660 38095 1698
rect 38061 1588 38095 1626
rect 38061 1516 38095 1554
rect 38061 1444 38095 1482
rect 38061 1372 38095 1410
rect 38061 1300 38095 1338
rect 38061 1228 38095 1266
rect 38061 1159 38095 1194
rect 38157 3100 38191 3135
rect 38157 3028 38191 3066
rect 38157 2956 38191 2994
rect 38157 2884 38191 2922
rect 38157 2812 38191 2850
rect 38157 2740 38191 2778
rect 38157 2668 38191 2706
rect 38157 2596 38191 2634
rect 38157 2524 38191 2562
rect 38157 2452 38191 2490
rect 38157 2380 38191 2418
rect 38157 2308 38191 2346
rect 38157 2236 38191 2274
rect 38157 2164 38191 2202
rect 38157 2092 38191 2130
rect 38157 2020 38191 2058
rect 38157 1948 38191 1986
rect 38157 1876 38191 1914
rect 38157 1804 38191 1842
rect 38157 1732 38191 1770
rect 38157 1660 38191 1698
rect 38157 1588 38191 1626
rect 38157 1516 38191 1554
rect 38157 1444 38191 1482
rect 38157 1372 38191 1410
rect 38157 1300 38191 1338
rect 38157 1228 38191 1266
rect 38157 1159 38191 1194
rect 38253 3100 38287 3135
rect 38253 3028 38287 3066
rect 38253 2956 38287 2994
rect 38253 2884 38287 2922
rect 38253 2812 38287 2850
rect 38253 2740 38287 2778
rect 38253 2668 38287 2706
rect 38253 2596 38287 2634
rect 38253 2524 38287 2562
rect 38253 2452 38287 2490
rect 38253 2380 38287 2418
rect 38253 2308 38287 2346
rect 38253 2236 38287 2274
rect 38253 2164 38287 2202
rect 38253 2092 38287 2130
rect 38253 2020 38287 2058
rect 38253 1948 38287 1986
rect 38253 1876 38287 1914
rect 38253 1804 38287 1842
rect 38253 1732 38287 1770
rect 38253 1660 38287 1698
rect 38253 1588 38287 1626
rect 38253 1516 38287 1554
rect 38253 1444 38287 1482
rect 38253 1372 38287 1410
rect 38253 1300 38287 1338
rect 38253 1228 38287 1266
rect 38253 1159 38287 1194
rect 38349 3100 38383 3135
rect 38349 3028 38383 3066
rect 38349 2956 38383 2994
rect 38349 2884 38383 2922
rect 38349 2812 38383 2850
rect 38349 2740 38383 2778
rect 38349 2668 38383 2706
rect 38349 2596 38383 2634
rect 38349 2524 38383 2562
rect 38349 2452 38383 2490
rect 38349 2380 38383 2418
rect 38349 2308 38383 2346
rect 38349 2236 38383 2274
rect 38349 2164 38383 2202
rect 38349 2092 38383 2130
rect 38349 2020 38383 2058
rect 38349 1948 38383 1986
rect 38349 1876 38383 1914
rect 38349 1804 38383 1842
rect 38349 1732 38383 1770
rect 38349 1660 38383 1698
rect 38349 1588 38383 1626
rect 38349 1516 38383 1554
rect 38349 1444 38383 1482
rect 38349 1372 38383 1410
rect 38349 1300 38383 1338
rect 38349 1228 38383 1266
rect 38349 1159 38383 1194
rect 38445 3100 38479 3135
rect 38445 3028 38479 3066
rect 38445 2956 38479 2994
rect 38445 2884 38479 2922
rect 38445 2812 38479 2850
rect 38445 2740 38479 2778
rect 38445 2668 38479 2706
rect 38445 2596 38479 2634
rect 38445 2524 38479 2562
rect 38445 2452 38479 2490
rect 38445 2380 38479 2418
rect 38445 2308 38479 2346
rect 38445 2236 38479 2274
rect 38445 2164 38479 2202
rect 38445 2092 38479 2130
rect 38445 2020 38479 2058
rect 38445 1948 38479 1986
rect 38445 1876 38479 1914
rect 38445 1804 38479 1842
rect 38445 1732 38479 1770
rect 38445 1660 38479 1698
rect 38445 1588 38479 1626
rect 38445 1516 38479 1554
rect 38445 1444 38479 1482
rect 38445 1372 38479 1410
rect 38445 1300 38479 1338
rect 38445 1228 38479 1266
rect 38445 1159 38479 1194
rect 38541 3100 38575 3135
rect 38541 3028 38575 3066
rect 38541 2956 38575 2994
rect 38541 2884 38575 2922
rect 38541 2812 38575 2850
rect 38541 2740 38575 2778
rect 38541 2668 38575 2706
rect 38541 2596 38575 2634
rect 38541 2524 38575 2562
rect 38541 2452 38575 2490
rect 38541 2380 38575 2418
rect 38541 2308 38575 2346
rect 38541 2236 38575 2274
rect 38541 2164 38575 2202
rect 38541 2092 38575 2130
rect 38541 2020 38575 2058
rect 38541 1948 38575 1986
rect 38541 1876 38575 1914
rect 38541 1804 38575 1842
rect 38541 1732 38575 1770
rect 38541 1660 38575 1698
rect 38541 1588 38575 1626
rect 38541 1516 38575 1554
rect 38541 1444 38575 1482
rect 38541 1372 38575 1410
rect 38541 1300 38575 1338
rect 38541 1228 38575 1266
rect 38541 1159 38575 1194
rect 38637 3099 38671 3134
rect 38637 3027 38671 3065
rect 38637 2955 38671 2993
rect 38637 2883 38671 2921
rect 38637 2811 38671 2849
rect 38637 2739 38671 2777
rect 38637 2667 38671 2705
rect 38637 2595 38671 2633
rect 38637 2523 38671 2561
rect 38637 2451 38671 2489
rect 38637 2379 38671 2417
rect 38637 2307 38671 2345
rect 38637 2235 38671 2273
rect 38637 2163 38671 2201
rect 38637 2091 38671 2129
rect 38637 2019 38671 2057
rect 38637 1947 38671 1985
rect 38637 1875 38671 1913
rect 38637 1803 38671 1841
rect 38637 1731 38671 1769
rect 38637 1659 38671 1697
rect 38637 1587 38671 1625
rect 38637 1515 38671 1553
rect 38637 1443 38671 1481
rect 38637 1371 38671 1409
rect 38637 1299 38671 1337
rect 38637 1227 38671 1265
rect 38637 1158 38671 1193
rect 29069 1099 38543 1109
rect 29069 1075 29100 1099
rect 29070 1065 29100 1075
rect 29134 1065 29172 1099
rect 29206 1065 29244 1099
rect 29278 1065 29316 1099
rect 29350 1065 29388 1099
rect 29422 1065 29460 1099
rect 29494 1065 29532 1099
rect 29566 1065 29604 1099
rect 29638 1065 29676 1099
rect 29710 1065 29748 1099
rect 29782 1065 29820 1099
rect 29854 1065 29892 1099
rect 29926 1065 29964 1099
rect 29998 1065 30036 1099
rect 30070 1065 30108 1099
rect 30142 1065 30180 1099
rect 30214 1065 30252 1099
rect 30286 1065 30324 1099
rect 30358 1065 30396 1099
rect 30430 1065 30468 1099
rect 30502 1065 30540 1099
rect 30574 1065 30612 1099
rect 30646 1065 30684 1099
rect 30718 1065 30756 1099
rect 30790 1065 30828 1099
rect 30862 1065 30900 1099
rect 30934 1065 30972 1099
rect 31006 1065 31044 1099
rect 31078 1065 31116 1099
rect 31150 1065 31188 1099
rect 31222 1065 31260 1099
rect 31294 1065 31332 1099
rect 31366 1065 31404 1099
rect 31438 1065 31476 1099
rect 31510 1065 31548 1099
rect 31582 1065 31620 1099
rect 31654 1065 31692 1099
rect 31726 1065 31764 1099
rect 31798 1065 31836 1099
rect 31870 1065 31908 1099
rect 31942 1065 31980 1099
rect 32014 1065 32052 1099
rect 32086 1065 32124 1099
rect 32158 1065 32196 1099
rect 32230 1065 32268 1099
rect 32302 1065 32340 1099
rect 32374 1065 32412 1099
rect 32446 1065 32484 1099
rect 32518 1065 32556 1099
rect 32590 1065 32628 1099
rect 32662 1065 32700 1099
rect 32734 1065 32772 1099
rect 32806 1065 32844 1099
rect 32878 1065 32916 1099
rect 32950 1065 32988 1099
rect 33022 1065 33060 1099
rect 33094 1065 33132 1099
rect 33166 1065 33204 1099
rect 33238 1065 33276 1099
rect 33310 1065 33348 1099
rect 33382 1065 33420 1099
rect 33454 1065 33492 1099
rect 33526 1065 33564 1099
rect 33598 1065 33636 1099
rect 33670 1065 33708 1099
rect 33742 1065 33780 1099
rect 33814 1065 33852 1099
rect 33886 1065 33924 1099
rect 33958 1065 33996 1099
rect 34030 1065 34068 1099
rect 34102 1065 34140 1099
rect 34174 1065 34212 1099
rect 34246 1065 34284 1099
rect 34318 1065 34356 1099
rect 34390 1065 34428 1099
rect 34462 1065 34500 1099
rect 34534 1065 34572 1099
rect 34606 1065 34644 1099
rect 34678 1065 34716 1099
rect 34750 1065 34788 1099
rect 34822 1065 34860 1099
rect 34894 1065 34932 1099
rect 34966 1065 35004 1099
rect 35038 1065 35076 1099
rect 35110 1065 35148 1099
rect 35182 1065 35220 1099
rect 35254 1065 35292 1099
rect 35326 1065 35364 1099
rect 35398 1065 35436 1099
rect 35470 1065 35508 1099
rect 35542 1065 35580 1099
rect 35614 1065 35652 1099
rect 35686 1065 35724 1099
rect 35758 1065 35796 1099
rect 35830 1065 35868 1099
rect 35902 1065 35940 1099
rect 35974 1065 36012 1099
rect 36046 1065 36084 1099
rect 36118 1065 36156 1099
rect 36190 1065 36228 1099
rect 36262 1065 36300 1099
rect 36334 1065 36372 1099
rect 36406 1065 36444 1099
rect 36478 1065 36516 1099
rect 36550 1065 36588 1099
rect 36622 1065 36660 1099
rect 36694 1065 36732 1099
rect 36766 1065 36804 1099
rect 36838 1065 36876 1099
rect 36910 1065 36948 1099
rect 36982 1065 37020 1099
rect 37054 1065 37092 1099
rect 37126 1065 37164 1099
rect 37198 1065 37236 1099
rect 37270 1065 37308 1099
rect 37342 1065 37380 1099
rect 37414 1065 37452 1099
rect 37486 1065 37524 1099
rect 37558 1065 37596 1099
rect 37630 1065 37668 1099
rect 37702 1065 37740 1099
rect 37774 1065 37812 1099
rect 37846 1065 37884 1099
rect 37918 1065 37956 1099
rect 37990 1065 38028 1099
rect 38062 1065 38100 1099
rect 38134 1065 38172 1099
rect 38206 1065 38244 1099
rect 38278 1065 38316 1099
rect 38350 1065 38388 1099
rect 38422 1065 38460 1099
rect 38494 1075 38543 1099
rect 38494 1065 38524 1075
rect 29070 1062 38524 1065
<< viali >>
rect 29200 3189 29234 3223
rect 29272 3189 29306 3223
rect 29344 3189 29378 3223
rect 29416 3189 29450 3223
rect 29488 3189 29522 3223
rect 29560 3189 29594 3223
rect 29632 3189 29666 3223
rect 29704 3189 29738 3223
rect 29776 3189 29810 3223
rect 29848 3189 29882 3223
rect 29920 3189 29954 3223
rect 29992 3189 30026 3223
rect 30064 3189 30098 3223
rect 30136 3189 30170 3223
rect 30208 3189 30242 3223
rect 30280 3189 30314 3223
rect 30352 3189 30386 3223
rect 30424 3189 30458 3223
rect 30496 3189 30530 3223
rect 30568 3189 30602 3223
rect 30640 3189 30674 3223
rect 30712 3189 30746 3223
rect 30784 3189 30818 3223
rect 30856 3189 30890 3223
rect 30928 3189 30962 3223
rect 31000 3189 31034 3223
rect 31072 3189 31106 3223
rect 31144 3189 31178 3223
rect 31216 3189 31250 3223
rect 31288 3189 31322 3223
rect 31360 3189 31394 3223
rect 31432 3189 31466 3223
rect 31504 3189 31538 3223
rect 31576 3189 31610 3223
rect 31648 3189 31682 3223
rect 31720 3189 31754 3223
rect 31792 3189 31826 3223
rect 31864 3189 31898 3223
rect 31936 3189 31970 3223
rect 32008 3189 32042 3223
rect 32080 3189 32114 3223
rect 32152 3189 32186 3223
rect 32224 3189 32258 3223
rect 32296 3189 32330 3223
rect 32368 3189 32402 3223
rect 32440 3189 32474 3223
rect 32512 3189 32546 3223
rect 32584 3189 32618 3223
rect 32656 3189 32690 3223
rect 32728 3189 32762 3223
rect 32800 3189 32834 3223
rect 32872 3189 32906 3223
rect 32944 3189 32978 3223
rect 33016 3189 33050 3223
rect 33088 3189 33122 3223
rect 33160 3189 33194 3223
rect 33232 3189 33266 3223
rect 33304 3189 33338 3223
rect 33376 3189 33410 3223
rect 33448 3189 33482 3223
rect 33520 3189 33554 3223
rect 33592 3189 33626 3223
rect 33664 3189 33698 3223
rect 33736 3189 33770 3223
rect 33808 3189 33842 3223
rect 33880 3189 33914 3223
rect 33952 3189 33986 3223
rect 34024 3189 34058 3223
rect 34096 3189 34130 3223
rect 34168 3189 34202 3223
rect 34240 3189 34274 3223
rect 34312 3189 34346 3223
rect 34384 3189 34418 3223
rect 34456 3189 34490 3223
rect 34528 3189 34562 3223
rect 34600 3189 34634 3223
rect 34672 3189 34706 3223
rect 34744 3189 34778 3223
rect 34816 3189 34850 3223
rect 34888 3189 34922 3223
rect 34960 3189 34994 3223
rect 35032 3189 35066 3223
rect 35104 3189 35138 3223
rect 35176 3189 35210 3223
rect 35248 3189 35282 3223
rect 35320 3189 35354 3223
rect 35392 3189 35426 3223
rect 35464 3189 35498 3223
rect 35536 3189 35570 3223
rect 35608 3189 35642 3223
rect 35680 3189 35714 3223
rect 35752 3189 35786 3223
rect 35824 3189 35858 3223
rect 35896 3189 35930 3223
rect 35968 3189 36002 3223
rect 36040 3189 36074 3223
rect 36112 3189 36146 3223
rect 36184 3189 36218 3223
rect 36256 3189 36290 3223
rect 36328 3189 36362 3223
rect 36400 3189 36434 3223
rect 36472 3189 36506 3223
rect 36544 3189 36578 3223
rect 36616 3189 36650 3223
rect 36688 3189 36722 3223
rect 36760 3189 36794 3223
rect 36832 3189 36866 3223
rect 36904 3189 36938 3223
rect 36976 3189 37010 3223
rect 37048 3189 37082 3223
rect 37120 3189 37154 3223
rect 37192 3189 37226 3223
rect 37264 3189 37298 3223
rect 37336 3189 37370 3223
rect 37408 3189 37442 3223
rect 37480 3189 37514 3223
rect 37552 3189 37586 3223
rect 37624 3189 37658 3223
rect 37696 3189 37730 3223
rect 37768 3189 37802 3223
rect 37840 3189 37874 3223
rect 37912 3189 37946 3223
rect 37984 3189 38018 3223
rect 38056 3189 38090 3223
rect 38128 3189 38162 3223
rect 38200 3189 38234 3223
rect 38272 3189 38306 3223
rect 38344 3189 38378 3223
rect 38416 3189 38450 3223
rect 38488 3189 38522 3223
rect 38560 3189 38594 3223
rect 29037 3066 29071 3100
rect 29037 2994 29071 3028
rect 29037 2922 29071 2956
rect 29037 2850 29071 2884
rect 29037 2778 29071 2812
rect 29037 2706 29071 2740
rect 29037 2634 29071 2668
rect 29037 2562 29071 2596
rect 29037 2490 29071 2524
rect 29037 2418 29071 2452
rect 29037 2346 29071 2380
rect 29037 2274 29071 2308
rect 29037 2202 29071 2236
rect 29037 2130 29071 2164
rect 29037 2058 29071 2092
rect 29037 1986 29071 2020
rect 29037 1914 29071 1948
rect 29037 1842 29071 1876
rect 29037 1770 29071 1804
rect 29037 1698 29071 1732
rect 29037 1626 29071 1660
rect 29037 1554 29071 1588
rect 29037 1482 29071 1516
rect 29037 1410 29071 1444
rect 29037 1338 29071 1372
rect 29037 1266 29071 1300
rect 29037 1194 29071 1228
rect 29133 3066 29167 3100
rect 29133 2994 29167 3028
rect 29133 2922 29167 2956
rect 29133 2850 29167 2884
rect 29133 2778 29167 2812
rect 29133 2706 29167 2740
rect 29133 2634 29167 2668
rect 29133 2562 29167 2596
rect 29133 2490 29167 2524
rect 29133 2418 29167 2452
rect 29133 2346 29167 2380
rect 29133 2274 29167 2308
rect 29133 2202 29167 2236
rect 29133 2130 29167 2164
rect 29133 2058 29167 2092
rect 29133 1986 29167 2020
rect 29133 1914 29167 1948
rect 29133 1842 29167 1876
rect 29133 1770 29167 1804
rect 29133 1698 29167 1732
rect 29133 1626 29167 1660
rect 29133 1554 29167 1588
rect 29133 1482 29167 1516
rect 29133 1410 29167 1444
rect 29133 1338 29167 1372
rect 29133 1266 29167 1300
rect 29133 1194 29167 1228
rect 29229 3066 29263 3100
rect 29229 2994 29263 3028
rect 29229 2922 29263 2956
rect 29229 2850 29263 2884
rect 29229 2778 29263 2812
rect 29229 2706 29263 2740
rect 29229 2634 29263 2668
rect 29229 2562 29263 2596
rect 29229 2490 29263 2524
rect 29229 2418 29263 2452
rect 29229 2346 29263 2380
rect 29229 2274 29263 2308
rect 29229 2202 29263 2236
rect 29229 2130 29263 2164
rect 29229 2058 29263 2092
rect 29229 1986 29263 2020
rect 29229 1914 29263 1948
rect 29229 1842 29263 1876
rect 29229 1770 29263 1804
rect 29229 1698 29263 1732
rect 29229 1626 29263 1660
rect 29229 1554 29263 1588
rect 29229 1482 29263 1516
rect 29229 1410 29263 1444
rect 29229 1338 29263 1372
rect 29229 1266 29263 1300
rect 29229 1194 29263 1228
rect 29325 3066 29359 3100
rect 29325 2994 29359 3028
rect 29325 2922 29359 2956
rect 29325 2850 29359 2884
rect 29325 2778 29359 2812
rect 29325 2706 29359 2740
rect 29325 2634 29359 2668
rect 29325 2562 29359 2596
rect 29325 2490 29359 2524
rect 29325 2418 29359 2452
rect 29325 2346 29359 2380
rect 29325 2274 29359 2308
rect 29325 2202 29359 2236
rect 29325 2130 29359 2164
rect 29325 2058 29359 2092
rect 29325 1986 29359 2020
rect 29325 1914 29359 1948
rect 29325 1842 29359 1876
rect 29325 1770 29359 1804
rect 29325 1698 29359 1732
rect 29325 1626 29359 1660
rect 29325 1554 29359 1588
rect 29325 1482 29359 1516
rect 29325 1410 29359 1444
rect 29325 1338 29359 1372
rect 29325 1266 29359 1300
rect 29325 1194 29359 1228
rect 29421 3066 29455 3100
rect 29421 2994 29455 3028
rect 29421 2922 29455 2956
rect 29421 2850 29455 2884
rect 29421 2778 29455 2812
rect 29421 2706 29455 2740
rect 29421 2634 29455 2668
rect 29421 2562 29455 2596
rect 29421 2490 29455 2524
rect 29421 2418 29455 2452
rect 29421 2346 29455 2380
rect 29421 2274 29455 2308
rect 29421 2202 29455 2236
rect 29421 2130 29455 2164
rect 29421 2058 29455 2092
rect 29421 1986 29455 2020
rect 29421 1914 29455 1948
rect 29421 1842 29455 1876
rect 29421 1770 29455 1804
rect 29421 1698 29455 1732
rect 29421 1626 29455 1660
rect 29421 1554 29455 1588
rect 29421 1482 29455 1516
rect 29421 1410 29455 1444
rect 29421 1338 29455 1372
rect 29421 1266 29455 1300
rect 29421 1194 29455 1228
rect 29517 3066 29551 3100
rect 29517 2994 29551 3028
rect 29517 2922 29551 2956
rect 29517 2850 29551 2884
rect 29517 2778 29551 2812
rect 29517 2706 29551 2740
rect 29517 2634 29551 2668
rect 29517 2562 29551 2596
rect 29517 2490 29551 2524
rect 29517 2418 29551 2452
rect 29517 2346 29551 2380
rect 29517 2274 29551 2308
rect 29517 2202 29551 2236
rect 29517 2130 29551 2164
rect 29517 2058 29551 2092
rect 29517 1986 29551 2020
rect 29517 1914 29551 1948
rect 29517 1842 29551 1876
rect 29517 1770 29551 1804
rect 29517 1698 29551 1732
rect 29517 1626 29551 1660
rect 29517 1554 29551 1588
rect 29517 1482 29551 1516
rect 29517 1410 29551 1444
rect 29517 1338 29551 1372
rect 29517 1266 29551 1300
rect 29517 1194 29551 1228
rect 29613 3066 29647 3100
rect 29613 2994 29647 3028
rect 29613 2922 29647 2956
rect 29613 2850 29647 2884
rect 29613 2778 29647 2812
rect 29613 2706 29647 2740
rect 29613 2634 29647 2668
rect 29613 2562 29647 2596
rect 29613 2490 29647 2524
rect 29613 2418 29647 2452
rect 29613 2346 29647 2380
rect 29613 2274 29647 2308
rect 29613 2202 29647 2236
rect 29613 2130 29647 2164
rect 29613 2058 29647 2092
rect 29613 1986 29647 2020
rect 29613 1914 29647 1948
rect 29613 1842 29647 1876
rect 29613 1770 29647 1804
rect 29613 1698 29647 1732
rect 29613 1626 29647 1660
rect 29613 1554 29647 1588
rect 29613 1482 29647 1516
rect 29613 1410 29647 1444
rect 29613 1338 29647 1372
rect 29613 1266 29647 1300
rect 29613 1194 29647 1228
rect 29709 3066 29743 3100
rect 29709 2994 29743 3028
rect 29709 2922 29743 2956
rect 29709 2850 29743 2884
rect 29709 2778 29743 2812
rect 29709 2706 29743 2740
rect 29709 2634 29743 2668
rect 29709 2562 29743 2596
rect 29709 2490 29743 2524
rect 29709 2418 29743 2452
rect 29709 2346 29743 2380
rect 29709 2274 29743 2308
rect 29709 2202 29743 2236
rect 29709 2130 29743 2164
rect 29709 2058 29743 2092
rect 29709 1986 29743 2020
rect 29709 1914 29743 1948
rect 29709 1842 29743 1876
rect 29709 1770 29743 1804
rect 29709 1698 29743 1732
rect 29709 1626 29743 1660
rect 29709 1554 29743 1588
rect 29709 1482 29743 1516
rect 29709 1410 29743 1444
rect 29709 1338 29743 1372
rect 29709 1266 29743 1300
rect 29709 1194 29743 1228
rect 29805 3066 29839 3100
rect 29805 2994 29839 3028
rect 29805 2922 29839 2956
rect 29805 2850 29839 2884
rect 29805 2778 29839 2812
rect 29805 2706 29839 2740
rect 29805 2634 29839 2668
rect 29805 2562 29839 2596
rect 29805 2490 29839 2524
rect 29805 2418 29839 2452
rect 29805 2346 29839 2380
rect 29805 2274 29839 2308
rect 29805 2202 29839 2236
rect 29805 2130 29839 2164
rect 29805 2058 29839 2092
rect 29805 1986 29839 2020
rect 29805 1914 29839 1948
rect 29805 1842 29839 1876
rect 29805 1770 29839 1804
rect 29805 1698 29839 1732
rect 29805 1626 29839 1660
rect 29805 1554 29839 1588
rect 29805 1482 29839 1516
rect 29805 1410 29839 1444
rect 29805 1338 29839 1372
rect 29805 1266 29839 1300
rect 29805 1194 29839 1228
rect 29901 3066 29935 3100
rect 29901 2994 29935 3028
rect 29901 2922 29935 2956
rect 29901 2850 29935 2884
rect 29901 2778 29935 2812
rect 29901 2706 29935 2740
rect 29901 2634 29935 2668
rect 29901 2562 29935 2596
rect 29901 2490 29935 2524
rect 29901 2418 29935 2452
rect 29901 2346 29935 2380
rect 29901 2274 29935 2308
rect 29901 2202 29935 2236
rect 29901 2130 29935 2164
rect 29901 2058 29935 2092
rect 29901 1986 29935 2020
rect 29901 1914 29935 1948
rect 29901 1842 29935 1876
rect 29901 1770 29935 1804
rect 29901 1698 29935 1732
rect 29901 1626 29935 1660
rect 29901 1554 29935 1588
rect 29901 1482 29935 1516
rect 29901 1410 29935 1444
rect 29901 1338 29935 1372
rect 29901 1266 29935 1300
rect 29901 1194 29935 1228
rect 29997 3066 30031 3100
rect 29997 2994 30031 3028
rect 29997 2922 30031 2956
rect 29997 2850 30031 2884
rect 29997 2778 30031 2812
rect 29997 2706 30031 2740
rect 29997 2634 30031 2668
rect 29997 2562 30031 2596
rect 29997 2490 30031 2524
rect 29997 2418 30031 2452
rect 29997 2346 30031 2380
rect 29997 2274 30031 2308
rect 29997 2202 30031 2236
rect 29997 2130 30031 2164
rect 29997 2058 30031 2092
rect 29997 1986 30031 2020
rect 29997 1914 30031 1948
rect 29997 1842 30031 1876
rect 29997 1770 30031 1804
rect 29997 1698 30031 1732
rect 29997 1626 30031 1660
rect 29997 1554 30031 1588
rect 29997 1482 30031 1516
rect 29997 1410 30031 1444
rect 29997 1338 30031 1372
rect 29997 1266 30031 1300
rect 29997 1194 30031 1228
rect 30093 3066 30127 3100
rect 30093 2994 30127 3028
rect 30093 2922 30127 2956
rect 30093 2850 30127 2884
rect 30093 2778 30127 2812
rect 30093 2706 30127 2740
rect 30093 2634 30127 2668
rect 30093 2562 30127 2596
rect 30093 2490 30127 2524
rect 30093 2418 30127 2452
rect 30093 2346 30127 2380
rect 30093 2274 30127 2308
rect 30093 2202 30127 2236
rect 30093 2130 30127 2164
rect 30093 2058 30127 2092
rect 30093 1986 30127 2020
rect 30093 1914 30127 1948
rect 30093 1842 30127 1876
rect 30093 1770 30127 1804
rect 30093 1698 30127 1732
rect 30093 1626 30127 1660
rect 30093 1554 30127 1588
rect 30093 1482 30127 1516
rect 30093 1410 30127 1444
rect 30093 1338 30127 1372
rect 30093 1266 30127 1300
rect 30093 1194 30127 1228
rect 30189 3066 30223 3100
rect 30189 2994 30223 3028
rect 30189 2922 30223 2956
rect 30189 2850 30223 2884
rect 30189 2778 30223 2812
rect 30189 2706 30223 2740
rect 30189 2634 30223 2668
rect 30189 2562 30223 2596
rect 30189 2490 30223 2524
rect 30189 2418 30223 2452
rect 30189 2346 30223 2380
rect 30189 2274 30223 2308
rect 30189 2202 30223 2236
rect 30189 2130 30223 2164
rect 30189 2058 30223 2092
rect 30189 1986 30223 2020
rect 30189 1914 30223 1948
rect 30189 1842 30223 1876
rect 30189 1770 30223 1804
rect 30189 1698 30223 1732
rect 30189 1626 30223 1660
rect 30189 1554 30223 1588
rect 30189 1482 30223 1516
rect 30189 1410 30223 1444
rect 30189 1338 30223 1372
rect 30189 1266 30223 1300
rect 30189 1194 30223 1228
rect 30285 3066 30319 3100
rect 30285 2994 30319 3028
rect 30285 2922 30319 2956
rect 30285 2850 30319 2884
rect 30285 2778 30319 2812
rect 30285 2706 30319 2740
rect 30285 2634 30319 2668
rect 30285 2562 30319 2596
rect 30285 2490 30319 2524
rect 30285 2418 30319 2452
rect 30285 2346 30319 2380
rect 30285 2274 30319 2308
rect 30285 2202 30319 2236
rect 30285 2130 30319 2164
rect 30285 2058 30319 2092
rect 30285 1986 30319 2020
rect 30285 1914 30319 1948
rect 30285 1842 30319 1876
rect 30285 1770 30319 1804
rect 30285 1698 30319 1732
rect 30285 1626 30319 1660
rect 30285 1554 30319 1588
rect 30285 1482 30319 1516
rect 30285 1410 30319 1444
rect 30285 1338 30319 1372
rect 30285 1266 30319 1300
rect 30285 1194 30319 1228
rect 30381 3066 30415 3100
rect 30381 2994 30415 3028
rect 30381 2922 30415 2956
rect 30381 2850 30415 2884
rect 30381 2778 30415 2812
rect 30381 2706 30415 2740
rect 30381 2634 30415 2668
rect 30381 2562 30415 2596
rect 30381 2490 30415 2524
rect 30381 2418 30415 2452
rect 30381 2346 30415 2380
rect 30381 2274 30415 2308
rect 30381 2202 30415 2236
rect 30381 2130 30415 2164
rect 30381 2058 30415 2092
rect 30381 1986 30415 2020
rect 30381 1914 30415 1948
rect 30381 1842 30415 1876
rect 30381 1770 30415 1804
rect 30381 1698 30415 1732
rect 30381 1626 30415 1660
rect 30381 1554 30415 1588
rect 30381 1482 30415 1516
rect 30381 1410 30415 1444
rect 30381 1338 30415 1372
rect 30381 1266 30415 1300
rect 30381 1194 30415 1228
rect 30477 3066 30511 3100
rect 30477 2994 30511 3028
rect 30477 2922 30511 2956
rect 30477 2850 30511 2884
rect 30477 2778 30511 2812
rect 30477 2706 30511 2740
rect 30477 2634 30511 2668
rect 30477 2562 30511 2596
rect 30477 2490 30511 2524
rect 30477 2418 30511 2452
rect 30477 2346 30511 2380
rect 30477 2274 30511 2308
rect 30477 2202 30511 2236
rect 30477 2130 30511 2164
rect 30477 2058 30511 2092
rect 30477 1986 30511 2020
rect 30477 1914 30511 1948
rect 30477 1842 30511 1876
rect 30477 1770 30511 1804
rect 30477 1698 30511 1732
rect 30477 1626 30511 1660
rect 30477 1554 30511 1588
rect 30477 1482 30511 1516
rect 30477 1410 30511 1444
rect 30477 1338 30511 1372
rect 30477 1266 30511 1300
rect 30477 1194 30511 1228
rect 30573 3066 30607 3100
rect 30573 2994 30607 3028
rect 30573 2922 30607 2956
rect 30573 2850 30607 2884
rect 30573 2778 30607 2812
rect 30573 2706 30607 2740
rect 30573 2634 30607 2668
rect 30573 2562 30607 2596
rect 30573 2490 30607 2524
rect 30573 2418 30607 2452
rect 30573 2346 30607 2380
rect 30573 2274 30607 2308
rect 30573 2202 30607 2236
rect 30573 2130 30607 2164
rect 30573 2058 30607 2092
rect 30573 1986 30607 2020
rect 30573 1914 30607 1948
rect 30573 1842 30607 1876
rect 30573 1770 30607 1804
rect 30573 1698 30607 1732
rect 30573 1626 30607 1660
rect 30573 1554 30607 1588
rect 30573 1482 30607 1516
rect 30573 1410 30607 1444
rect 30573 1338 30607 1372
rect 30573 1266 30607 1300
rect 30573 1194 30607 1228
rect 30669 3066 30703 3100
rect 30669 2994 30703 3028
rect 30669 2922 30703 2956
rect 30669 2850 30703 2884
rect 30669 2778 30703 2812
rect 30669 2706 30703 2740
rect 30669 2634 30703 2668
rect 30669 2562 30703 2596
rect 30669 2490 30703 2524
rect 30669 2418 30703 2452
rect 30669 2346 30703 2380
rect 30669 2274 30703 2308
rect 30669 2202 30703 2236
rect 30669 2130 30703 2164
rect 30669 2058 30703 2092
rect 30669 1986 30703 2020
rect 30669 1914 30703 1948
rect 30669 1842 30703 1876
rect 30669 1770 30703 1804
rect 30669 1698 30703 1732
rect 30669 1626 30703 1660
rect 30669 1554 30703 1588
rect 30669 1482 30703 1516
rect 30669 1410 30703 1444
rect 30669 1338 30703 1372
rect 30669 1266 30703 1300
rect 30669 1194 30703 1228
rect 30765 3066 30799 3100
rect 30765 2994 30799 3028
rect 30765 2922 30799 2956
rect 30765 2850 30799 2884
rect 30765 2778 30799 2812
rect 30765 2706 30799 2740
rect 30765 2634 30799 2668
rect 30765 2562 30799 2596
rect 30765 2490 30799 2524
rect 30765 2418 30799 2452
rect 30765 2346 30799 2380
rect 30765 2274 30799 2308
rect 30765 2202 30799 2236
rect 30765 2130 30799 2164
rect 30765 2058 30799 2092
rect 30765 1986 30799 2020
rect 30765 1914 30799 1948
rect 30765 1842 30799 1876
rect 30765 1770 30799 1804
rect 30765 1698 30799 1732
rect 30765 1626 30799 1660
rect 30765 1554 30799 1588
rect 30765 1482 30799 1516
rect 30765 1410 30799 1444
rect 30765 1338 30799 1372
rect 30765 1266 30799 1300
rect 30765 1194 30799 1228
rect 30861 3066 30895 3100
rect 30861 2994 30895 3028
rect 30861 2922 30895 2956
rect 30861 2850 30895 2884
rect 30861 2778 30895 2812
rect 30861 2706 30895 2740
rect 30861 2634 30895 2668
rect 30861 2562 30895 2596
rect 30861 2490 30895 2524
rect 30861 2418 30895 2452
rect 30861 2346 30895 2380
rect 30861 2274 30895 2308
rect 30861 2202 30895 2236
rect 30861 2130 30895 2164
rect 30861 2058 30895 2092
rect 30861 1986 30895 2020
rect 30861 1914 30895 1948
rect 30861 1842 30895 1876
rect 30861 1770 30895 1804
rect 30861 1698 30895 1732
rect 30861 1626 30895 1660
rect 30861 1554 30895 1588
rect 30861 1482 30895 1516
rect 30861 1410 30895 1444
rect 30861 1338 30895 1372
rect 30861 1266 30895 1300
rect 30861 1194 30895 1228
rect 30957 3066 30991 3100
rect 30957 2994 30991 3028
rect 30957 2922 30991 2956
rect 30957 2850 30991 2884
rect 30957 2778 30991 2812
rect 30957 2706 30991 2740
rect 30957 2634 30991 2668
rect 30957 2562 30991 2596
rect 30957 2490 30991 2524
rect 30957 2418 30991 2452
rect 30957 2346 30991 2380
rect 30957 2274 30991 2308
rect 30957 2202 30991 2236
rect 30957 2130 30991 2164
rect 30957 2058 30991 2092
rect 30957 1986 30991 2020
rect 30957 1914 30991 1948
rect 30957 1842 30991 1876
rect 30957 1770 30991 1804
rect 30957 1698 30991 1732
rect 30957 1626 30991 1660
rect 30957 1554 30991 1588
rect 30957 1482 30991 1516
rect 30957 1410 30991 1444
rect 30957 1338 30991 1372
rect 30957 1266 30991 1300
rect 30957 1194 30991 1228
rect 31053 3066 31087 3100
rect 31053 2994 31087 3028
rect 31053 2922 31087 2956
rect 31053 2850 31087 2884
rect 31053 2778 31087 2812
rect 31053 2706 31087 2740
rect 31053 2634 31087 2668
rect 31053 2562 31087 2596
rect 31053 2490 31087 2524
rect 31053 2418 31087 2452
rect 31053 2346 31087 2380
rect 31053 2274 31087 2308
rect 31053 2202 31087 2236
rect 31053 2130 31087 2164
rect 31053 2058 31087 2092
rect 31053 1986 31087 2020
rect 31053 1914 31087 1948
rect 31053 1842 31087 1876
rect 31053 1770 31087 1804
rect 31053 1698 31087 1732
rect 31053 1626 31087 1660
rect 31053 1554 31087 1588
rect 31053 1482 31087 1516
rect 31053 1410 31087 1444
rect 31053 1338 31087 1372
rect 31053 1266 31087 1300
rect 31053 1194 31087 1228
rect 31149 3066 31183 3100
rect 31149 2994 31183 3028
rect 31149 2922 31183 2956
rect 31149 2850 31183 2884
rect 31149 2778 31183 2812
rect 31149 2706 31183 2740
rect 31149 2634 31183 2668
rect 31149 2562 31183 2596
rect 31149 2490 31183 2524
rect 31149 2418 31183 2452
rect 31149 2346 31183 2380
rect 31149 2274 31183 2308
rect 31149 2202 31183 2236
rect 31149 2130 31183 2164
rect 31149 2058 31183 2092
rect 31149 1986 31183 2020
rect 31149 1914 31183 1948
rect 31149 1842 31183 1876
rect 31149 1770 31183 1804
rect 31149 1698 31183 1732
rect 31149 1626 31183 1660
rect 31149 1554 31183 1588
rect 31149 1482 31183 1516
rect 31149 1410 31183 1444
rect 31149 1338 31183 1372
rect 31149 1266 31183 1300
rect 31149 1194 31183 1228
rect 31245 3066 31279 3100
rect 31245 2994 31279 3028
rect 31245 2922 31279 2956
rect 31245 2850 31279 2884
rect 31245 2778 31279 2812
rect 31245 2706 31279 2740
rect 31245 2634 31279 2668
rect 31245 2562 31279 2596
rect 31245 2490 31279 2524
rect 31245 2418 31279 2452
rect 31245 2346 31279 2380
rect 31245 2274 31279 2308
rect 31245 2202 31279 2236
rect 31245 2130 31279 2164
rect 31245 2058 31279 2092
rect 31245 1986 31279 2020
rect 31245 1914 31279 1948
rect 31245 1842 31279 1876
rect 31245 1770 31279 1804
rect 31245 1698 31279 1732
rect 31245 1626 31279 1660
rect 31245 1554 31279 1588
rect 31245 1482 31279 1516
rect 31245 1410 31279 1444
rect 31245 1338 31279 1372
rect 31245 1266 31279 1300
rect 31245 1194 31279 1228
rect 31341 3066 31375 3100
rect 31341 2994 31375 3028
rect 31341 2922 31375 2956
rect 31341 2850 31375 2884
rect 31341 2778 31375 2812
rect 31341 2706 31375 2740
rect 31341 2634 31375 2668
rect 31341 2562 31375 2596
rect 31341 2490 31375 2524
rect 31341 2418 31375 2452
rect 31341 2346 31375 2380
rect 31341 2274 31375 2308
rect 31341 2202 31375 2236
rect 31341 2130 31375 2164
rect 31341 2058 31375 2092
rect 31341 1986 31375 2020
rect 31341 1914 31375 1948
rect 31341 1842 31375 1876
rect 31341 1770 31375 1804
rect 31341 1698 31375 1732
rect 31341 1626 31375 1660
rect 31341 1554 31375 1588
rect 31341 1482 31375 1516
rect 31341 1410 31375 1444
rect 31341 1338 31375 1372
rect 31341 1266 31375 1300
rect 31341 1194 31375 1228
rect 31437 3066 31471 3100
rect 31437 2994 31471 3028
rect 31437 2922 31471 2956
rect 31437 2850 31471 2884
rect 31437 2778 31471 2812
rect 31437 2706 31471 2740
rect 31437 2634 31471 2668
rect 31437 2562 31471 2596
rect 31437 2490 31471 2524
rect 31437 2418 31471 2452
rect 31437 2346 31471 2380
rect 31437 2274 31471 2308
rect 31437 2202 31471 2236
rect 31437 2130 31471 2164
rect 31437 2058 31471 2092
rect 31437 1986 31471 2020
rect 31437 1914 31471 1948
rect 31437 1842 31471 1876
rect 31437 1770 31471 1804
rect 31437 1698 31471 1732
rect 31437 1626 31471 1660
rect 31437 1554 31471 1588
rect 31437 1482 31471 1516
rect 31437 1410 31471 1444
rect 31437 1338 31471 1372
rect 31437 1266 31471 1300
rect 31437 1194 31471 1228
rect 31533 3066 31567 3100
rect 31533 2994 31567 3028
rect 31533 2922 31567 2956
rect 31533 2850 31567 2884
rect 31533 2778 31567 2812
rect 31533 2706 31567 2740
rect 31533 2634 31567 2668
rect 31533 2562 31567 2596
rect 31533 2490 31567 2524
rect 31533 2418 31567 2452
rect 31533 2346 31567 2380
rect 31533 2274 31567 2308
rect 31533 2202 31567 2236
rect 31533 2130 31567 2164
rect 31533 2058 31567 2092
rect 31533 1986 31567 2020
rect 31533 1914 31567 1948
rect 31533 1842 31567 1876
rect 31533 1770 31567 1804
rect 31533 1698 31567 1732
rect 31533 1626 31567 1660
rect 31533 1554 31567 1588
rect 31533 1482 31567 1516
rect 31533 1410 31567 1444
rect 31533 1338 31567 1372
rect 31533 1266 31567 1300
rect 31533 1194 31567 1228
rect 31629 3066 31663 3100
rect 31629 2994 31663 3028
rect 31629 2922 31663 2956
rect 31629 2850 31663 2884
rect 31629 2778 31663 2812
rect 31629 2706 31663 2740
rect 31629 2634 31663 2668
rect 31629 2562 31663 2596
rect 31629 2490 31663 2524
rect 31629 2418 31663 2452
rect 31629 2346 31663 2380
rect 31629 2274 31663 2308
rect 31629 2202 31663 2236
rect 31629 2130 31663 2164
rect 31629 2058 31663 2092
rect 31629 1986 31663 2020
rect 31629 1914 31663 1948
rect 31629 1842 31663 1876
rect 31629 1770 31663 1804
rect 31629 1698 31663 1732
rect 31629 1626 31663 1660
rect 31629 1554 31663 1588
rect 31629 1482 31663 1516
rect 31629 1410 31663 1444
rect 31629 1338 31663 1372
rect 31629 1266 31663 1300
rect 31629 1194 31663 1228
rect 31725 3066 31759 3100
rect 31725 2994 31759 3028
rect 31725 2922 31759 2956
rect 31725 2850 31759 2884
rect 31725 2778 31759 2812
rect 31725 2706 31759 2740
rect 31725 2634 31759 2668
rect 31725 2562 31759 2596
rect 31725 2490 31759 2524
rect 31725 2418 31759 2452
rect 31725 2346 31759 2380
rect 31725 2274 31759 2308
rect 31725 2202 31759 2236
rect 31725 2130 31759 2164
rect 31725 2058 31759 2092
rect 31725 1986 31759 2020
rect 31725 1914 31759 1948
rect 31725 1842 31759 1876
rect 31725 1770 31759 1804
rect 31725 1698 31759 1732
rect 31725 1626 31759 1660
rect 31725 1554 31759 1588
rect 31725 1482 31759 1516
rect 31725 1410 31759 1444
rect 31725 1338 31759 1372
rect 31725 1266 31759 1300
rect 31725 1194 31759 1228
rect 31821 3066 31855 3100
rect 31821 2994 31855 3028
rect 31821 2922 31855 2956
rect 31821 2850 31855 2884
rect 31821 2778 31855 2812
rect 31821 2706 31855 2740
rect 31821 2634 31855 2668
rect 31821 2562 31855 2596
rect 31821 2490 31855 2524
rect 31821 2418 31855 2452
rect 31821 2346 31855 2380
rect 31821 2274 31855 2308
rect 31821 2202 31855 2236
rect 31821 2130 31855 2164
rect 31821 2058 31855 2092
rect 31821 1986 31855 2020
rect 31821 1914 31855 1948
rect 31821 1842 31855 1876
rect 31821 1770 31855 1804
rect 31821 1698 31855 1732
rect 31821 1626 31855 1660
rect 31821 1554 31855 1588
rect 31821 1482 31855 1516
rect 31821 1410 31855 1444
rect 31821 1338 31855 1372
rect 31821 1266 31855 1300
rect 31821 1194 31855 1228
rect 31917 3066 31951 3100
rect 31917 2994 31951 3028
rect 31917 2922 31951 2956
rect 31917 2850 31951 2884
rect 31917 2778 31951 2812
rect 31917 2706 31951 2740
rect 31917 2634 31951 2668
rect 31917 2562 31951 2596
rect 31917 2490 31951 2524
rect 31917 2418 31951 2452
rect 31917 2346 31951 2380
rect 31917 2274 31951 2308
rect 31917 2202 31951 2236
rect 31917 2130 31951 2164
rect 31917 2058 31951 2092
rect 31917 1986 31951 2020
rect 31917 1914 31951 1948
rect 31917 1842 31951 1876
rect 31917 1770 31951 1804
rect 31917 1698 31951 1732
rect 31917 1626 31951 1660
rect 31917 1554 31951 1588
rect 31917 1482 31951 1516
rect 31917 1410 31951 1444
rect 31917 1338 31951 1372
rect 31917 1266 31951 1300
rect 31917 1194 31951 1228
rect 32013 3066 32047 3100
rect 32013 2994 32047 3028
rect 32013 2922 32047 2956
rect 32013 2850 32047 2884
rect 32013 2778 32047 2812
rect 32013 2706 32047 2740
rect 32013 2634 32047 2668
rect 32013 2562 32047 2596
rect 32013 2490 32047 2524
rect 32013 2418 32047 2452
rect 32013 2346 32047 2380
rect 32013 2274 32047 2308
rect 32013 2202 32047 2236
rect 32013 2130 32047 2164
rect 32013 2058 32047 2092
rect 32013 1986 32047 2020
rect 32013 1914 32047 1948
rect 32013 1842 32047 1876
rect 32013 1770 32047 1804
rect 32013 1698 32047 1732
rect 32013 1626 32047 1660
rect 32013 1554 32047 1588
rect 32013 1482 32047 1516
rect 32013 1410 32047 1444
rect 32013 1338 32047 1372
rect 32013 1266 32047 1300
rect 32013 1194 32047 1228
rect 32109 3066 32143 3100
rect 32109 2994 32143 3028
rect 32109 2922 32143 2956
rect 32109 2850 32143 2884
rect 32109 2778 32143 2812
rect 32109 2706 32143 2740
rect 32109 2634 32143 2668
rect 32109 2562 32143 2596
rect 32109 2490 32143 2524
rect 32109 2418 32143 2452
rect 32109 2346 32143 2380
rect 32109 2274 32143 2308
rect 32109 2202 32143 2236
rect 32109 2130 32143 2164
rect 32109 2058 32143 2092
rect 32109 1986 32143 2020
rect 32109 1914 32143 1948
rect 32109 1842 32143 1876
rect 32109 1770 32143 1804
rect 32109 1698 32143 1732
rect 32109 1626 32143 1660
rect 32109 1554 32143 1588
rect 32109 1482 32143 1516
rect 32109 1410 32143 1444
rect 32109 1338 32143 1372
rect 32109 1266 32143 1300
rect 32109 1194 32143 1228
rect 32205 3066 32239 3100
rect 32205 2994 32239 3028
rect 32205 2922 32239 2956
rect 32205 2850 32239 2884
rect 32205 2778 32239 2812
rect 32205 2706 32239 2740
rect 32205 2634 32239 2668
rect 32205 2562 32239 2596
rect 32205 2490 32239 2524
rect 32205 2418 32239 2452
rect 32205 2346 32239 2380
rect 32205 2274 32239 2308
rect 32205 2202 32239 2236
rect 32205 2130 32239 2164
rect 32205 2058 32239 2092
rect 32205 1986 32239 2020
rect 32205 1914 32239 1948
rect 32205 1842 32239 1876
rect 32205 1770 32239 1804
rect 32205 1698 32239 1732
rect 32205 1626 32239 1660
rect 32205 1554 32239 1588
rect 32205 1482 32239 1516
rect 32205 1410 32239 1444
rect 32205 1338 32239 1372
rect 32205 1266 32239 1300
rect 32205 1194 32239 1228
rect 32301 3066 32335 3100
rect 32301 2994 32335 3028
rect 32301 2922 32335 2956
rect 32301 2850 32335 2884
rect 32301 2778 32335 2812
rect 32301 2706 32335 2740
rect 32301 2634 32335 2668
rect 32301 2562 32335 2596
rect 32301 2490 32335 2524
rect 32301 2418 32335 2452
rect 32301 2346 32335 2380
rect 32301 2274 32335 2308
rect 32301 2202 32335 2236
rect 32301 2130 32335 2164
rect 32301 2058 32335 2092
rect 32301 1986 32335 2020
rect 32301 1914 32335 1948
rect 32301 1842 32335 1876
rect 32301 1770 32335 1804
rect 32301 1698 32335 1732
rect 32301 1626 32335 1660
rect 32301 1554 32335 1588
rect 32301 1482 32335 1516
rect 32301 1410 32335 1444
rect 32301 1338 32335 1372
rect 32301 1266 32335 1300
rect 32301 1194 32335 1228
rect 32397 3066 32431 3100
rect 32397 2994 32431 3028
rect 32397 2922 32431 2956
rect 32397 2850 32431 2884
rect 32397 2778 32431 2812
rect 32397 2706 32431 2740
rect 32397 2634 32431 2668
rect 32397 2562 32431 2596
rect 32397 2490 32431 2524
rect 32397 2418 32431 2452
rect 32397 2346 32431 2380
rect 32397 2274 32431 2308
rect 32397 2202 32431 2236
rect 32397 2130 32431 2164
rect 32397 2058 32431 2092
rect 32397 1986 32431 2020
rect 32397 1914 32431 1948
rect 32397 1842 32431 1876
rect 32397 1770 32431 1804
rect 32397 1698 32431 1732
rect 32397 1626 32431 1660
rect 32397 1554 32431 1588
rect 32397 1482 32431 1516
rect 32397 1410 32431 1444
rect 32397 1338 32431 1372
rect 32397 1266 32431 1300
rect 32397 1194 32431 1228
rect 32493 3066 32527 3100
rect 32493 2994 32527 3028
rect 32493 2922 32527 2956
rect 32493 2850 32527 2884
rect 32493 2778 32527 2812
rect 32493 2706 32527 2740
rect 32493 2634 32527 2668
rect 32493 2562 32527 2596
rect 32493 2490 32527 2524
rect 32493 2418 32527 2452
rect 32493 2346 32527 2380
rect 32493 2274 32527 2308
rect 32493 2202 32527 2236
rect 32493 2130 32527 2164
rect 32493 2058 32527 2092
rect 32493 1986 32527 2020
rect 32493 1914 32527 1948
rect 32493 1842 32527 1876
rect 32493 1770 32527 1804
rect 32493 1698 32527 1732
rect 32493 1626 32527 1660
rect 32493 1554 32527 1588
rect 32493 1482 32527 1516
rect 32493 1410 32527 1444
rect 32493 1338 32527 1372
rect 32493 1266 32527 1300
rect 32493 1194 32527 1228
rect 32589 3066 32623 3100
rect 32589 2994 32623 3028
rect 32589 2922 32623 2956
rect 32589 2850 32623 2884
rect 32589 2778 32623 2812
rect 32589 2706 32623 2740
rect 32589 2634 32623 2668
rect 32589 2562 32623 2596
rect 32589 2490 32623 2524
rect 32589 2418 32623 2452
rect 32589 2346 32623 2380
rect 32589 2274 32623 2308
rect 32589 2202 32623 2236
rect 32589 2130 32623 2164
rect 32589 2058 32623 2092
rect 32589 1986 32623 2020
rect 32589 1914 32623 1948
rect 32589 1842 32623 1876
rect 32589 1770 32623 1804
rect 32589 1698 32623 1732
rect 32589 1626 32623 1660
rect 32589 1554 32623 1588
rect 32589 1482 32623 1516
rect 32589 1410 32623 1444
rect 32589 1338 32623 1372
rect 32589 1266 32623 1300
rect 32589 1194 32623 1228
rect 32685 3066 32719 3100
rect 32685 2994 32719 3028
rect 32685 2922 32719 2956
rect 32685 2850 32719 2884
rect 32685 2778 32719 2812
rect 32685 2706 32719 2740
rect 32685 2634 32719 2668
rect 32685 2562 32719 2596
rect 32685 2490 32719 2524
rect 32685 2418 32719 2452
rect 32685 2346 32719 2380
rect 32685 2274 32719 2308
rect 32685 2202 32719 2236
rect 32685 2130 32719 2164
rect 32685 2058 32719 2092
rect 32685 1986 32719 2020
rect 32685 1914 32719 1948
rect 32685 1842 32719 1876
rect 32685 1770 32719 1804
rect 32685 1698 32719 1732
rect 32685 1626 32719 1660
rect 32685 1554 32719 1588
rect 32685 1482 32719 1516
rect 32685 1410 32719 1444
rect 32685 1338 32719 1372
rect 32685 1266 32719 1300
rect 32685 1194 32719 1228
rect 32781 3066 32815 3100
rect 32781 2994 32815 3028
rect 32781 2922 32815 2956
rect 32781 2850 32815 2884
rect 32781 2778 32815 2812
rect 32781 2706 32815 2740
rect 32781 2634 32815 2668
rect 32781 2562 32815 2596
rect 32781 2490 32815 2524
rect 32781 2418 32815 2452
rect 32781 2346 32815 2380
rect 32781 2274 32815 2308
rect 32781 2202 32815 2236
rect 32781 2130 32815 2164
rect 32781 2058 32815 2092
rect 32781 1986 32815 2020
rect 32781 1914 32815 1948
rect 32781 1842 32815 1876
rect 32781 1770 32815 1804
rect 32781 1698 32815 1732
rect 32781 1626 32815 1660
rect 32781 1554 32815 1588
rect 32781 1482 32815 1516
rect 32781 1410 32815 1444
rect 32781 1338 32815 1372
rect 32781 1266 32815 1300
rect 32781 1194 32815 1228
rect 32877 3066 32911 3100
rect 32877 2994 32911 3028
rect 32877 2922 32911 2956
rect 32877 2850 32911 2884
rect 32877 2778 32911 2812
rect 32877 2706 32911 2740
rect 32877 2634 32911 2668
rect 32877 2562 32911 2596
rect 32877 2490 32911 2524
rect 32877 2418 32911 2452
rect 32877 2346 32911 2380
rect 32877 2274 32911 2308
rect 32877 2202 32911 2236
rect 32877 2130 32911 2164
rect 32877 2058 32911 2092
rect 32877 1986 32911 2020
rect 32877 1914 32911 1948
rect 32877 1842 32911 1876
rect 32877 1770 32911 1804
rect 32877 1698 32911 1732
rect 32877 1626 32911 1660
rect 32877 1554 32911 1588
rect 32877 1482 32911 1516
rect 32877 1410 32911 1444
rect 32877 1338 32911 1372
rect 32877 1266 32911 1300
rect 32877 1194 32911 1228
rect 32973 3066 33007 3100
rect 32973 2994 33007 3028
rect 32973 2922 33007 2956
rect 32973 2850 33007 2884
rect 32973 2778 33007 2812
rect 32973 2706 33007 2740
rect 32973 2634 33007 2668
rect 32973 2562 33007 2596
rect 32973 2490 33007 2524
rect 32973 2418 33007 2452
rect 32973 2346 33007 2380
rect 32973 2274 33007 2308
rect 32973 2202 33007 2236
rect 32973 2130 33007 2164
rect 32973 2058 33007 2092
rect 32973 1986 33007 2020
rect 32973 1914 33007 1948
rect 32973 1842 33007 1876
rect 32973 1770 33007 1804
rect 32973 1698 33007 1732
rect 32973 1626 33007 1660
rect 32973 1554 33007 1588
rect 32973 1482 33007 1516
rect 32973 1410 33007 1444
rect 32973 1338 33007 1372
rect 32973 1266 33007 1300
rect 32973 1194 33007 1228
rect 33069 3066 33103 3100
rect 33069 2994 33103 3028
rect 33069 2922 33103 2956
rect 33069 2850 33103 2884
rect 33069 2778 33103 2812
rect 33069 2706 33103 2740
rect 33069 2634 33103 2668
rect 33069 2562 33103 2596
rect 33069 2490 33103 2524
rect 33069 2418 33103 2452
rect 33069 2346 33103 2380
rect 33069 2274 33103 2308
rect 33069 2202 33103 2236
rect 33069 2130 33103 2164
rect 33069 2058 33103 2092
rect 33069 1986 33103 2020
rect 33069 1914 33103 1948
rect 33069 1842 33103 1876
rect 33069 1770 33103 1804
rect 33069 1698 33103 1732
rect 33069 1626 33103 1660
rect 33069 1554 33103 1588
rect 33069 1482 33103 1516
rect 33069 1410 33103 1444
rect 33069 1338 33103 1372
rect 33069 1266 33103 1300
rect 33069 1194 33103 1228
rect 33165 3066 33199 3100
rect 33165 2994 33199 3028
rect 33165 2922 33199 2956
rect 33165 2850 33199 2884
rect 33165 2778 33199 2812
rect 33165 2706 33199 2740
rect 33165 2634 33199 2668
rect 33165 2562 33199 2596
rect 33165 2490 33199 2524
rect 33165 2418 33199 2452
rect 33165 2346 33199 2380
rect 33165 2274 33199 2308
rect 33165 2202 33199 2236
rect 33165 2130 33199 2164
rect 33165 2058 33199 2092
rect 33165 1986 33199 2020
rect 33165 1914 33199 1948
rect 33165 1842 33199 1876
rect 33165 1770 33199 1804
rect 33165 1698 33199 1732
rect 33165 1626 33199 1660
rect 33165 1554 33199 1588
rect 33165 1482 33199 1516
rect 33165 1410 33199 1444
rect 33165 1338 33199 1372
rect 33165 1266 33199 1300
rect 33165 1194 33199 1228
rect 33261 3066 33295 3100
rect 33261 2994 33295 3028
rect 33261 2922 33295 2956
rect 33261 2850 33295 2884
rect 33261 2778 33295 2812
rect 33261 2706 33295 2740
rect 33261 2634 33295 2668
rect 33261 2562 33295 2596
rect 33261 2490 33295 2524
rect 33261 2418 33295 2452
rect 33261 2346 33295 2380
rect 33261 2274 33295 2308
rect 33261 2202 33295 2236
rect 33261 2130 33295 2164
rect 33261 2058 33295 2092
rect 33261 1986 33295 2020
rect 33261 1914 33295 1948
rect 33261 1842 33295 1876
rect 33261 1770 33295 1804
rect 33261 1698 33295 1732
rect 33261 1626 33295 1660
rect 33261 1554 33295 1588
rect 33261 1482 33295 1516
rect 33261 1410 33295 1444
rect 33261 1338 33295 1372
rect 33261 1266 33295 1300
rect 33261 1194 33295 1228
rect 33357 3066 33391 3100
rect 33357 2994 33391 3028
rect 33357 2922 33391 2956
rect 33357 2850 33391 2884
rect 33357 2778 33391 2812
rect 33357 2706 33391 2740
rect 33357 2634 33391 2668
rect 33357 2562 33391 2596
rect 33357 2490 33391 2524
rect 33357 2418 33391 2452
rect 33357 2346 33391 2380
rect 33357 2274 33391 2308
rect 33357 2202 33391 2236
rect 33357 2130 33391 2164
rect 33357 2058 33391 2092
rect 33357 1986 33391 2020
rect 33357 1914 33391 1948
rect 33357 1842 33391 1876
rect 33357 1770 33391 1804
rect 33357 1698 33391 1732
rect 33357 1626 33391 1660
rect 33357 1554 33391 1588
rect 33357 1482 33391 1516
rect 33357 1410 33391 1444
rect 33357 1338 33391 1372
rect 33357 1266 33391 1300
rect 33357 1194 33391 1228
rect 33453 3066 33487 3100
rect 33453 2994 33487 3028
rect 33453 2922 33487 2956
rect 33453 2850 33487 2884
rect 33453 2778 33487 2812
rect 33453 2706 33487 2740
rect 33453 2634 33487 2668
rect 33453 2562 33487 2596
rect 33453 2490 33487 2524
rect 33453 2418 33487 2452
rect 33453 2346 33487 2380
rect 33453 2274 33487 2308
rect 33453 2202 33487 2236
rect 33453 2130 33487 2164
rect 33453 2058 33487 2092
rect 33453 1986 33487 2020
rect 33453 1914 33487 1948
rect 33453 1842 33487 1876
rect 33453 1770 33487 1804
rect 33453 1698 33487 1732
rect 33453 1626 33487 1660
rect 33453 1554 33487 1588
rect 33453 1482 33487 1516
rect 33453 1410 33487 1444
rect 33453 1338 33487 1372
rect 33453 1266 33487 1300
rect 33453 1194 33487 1228
rect 33549 3066 33583 3100
rect 33549 2994 33583 3028
rect 33549 2922 33583 2956
rect 33549 2850 33583 2884
rect 33549 2778 33583 2812
rect 33549 2706 33583 2740
rect 33549 2634 33583 2668
rect 33549 2562 33583 2596
rect 33549 2490 33583 2524
rect 33549 2418 33583 2452
rect 33549 2346 33583 2380
rect 33549 2274 33583 2308
rect 33549 2202 33583 2236
rect 33549 2130 33583 2164
rect 33549 2058 33583 2092
rect 33549 1986 33583 2020
rect 33549 1914 33583 1948
rect 33549 1842 33583 1876
rect 33549 1770 33583 1804
rect 33549 1698 33583 1732
rect 33549 1626 33583 1660
rect 33549 1554 33583 1588
rect 33549 1482 33583 1516
rect 33549 1410 33583 1444
rect 33549 1338 33583 1372
rect 33549 1266 33583 1300
rect 33549 1194 33583 1228
rect 33645 3066 33679 3100
rect 33645 2994 33679 3028
rect 33645 2922 33679 2956
rect 33645 2850 33679 2884
rect 33645 2778 33679 2812
rect 33645 2706 33679 2740
rect 33645 2634 33679 2668
rect 33645 2562 33679 2596
rect 33645 2490 33679 2524
rect 33645 2418 33679 2452
rect 33645 2346 33679 2380
rect 33645 2274 33679 2308
rect 33645 2202 33679 2236
rect 33645 2130 33679 2164
rect 33645 2058 33679 2092
rect 33645 1986 33679 2020
rect 33645 1914 33679 1948
rect 33645 1842 33679 1876
rect 33645 1770 33679 1804
rect 33645 1698 33679 1732
rect 33645 1626 33679 1660
rect 33645 1554 33679 1588
rect 33645 1482 33679 1516
rect 33645 1410 33679 1444
rect 33645 1338 33679 1372
rect 33645 1266 33679 1300
rect 33645 1194 33679 1228
rect 33741 3066 33775 3100
rect 33741 2994 33775 3028
rect 33741 2922 33775 2956
rect 33741 2850 33775 2884
rect 33741 2778 33775 2812
rect 33741 2706 33775 2740
rect 33741 2634 33775 2668
rect 33741 2562 33775 2596
rect 33741 2490 33775 2524
rect 33741 2418 33775 2452
rect 33741 2346 33775 2380
rect 33741 2274 33775 2308
rect 33741 2202 33775 2236
rect 33741 2130 33775 2164
rect 33741 2058 33775 2092
rect 33741 1986 33775 2020
rect 33741 1914 33775 1948
rect 33741 1842 33775 1876
rect 33741 1770 33775 1804
rect 33741 1698 33775 1732
rect 33741 1626 33775 1660
rect 33741 1554 33775 1588
rect 33741 1482 33775 1516
rect 33741 1410 33775 1444
rect 33741 1338 33775 1372
rect 33741 1266 33775 1300
rect 33741 1194 33775 1228
rect 33837 3066 33871 3100
rect 33837 2994 33871 3028
rect 33837 2922 33871 2956
rect 33837 2850 33871 2884
rect 33837 2778 33871 2812
rect 33837 2706 33871 2740
rect 33837 2634 33871 2668
rect 33837 2562 33871 2596
rect 33837 2490 33871 2524
rect 33837 2418 33871 2452
rect 33837 2346 33871 2380
rect 33837 2274 33871 2308
rect 33837 2202 33871 2236
rect 33837 2130 33871 2164
rect 33837 2058 33871 2092
rect 33837 1986 33871 2020
rect 33837 1914 33871 1948
rect 33837 1842 33871 1876
rect 33837 1770 33871 1804
rect 33837 1698 33871 1732
rect 33837 1626 33871 1660
rect 33837 1554 33871 1588
rect 33837 1482 33871 1516
rect 33837 1410 33871 1444
rect 33837 1338 33871 1372
rect 33837 1266 33871 1300
rect 33837 1194 33871 1228
rect 33933 3066 33967 3100
rect 33933 2994 33967 3028
rect 33933 2922 33967 2956
rect 33933 2850 33967 2884
rect 33933 2778 33967 2812
rect 33933 2706 33967 2740
rect 33933 2634 33967 2668
rect 33933 2562 33967 2596
rect 33933 2490 33967 2524
rect 33933 2418 33967 2452
rect 33933 2346 33967 2380
rect 33933 2274 33967 2308
rect 33933 2202 33967 2236
rect 33933 2130 33967 2164
rect 33933 2058 33967 2092
rect 33933 1986 33967 2020
rect 33933 1914 33967 1948
rect 33933 1842 33967 1876
rect 33933 1770 33967 1804
rect 33933 1698 33967 1732
rect 33933 1626 33967 1660
rect 33933 1554 33967 1588
rect 33933 1482 33967 1516
rect 33933 1410 33967 1444
rect 33933 1338 33967 1372
rect 33933 1266 33967 1300
rect 33933 1194 33967 1228
rect 34029 3066 34063 3100
rect 34029 2994 34063 3028
rect 34029 2922 34063 2956
rect 34029 2850 34063 2884
rect 34029 2778 34063 2812
rect 34029 2706 34063 2740
rect 34029 2634 34063 2668
rect 34029 2562 34063 2596
rect 34029 2490 34063 2524
rect 34029 2418 34063 2452
rect 34029 2346 34063 2380
rect 34029 2274 34063 2308
rect 34029 2202 34063 2236
rect 34029 2130 34063 2164
rect 34029 2058 34063 2092
rect 34029 1986 34063 2020
rect 34029 1914 34063 1948
rect 34029 1842 34063 1876
rect 34029 1770 34063 1804
rect 34029 1698 34063 1732
rect 34029 1626 34063 1660
rect 34029 1554 34063 1588
rect 34029 1482 34063 1516
rect 34029 1410 34063 1444
rect 34029 1338 34063 1372
rect 34029 1266 34063 1300
rect 34029 1194 34063 1228
rect 34125 3066 34159 3100
rect 34125 2994 34159 3028
rect 34125 2922 34159 2956
rect 34125 2850 34159 2884
rect 34125 2778 34159 2812
rect 34125 2706 34159 2740
rect 34125 2634 34159 2668
rect 34125 2562 34159 2596
rect 34125 2490 34159 2524
rect 34125 2418 34159 2452
rect 34125 2346 34159 2380
rect 34125 2274 34159 2308
rect 34125 2202 34159 2236
rect 34125 2130 34159 2164
rect 34125 2058 34159 2092
rect 34125 1986 34159 2020
rect 34125 1914 34159 1948
rect 34125 1842 34159 1876
rect 34125 1770 34159 1804
rect 34125 1698 34159 1732
rect 34125 1626 34159 1660
rect 34125 1554 34159 1588
rect 34125 1482 34159 1516
rect 34125 1410 34159 1444
rect 34125 1338 34159 1372
rect 34125 1266 34159 1300
rect 34125 1194 34159 1228
rect 34221 3066 34255 3100
rect 34221 2994 34255 3028
rect 34221 2922 34255 2956
rect 34221 2850 34255 2884
rect 34221 2778 34255 2812
rect 34221 2706 34255 2740
rect 34221 2634 34255 2668
rect 34221 2562 34255 2596
rect 34221 2490 34255 2524
rect 34221 2418 34255 2452
rect 34221 2346 34255 2380
rect 34221 2274 34255 2308
rect 34221 2202 34255 2236
rect 34221 2130 34255 2164
rect 34221 2058 34255 2092
rect 34221 1986 34255 2020
rect 34221 1914 34255 1948
rect 34221 1842 34255 1876
rect 34221 1770 34255 1804
rect 34221 1698 34255 1732
rect 34221 1626 34255 1660
rect 34221 1554 34255 1588
rect 34221 1482 34255 1516
rect 34221 1410 34255 1444
rect 34221 1338 34255 1372
rect 34221 1266 34255 1300
rect 34221 1194 34255 1228
rect 34317 3066 34351 3100
rect 34317 2994 34351 3028
rect 34317 2922 34351 2956
rect 34317 2850 34351 2884
rect 34317 2778 34351 2812
rect 34317 2706 34351 2740
rect 34317 2634 34351 2668
rect 34317 2562 34351 2596
rect 34317 2490 34351 2524
rect 34317 2418 34351 2452
rect 34317 2346 34351 2380
rect 34317 2274 34351 2308
rect 34317 2202 34351 2236
rect 34317 2130 34351 2164
rect 34317 2058 34351 2092
rect 34317 1986 34351 2020
rect 34317 1914 34351 1948
rect 34317 1842 34351 1876
rect 34317 1770 34351 1804
rect 34317 1698 34351 1732
rect 34317 1626 34351 1660
rect 34317 1554 34351 1588
rect 34317 1482 34351 1516
rect 34317 1410 34351 1444
rect 34317 1338 34351 1372
rect 34317 1266 34351 1300
rect 34317 1194 34351 1228
rect 34413 3066 34447 3100
rect 34413 2994 34447 3028
rect 34413 2922 34447 2956
rect 34413 2850 34447 2884
rect 34413 2778 34447 2812
rect 34413 2706 34447 2740
rect 34413 2634 34447 2668
rect 34413 2562 34447 2596
rect 34413 2490 34447 2524
rect 34413 2418 34447 2452
rect 34413 2346 34447 2380
rect 34413 2274 34447 2308
rect 34413 2202 34447 2236
rect 34413 2130 34447 2164
rect 34413 2058 34447 2092
rect 34413 1986 34447 2020
rect 34413 1914 34447 1948
rect 34413 1842 34447 1876
rect 34413 1770 34447 1804
rect 34413 1698 34447 1732
rect 34413 1626 34447 1660
rect 34413 1554 34447 1588
rect 34413 1482 34447 1516
rect 34413 1410 34447 1444
rect 34413 1338 34447 1372
rect 34413 1266 34447 1300
rect 34413 1194 34447 1228
rect 34509 3066 34543 3100
rect 34509 2994 34543 3028
rect 34509 2922 34543 2956
rect 34509 2850 34543 2884
rect 34509 2778 34543 2812
rect 34509 2706 34543 2740
rect 34509 2634 34543 2668
rect 34509 2562 34543 2596
rect 34509 2490 34543 2524
rect 34509 2418 34543 2452
rect 34509 2346 34543 2380
rect 34509 2274 34543 2308
rect 34509 2202 34543 2236
rect 34509 2130 34543 2164
rect 34509 2058 34543 2092
rect 34509 1986 34543 2020
rect 34509 1914 34543 1948
rect 34509 1842 34543 1876
rect 34509 1770 34543 1804
rect 34509 1698 34543 1732
rect 34509 1626 34543 1660
rect 34509 1554 34543 1588
rect 34509 1482 34543 1516
rect 34509 1410 34543 1444
rect 34509 1338 34543 1372
rect 34509 1266 34543 1300
rect 34509 1194 34543 1228
rect 34605 3066 34639 3100
rect 34605 2994 34639 3028
rect 34605 2922 34639 2956
rect 34605 2850 34639 2884
rect 34605 2778 34639 2812
rect 34605 2706 34639 2740
rect 34605 2634 34639 2668
rect 34605 2562 34639 2596
rect 34605 2490 34639 2524
rect 34605 2418 34639 2452
rect 34605 2346 34639 2380
rect 34605 2274 34639 2308
rect 34605 2202 34639 2236
rect 34605 2130 34639 2164
rect 34605 2058 34639 2092
rect 34605 1986 34639 2020
rect 34605 1914 34639 1948
rect 34605 1842 34639 1876
rect 34605 1770 34639 1804
rect 34605 1698 34639 1732
rect 34605 1626 34639 1660
rect 34605 1554 34639 1588
rect 34605 1482 34639 1516
rect 34605 1410 34639 1444
rect 34605 1338 34639 1372
rect 34605 1266 34639 1300
rect 34605 1194 34639 1228
rect 34701 3066 34735 3100
rect 34701 2994 34735 3028
rect 34701 2922 34735 2956
rect 34701 2850 34735 2884
rect 34701 2778 34735 2812
rect 34701 2706 34735 2740
rect 34701 2634 34735 2668
rect 34701 2562 34735 2596
rect 34701 2490 34735 2524
rect 34701 2418 34735 2452
rect 34701 2346 34735 2380
rect 34701 2274 34735 2308
rect 34701 2202 34735 2236
rect 34701 2130 34735 2164
rect 34701 2058 34735 2092
rect 34701 1986 34735 2020
rect 34701 1914 34735 1948
rect 34701 1842 34735 1876
rect 34701 1770 34735 1804
rect 34701 1698 34735 1732
rect 34701 1626 34735 1660
rect 34701 1554 34735 1588
rect 34701 1482 34735 1516
rect 34701 1410 34735 1444
rect 34701 1338 34735 1372
rect 34701 1266 34735 1300
rect 34701 1194 34735 1228
rect 34797 3066 34831 3100
rect 34797 2994 34831 3028
rect 34797 2922 34831 2956
rect 34797 2850 34831 2884
rect 34797 2778 34831 2812
rect 34797 2706 34831 2740
rect 34797 2634 34831 2668
rect 34797 2562 34831 2596
rect 34797 2490 34831 2524
rect 34797 2418 34831 2452
rect 34797 2346 34831 2380
rect 34797 2274 34831 2308
rect 34797 2202 34831 2236
rect 34797 2130 34831 2164
rect 34797 2058 34831 2092
rect 34797 1986 34831 2020
rect 34797 1914 34831 1948
rect 34797 1842 34831 1876
rect 34797 1770 34831 1804
rect 34797 1698 34831 1732
rect 34797 1626 34831 1660
rect 34797 1554 34831 1588
rect 34797 1482 34831 1516
rect 34797 1410 34831 1444
rect 34797 1338 34831 1372
rect 34797 1266 34831 1300
rect 34797 1194 34831 1228
rect 34893 3066 34927 3100
rect 34893 2994 34927 3028
rect 34893 2922 34927 2956
rect 34893 2850 34927 2884
rect 34893 2778 34927 2812
rect 34893 2706 34927 2740
rect 34893 2634 34927 2668
rect 34893 2562 34927 2596
rect 34893 2490 34927 2524
rect 34893 2418 34927 2452
rect 34893 2346 34927 2380
rect 34893 2274 34927 2308
rect 34893 2202 34927 2236
rect 34893 2130 34927 2164
rect 34893 2058 34927 2092
rect 34893 1986 34927 2020
rect 34893 1914 34927 1948
rect 34893 1842 34927 1876
rect 34893 1770 34927 1804
rect 34893 1698 34927 1732
rect 34893 1626 34927 1660
rect 34893 1554 34927 1588
rect 34893 1482 34927 1516
rect 34893 1410 34927 1444
rect 34893 1338 34927 1372
rect 34893 1266 34927 1300
rect 34893 1194 34927 1228
rect 34989 3066 35023 3100
rect 34989 2994 35023 3028
rect 34989 2922 35023 2956
rect 34989 2850 35023 2884
rect 34989 2778 35023 2812
rect 34989 2706 35023 2740
rect 34989 2634 35023 2668
rect 34989 2562 35023 2596
rect 34989 2490 35023 2524
rect 34989 2418 35023 2452
rect 34989 2346 35023 2380
rect 34989 2274 35023 2308
rect 34989 2202 35023 2236
rect 34989 2130 35023 2164
rect 34989 2058 35023 2092
rect 34989 1986 35023 2020
rect 34989 1914 35023 1948
rect 34989 1842 35023 1876
rect 34989 1770 35023 1804
rect 34989 1698 35023 1732
rect 34989 1626 35023 1660
rect 34989 1554 35023 1588
rect 34989 1482 35023 1516
rect 34989 1410 35023 1444
rect 34989 1338 35023 1372
rect 34989 1266 35023 1300
rect 34989 1194 35023 1228
rect 35085 3066 35119 3100
rect 35085 2994 35119 3028
rect 35085 2922 35119 2956
rect 35085 2850 35119 2884
rect 35085 2778 35119 2812
rect 35085 2706 35119 2740
rect 35085 2634 35119 2668
rect 35085 2562 35119 2596
rect 35085 2490 35119 2524
rect 35085 2418 35119 2452
rect 35085 2346 35119 2380
rect 35085 2274 35119 2308
rect 35085 2202 35119 2236
rect 35085 2130 35119 2164
rect 35085 2058 35119 2092
rect 35085 1986 35119 2020
rect 35085 1914 35119 1948
rect 35085 1842 35119 1876
rect 35085 1770 35119 1804
rect 35085 1698 35119 1732
rect 35085 1626 35119 1660
rect 35085 1554 35119 1588
rect 35085 1482 35119 1516
rect 35085 1410 35119 1444
rect 35085 1338 35119 1372
rect 35085 1266 35119 1300
rect 35085 1194 35119 1228
rect 35181 3066 35215 3100
rect 35181 2994 35215 3028
rect 35181 2922 35215 2956
rect 35181 2850 35215 2884
rect 35181 2778 35215 2812
rect 35181 2706 35215 2740
rect 35181 2634 35215 2668
rect 35181 2562 35215 2596
rect 35181 2490 35215 2524
rect 35181 2418 35215 2452
rect 35181 2346 35215 2380
rect 35181 2274 35215 2308
rect 35181 2202 35215 2236
rect 35181 2130 35215 2164
rect 35181 2058 35215 2092
rect 35181 1986 35215 2020
rect 35181 1914 35215 1948
rect 35181 1842 35215 1876
rect 35181 1770 35215 1804
rect 35181 1698 35215 1732
rect 35181 1626 35215 1660
rect 35181 1554 35215 1588
rect 35181 1482 35215 1516
rect 35181 1410 35215 1444
rect 35181 1338 35215 1372
rect 35181 1266 35215 1300
rect 35181 1194 35215 1228
rect 35277 3066 35311 3100
rect 35277 2994 35311 3028
rect 35277 2922 35311 2956
rect 35277 2850 35311 2884
rect 35277 2778 35311 2812
rect 35277 2706 35311 2740
rect 35277 2634 35311 2668
rect 35277 2562 35311 2596
rect 35277 2490 35311 2524
rect 35277 2418 35311 2452
rect 35277 2346 35311 2380
rect 35277 2274 35311 2308
rect 35277 2202 35311 2236
rect 35277 2130 35311 2164
rect 35277 2058 35311 2092
rect 35277 1986 35311 2020
rect 35277 1914 35311 1948
rect 35277 1842 35311 1876
rect 35277 1770 35311 1804
rect 35277 1698 35311 1732
rect 35277 1626 35311 1660
rect 35277 1554 35311 1588
rect 35277 1482 35311 1516
rect 35277 1410 35311 1444
rect 35277 1338 35311 1372
rect 35277 1266 35311 1300
rect 35277 1194 35311 1228
rect 35373 3066 35407 3100
rect 35373 2994 35407 3028
rect 35373 2922 35407 2956
rect 35373 2850 35407 2884
rect 35373 2778 35407 2812
rect 35373 2706 35407 2740
rect 35373 2634 35407 2668
rect 35373 2562 35407 2596
rect 35373 2490 35407 2524
rect 35373 2418 35407 2452
rect 35373 2346 35407 2380
rect 35373 2274 35407 2308
rect 35373 2202 35407 2236
rect 35373 2130 35407 2164
rect 35373 2058 35407 2092
rect 35373 1986 35407 2020
rect 35373 1914 35407 1948
rect 35373 1842 35407 1876
rect 35373 1770 35407 1804
rect 35373 1698 35407 1732
rect 35373 1626 35407 1660
rect 35373 1554 35407 1588
rect 35373 1482 35407 1516
rect 35373 1410 35407 1444
rect 35373 1338 35407 1372
rect 35373 1266 35407 1300
rect 35373 1194 35407 1228
rect 35469 3066 35503 3100
rect 35469 2994 35503 3028
rect 35469 2922 35503 2956
rect 35469 2850 35503 2884
rect 35469 2778 35503 2812
rect 35469 2706 35503 2740
rect 35469 2634 35503 2668
rect 35469 2562 35503 2596
rect 35469 2490 35503 2524
rect 35469 2418 35503 2452
rect 35469 2346 35503 2380
rect 35469 2274 35503 2308
rect 35469 2202 35503 2236
rect 35469 2130 35503 2164
rect 35469 2058 35503 2092
rect 35469 1986 35503 2020
rect 35469 1914 35503 1948
rect 35469 1842 35503 1876
rect 35469 1770 35503 1804
rect 35469 1698 35503 1732
rect 35469 1626 35503 1660
rect 35469 1554 35503 1588
rect 35469 1482 35503 1516
rect 35469 1410 35503 1444
rect 35469 1338 35503 1372
rect 35469 1266 35503 1300
rect 35469 1194 35503 1228
rect 35565 3066 35599 3100
rect 35565 2994 35599 3028
rect 35565 2922 35599 2956
rect 35565 2850 35599 2884
rect 35565 2778 35599 2812
rect 35565 2706 35599 2740
rect 35565 2634 35599 2668
rect 35565 2562 35599 2596
rect 35565 2490 35599 2524
rect 35565 2418 35599 2452
rect 35565 2346 35599 2380
rect 35565 2274 35599 2308
rect 35565 2202 35599 2236
rect 35565 2130 35599 2164
rect 35565 2058 35599 2092
rect 35565 1986 35599 2020
rect 35565 1914 35599 1948
rect 35565 1842 35599 1876
rect 35565 1770 35599 1804
rect 35565 1698 35599 1732
rect 35565 1626 35599 1660
rect 35565 1554 35599 1588
rect 35565 1482 35599 1516
rect 35565 1410 35599 1444
rect 35565 1338 35599 1372
rect 35565 1266 35599 1300
rect 35565 1194 35599 1228
rect 35661 3066 35695 3100
rect 35661 2994 35695 3028
rect 35661 2922 35695 2956
rect 35661 2850 35695 2884
rect 35661 2778 35695 2812
rect 35661 2706 35695 2740
rect 35661 2634 35695 2668
rect 35661 2562 35695 2596
rect 35661 2490 35695 2524
rect 35661 2418 35695 2452
rect 35661 2346 35695 2380
rect 35661 2274 35695 2308
rect 35661 2202 35695 2236
rect 35661 2130 35695 2164
rect 35661 2058 35695 2092
rect 35661 1986 35695 2020
rect 35661 1914 35695 1948
rect 35661 1842 35695 1876
rect 35661 1770 35695 1804
rect 35661 1698 35695 1732
rect 35661 1626 35695 1660
rect 35661 1554 35695 1588
rect 35661 1482 35695 1516
rect 35661 1410 35695 1444
rect 35661 1338 35695 1372
rect 35661 1266 35695 1300
rect 35661 1194 35695 1228
rect 35757 3066 35791 3100
rect 35757 2994 35791 3028
rect 35757 2922 35791 2956
rect 35757 2850 35791 2884
rect 35757 2778 35791 2812
rect 35757 2706 35791 2740
rect 35757 2634 35791 2668
rect 35757 2562 35791 2596
rect 35757 2490 35791 2524
rect 35757 2418 35791 2452
rect 35757 2346 35791 2380
rect 35757 2274 35791 2308
rect 35757 2202 35791 2236
rect 35757 2130 35791 2164
rect 35757 2058 35791 2092
rect 35757 1986 35791 2020
rect 35757 1914 35791 1948
rect 35757 1842 35791 1876
rect 35757 1770 35791 1804
rect 35757 1698 35791 1732
rect 35757 1626 35791 1660
rect 35757 1554 35791 1588
rect 35757 1482 35791 1516
rect 35757 1410 35791 1444
rect 35757 1338 35791 1372
rect 35757 1266 35791 1300
rect 35757 1194 35791 1228
rect 35853 3066 35887 3100
rect 35853 2994 35887 3028
rect 35853 2922 35887 2956
rect 35853 2850 35887 2884
rect 35853 2778 35887 2812
rect 35853 2706 35887 2740
rect 35853 2634 35887 2668
rect 35853 2562 35887 2596
rect 35853 2490 35887 2524
rect 35853 2418 35887 2452
rect 35853 2346 35887 2380
rect 35853 2274 35887 2308
rect 35853 2202 35887 2236
rect 35853 2130 35887 2164
rect 35853 2058 35887 2092
rect 35853 1986 35887 2020
rect 35853 1914 35887 1948
rect 35853 1842 35887 1876
rect 35853 1770 35887 1804
rect 35853 1698 35887 1732
rect 35853 1626 35887 1660
rect 35853 1554 35887 1588
rect 35853 1482 35887 1516
rect 35853 1410 35887 1444
rect 35853 1338 35887 1372
rect 35853 1266 35887 1300
rect 35853 1194 35887 1228
rect 35949 3066 35983 3100
rect 35949 2994 35983 3028
rect 35949 2922 35983 2956
rect 35949 2850 35983 2884
rect 35949 2778 35983 2812
rect 35949 2706 35983 2740
rect 35949 2634 35983 2668
rect 35949 2562 35983 2596
rect 35949 2490 35983 2524
rect 35949 2418 35983 2452
rect 35949 2346 35983 2380
rect 35949 2274 35983 2308
rect 35949 2202 35983 2236
rect 35949 2130 35983 2164
rect 35949 2058 35983 2092
rect 35949 1986 35983 2020
rect 35949 1914 35983 1948
rect 35949 1842 35983 1876
rect 35949 1770 35983 1804
rect 35949 1698 35983 1732
rect 35949 1626 35983 1660
rect 35949 1554 35983 1588
rect 35949 1482 35983 1516
rect 35949 1410 35983 1444
rect 35949 1338 35983 1372
rect 35949 1266 35983 1300
rect 35949 1194 35983 1228
rect 36045 3066 36079 3100
rect 36045 2994 36079 3028
rect 36045 2922 36079 2956
rect 36045 2850 36079 2884
rect 36045 2778 36079 2812
rect 36045 2706 36079 2740
rect 36045 2634 36079 2668
rect 36045 2562 36079 2596
rect 36045 2490 36079 2524
rect 36045 2418 36079 2452
rect 36045 2346 36079 2380
rect 36045 2274 36079 2308
rect 36045 2202 36079 2236
rect 36045 2130 36079 2164
rect 36045 2058 36079 2092
rect 36045 1986 36079 2020
rect 36045 1914 36079 1948
rect 36045 1842 36079 1876
rect 36045 1770 36079 1804
rect 36045 1698 36079 1732
rect 36045 1626 36079 1660
rect 36045 1554 36079 1588
rect 36045 1482 36079 1516
rect 36045 1410 36079 1444
rect 36045 1338 36079 1372
rect 36045 1266 36079 1300
rect 36045 1194 36079 1228
rect 36141 3066 36175 3100
rect 36141 2994 36175 3028
rect 36141 2922 36175 2956
rect 36141 2850 36175 2884
rect 36141 2778 36175 2812
rect 36141 2706 36175 2740
rect 36141 2634 36175 2668
rect 36141 2562 36175 2596
rect 36141 2490 36175 2524
rect 36141 2418 36175 2452
rect 36141 2346 36175 2380
rect 36141 2274 36175 2308
rect 36141 2202 36175 2236
rect 36141 2130 36175 2164
rect 36141 2058 36175 2092
rect 36141 1986 36175 2020
rect 36141 1914 36175 1948
rect 36141 1842 36175 1876
rect 36141 1770 36175 1804
rect 36141 1698 36175 1732
rect 36141 1626 36175 1660
rect 36141 1554 36175 1588
rect 36141 1482 36175 1516
rect 36141 1410 36175 1444
rect 36141 1338 36175 1372
rect 36141 1266 36175 1300
rect 36141 1194 36175 1228
rect 36237 3066 36271 3100
rect 36237 2994 36271 3028
rect 36237 2922 36271 2956
rect 36237 2850 36271 2884
rect 36237 2778 36271 2812
rect 36237 2706 36271 2740
rect 36237 2634 36271 2668
rect 36237 2562 36271 2596
rect 36237 2490 36271 2524
rect 36237 2418 36271 2452
rect 36237 2346 36271 2380
rect 36237 2274 36271 2308
rect 36237 2202 36271 2236
rect 36237 2130 36271 2164
rect 36237 2058 36271 2092
rect 36237 1986 36271 2020
rect 36237 1914 36271 1948
rect 36237 1842 36271 1876
rect 36237 1770 36271 1804
rect 36237 1698 36271 1732
rect 36237 1626 36271 1660
rect 36237 1554 36271 1588
rect 36237 1482 36271 1516
rect 36237 1410 36271 1444
rect 36237 1338 36271 1372
rect 36237 1266 36271 1300
rect 36237 1194 36271 1228
rect 36333 3066 36367 3100
rect 36333 2994 36367 3028
rect 36333 2922 36367 2956
rect 36333 2850 36367 2884
rect 36333 2778 36367 2812
rect 36333 2706 36367 2740
rect 36333 2634 36367 2668
rect 36333 2562 36367 2596
rect 36333 2490 36367 2524
rect 36333 2418 36367 2452
rect 36333 2346 36367 2380
rect 36333 2274 36367 2308
rect 36333 2202 36367 2236
rect 36333 2130 36367 2164
rect 36333 2058 36367 2092
rect 36333 1986 36367 2020
rect 36333 1914 36367 1948
rect 36333 1842 36367 1876
rect 36333 1770 36367 1804
rect 36333 1698 36367 1732
rect 36333 1626 36367 1660
rect 36333 1554 36367 1588
rect 36333 1482 36367 1516
rect 36333 1410 36367 1444
rect 36333 1338 36367 1372
rect 36333 1266 36367 1300
rect 36333 1194 36367 1228
rect 36429 3066 36463 3100
rect 36429 2994 36463 3028
rect 36429 2922 36463 2956
rect 36429 2850 36463 2884
rect 36429 2778 36463 2812
rect 36429 2706 36463 2740
rect 36429 2634 36463 2668
rect 36429 2562 36463 2596
rect 36429 2490 36463 2524
rect 36429 2418 36463 2452
rect 36429 2346 36463 2380
rect 36429 2274 36463 2308
rect 36429 2202 36463 2236
rect 36429 2130 36463 2164
rect 36429 2058 36463 2092
rect 36429 1986 36463 2020
rect 36429 1914 36463 1948
rect 36429 1842 36463 1876
rect 36429 1770 36463 1804
rect 36429 1698 36463 1732
rect 36429 1626 36463 1660
rect 36429 1554 36463 1588
rect 36429 1482 36463 1516
rect 36429 1410 36463 1444
rect 36429 1338 36463 1372
rect 36429 1266 36463 1300
rect 36429 1194 36463 1228
rect 36525 3066 36559 3100
rect 36525 2994 36559 3028
rect 36525 2922 36559 2956
rect 36525 2850 36559 2884
rect 36525 2778 36559 2812
rect 36525 2706 36559 2740
rect 36525 2634 36559 2668
rect 36525 2562 36559 2596
rect 36525 2490 36559 2524
rect 36525 2418 36559 2452
rect 36525 2346 36559 2380
rect 36525 2274 36559 2308
rect 36525 2202 36559 2236
rect 36525 2130 36559 2164
rect 36525 2058 36559 2092
rect 36525 1986 36559 2020
rect 36525 1914 36559 1948
rect 36525 1842 36559 1876
rect 36525 1770 36559 1804
rect 36525 1698 36559 1732
rect 36525 1626 36559 1660
rect 36525 1554 36559 1588
rect 36525 1482 36559 1516
rect 36525 1410 36559 1444
rect 36525 1338 36559 1372
rect 36525 1266 36559 1300
rect 36525 1194 36559 1228
rect 36621 3066 36655 3100
rect 36621 2994 36655 3028
rect 36621 2922 36655 2956
rect 36621 2850 36655 2884
rect 36621 2778 36655 2812
rect 36621 2706 36655 2740
rect 36621 2634 36655 2668
rect 36621 2562 36655 2596
rect 36621 2490 36655 2524
rect 36621 2418 36655 2452
rect 36621 2346 36655 2380
rect 36621 2274 36655 2308
rect 36621 2202 36655 2236
rect 36621 2130 36655 2164
rect 36621 2058 36655 2092
rect 36621 1986 36655 2020
rect 36621 1914 36655 1948
rect 36621 1842 36655 1876
rect 36621 1770 36655 1804
rect 36621 1698 36655 1732
rect 36621 1626 36655 1660
rect 36621 1554 36655 1588
rect 36621 1482 36655 1516
rect 36621 1410 36655 1444
rect 36621 1338 36655 1372
rect 36621 1266 36655 1300
rect 36621 1194 36655 1228
rect 36717 3066 36751 3100
rect 36717 2994 36751 3028
rect 36717 2922 36751 2956
rect 36717 2850 36751 2884
rect 36717 2778 36751 2812
rect 36717 2706 36751 2740
rect 36717 2634 36751 2668
rect 36717 2562 36751 2596
rect 36717 2490 36751 2524
rect 36717 2418 36751 2452
rect 36717 2346 36751 2380
rect 36717 2274 36751 2308
rect 36717 2202 36751 2236
rect 36717 2130 36751 2164
rect 36717 2058 36751 2092
rect 36717 1986 36751 2020
rect 36717 1914 36751 1948
rect 36717 1842 36751 1876
rect 36717 1770 36751 1804
rect 36717 1698 36751 1732
rect 36717 1626 36751 1660
rect 36717 1554 36751 1588
rect 36717 1482 36751 1516
rect 36717 1410 36751 1444
rect 36717 1338 36751 1372
rect 36717 1266 36751 1300
rect 36717 1194 36751 1228
rect 36813 3066 36847 3100
rect 36813 2994 36847 3028
rect 36813 2922 36847 2956
rect 36813 2850 36847 2884
rect 36813 2778 36847 2812
rect 36813 2706 36847 2740
rect 36813 2634 36847 2668
rect 36813 2562 36847 2596
rect 36813 2490 36847 2524
rect 36813 2418 36847 2452
rect 36813 2346 36847 2380
rect 36813 2274 36847 2308
rect 36813 2202 36847 2236
rect 36813 2130 36847 2164
rect 36813 2058 36847 2092
rect 36813 1986 36847 2020
rect 36813 1914 36847 1948
rect 36813 1842 36847 1876
rect 36813 1770 36847 1804
rect 36813 1698 36847 1732
rect 36813 1626 36847 1660
rect 36813 1554 36847 1588
rect 36813 1482 36847 1516
rect 36813 1410 36847 1444
rect 36813 1338 36847 1372
rect 36813 1266 36847 1300
rect 36813 1194 36847 1228
rect 36909 3066 36943 3100
rect 36909 2994 36943 3028
rect 36909 2922 36943 2956
rect 36909 2850 36943 2884
rect 36909 2778 36943 2812
rect 36909 2706 36943 2740
rect 36909 2634 36943 2668
rect 36909 2562 36943 2596
rect 36909 2490 36943 2524
rect 36909 2418 36943 2452
rect 36909 2346 36943 2380
rect 36909 2274 36943 2308
rect 36909 2202 36943 2236
rect 36909 2130 36943 2164
rect 36909 2058 36943 2092
rect 36909 1986 36943 2020
rect 36909 1914 36943 1948
rect 36909 1842 36943 1876
rect 36909 1770 36943 1804
rect 36909 1698 36943 1732
rect 36909 1626 36943 1660
rect 36909 1554 36943 1588
rect 36909 1482 36943 1516
rect 36909 1410 36943 1444
rect 36909 1338 36943 1372
rect 36909 1266 36943 1300
rect 36909 1194 36943 1228
rect 37005 3066 37039 3100
rect 37005 2994 37039 3028
rect 37005 2922 37039 2956
rect 37005 2850 37039 2884
rect 37005 2778 37039 2812
rect 37005 2706 37039 2740
rect 37005 2634 37039 2668
rect 37005 2562 37039 2596
rect 37005 2490 37039 2524
rect 37005 2418 37039 2452
rect 37005 2346 37039 2380
rect 37005 2274 37039 2308
rect 37005 2202 37039 2236
rect 37005 2130 37039 2164
rect 37005 2058 37039 2092
rect 37005 1986 37039 2020
rect 37005 1914 37039 1948
rect 37005 1842 37039 1876
rect 37005 1770 37039 1804
rect 37005 1698 37039 1732
rect 37005 1626 37039 1660
rect 37005 1554 37039 1588
rect 37005 1482 37039 1516
rect 37005 1410 37039 1444
rect 37005 1338 37039 1372
rect 37005 1266 37039 1300
rect 37005 1194 37039 1228
rect 37101 3066 37135 3100
rect 37101 2994 37135 3028
rect 37101 2922 37135 2956
rect 37101 2850 37135 2884
rect 37101 2778 37135 2812
rect 37101 2706 37135 2740
rect 37101 2634 37135 2668
rect 37101 2562 37135 2596
rect 37101 2490 37135 2524
rect 37101 2418 37135 2452
rect 37101 2346 37135 2380
rect 37101 2274 37135 2308
rect 37101 2202 37135 2236
rect 37101 2130 37135 2164
rect 37101 2058 37135 2092
rect 37101 1986 37135 2020
rect 37101 1914 37135 1948
rect 37101 1842 37135 1876
rect 37101 1770 37135 1804
rect 37101 1698 37135 1732
rect 37101 1626 37135 1660
rect 37101 1554 37135 1588
rect 37101 1482 37135 1516
rect 37101 1410 37135 1444
rect 37101 1338 37135 1372
rect 37101 1266 37135 1300
rect 37101 1194 37135 1228
rect 37197 3066 37231 3100
rect 37197 2994 37231 3028
rect 37197 2922 37231 2956
rect 37197 2850 37231 2884
rect 37197 2778 37231 2812
rect 37197 2706 37231 2740
rect 37197 2634 37231 2668
rect 37197 2562 37231 2596
rect 37197 2490 37231 2524
rect 37197 2418 37231 2452
rect 37197 2346 37231 2380
rect 37197 2274 37231 2308
rect 37197 2202 37231 2236
rect 37197 2130 37231 2164
rect 37197 2058 37231 2092
rect 37197 1986 37231 2020
rect 37197 1914 37231 1948
rect 37197 1842 37231 1876
rect 37197 1770 37231 1804
rect 37197 1698 37231 1732
rect 37197 1626 37231 1660
rect 37197 1554 37231 1588
rect 37197 1482 37231 1516
rect 37197 1410 37231 1444
rect 37197 1338 37231 1372
rect 37197 1266 37231 1300
rect 37197 1194 37231 1228
rect 37293 3066 37327 3100
rect 37293 2994 37327 3028
rect 37293 2922 37327 2956
rect 37293 2850 37327 2884
rect 37293 2778 37327 2812
rect 37293 2706 37327 2740
rect 37293 2634 37327 2668
rect 37293 2562 37327 2596
rect 37293 2490 37327 2524
rect 37293 2418 37327 2452
rect 37293 2346 37327 2380
rect 37293 2274 37327 2308
rect 37293 2202 37327 2236
rect 37293 2130 37327 2164
rect 37293 2058 37327 2092
rect 37293 1986 37327 2020
rect 37293 1914 37327 1948
rect 37293 1842 37327 1876
rect 37293 1770 37327 1804
rect 37293 1698 37327 1732
rect 37293 1626 37327 1660
rect 37293 1554 37327 1588
rect 37293 1482 37327 1516
rect 37293 1410 37327 1444
rect 37293 1338 37327 1372
rect 37293 1266 37327 1300
rect 37293 1194 37327 1228
rect 37389 3066 37423 3100
rect 37389 2994 37423 3028
rect 37389 2922 37423 2956
rect 37389 2850 37423 2884
rect 37389 2778 37423 2812
rect 37389 2706 37423 2740
rect 37389 2634 37423 2668
rect 37389 2562 37423 2596
rect 37389 2490 37423 2524
rect 37389 2418 37423 2452
rect 37389 2346 37423 2380
rect 37389 2274 37423 2308
rect 37389 2202 37423 2236
rect 37389 2130 37423 2164
rect 37389 2058 37423 2092
rect 37389 1986 37423 2020
rect 37389 1914 37423 1948
rect 37389 1842 37423 1876
rect 37389 1770 37423 1804
rect 37389 1698 37423 1732
rect 37389 1626 37423 1660
rect 37389 1554 37423 1588
rect 37389 1482 37423 1516
rect 37389 1410 37423 1444
rect 37389 1338 37423 1372
rect 37389 1266 37423 1300
rect 37389 1194 37423 1228
rect 37485 3066 37519 3100
rect 37485 2994 37519 3028
rect 37485 2922 37519 2956
rect 37485 2850 37519 2884
rect 37485 2778 37519 2812
rect 37485 2706 37519 2740
rect 37485 2634 37519 2668
rect 37485 2562 37519 2596
rect 37485 2490 37519 2524
rect 37485 2418 37519 2452
rect 37485 2346 37519 2380
rect 37485 2274 37519 2308
rect 37485 2202 37519 2236
rect 37485 2130 37519 2164
rect 37485 2058 37519 2092
rect 37485 1986 37519 2020
rect 37485 1914 37519 1948
rect 37485 1842 37519 1876
rect 37485 1770 37519 1804
rect 37485 1698 37519 1732
rect 37485 1626 37519 1660
rect 37485 1554 37519 1588
rect 37485 1482 37519 1516
rect 37485 1410 37519 1444
rect 37485 1338 37519 1372
rect 37485 1266 37519 1300
rect 37485 1194 37519 1228
rect 37581 3066 37615 3100
rect 37581 2994 37615 3028
rect 37581 2922 37615 2956
rect 37581 2850 37615 2884
rect 37581 2778 37615 2812
rect 37581 2706 37615 2740
rect 37581 2634 37615 2668
rect 37581 2562 37615 2596
rect 37581 2490 37615 2524
rect 37581 2418 37615 2452
rect 37581 2346 37615 2380
rect 37581 2274 37615 2308
rect 37581 2202 37615 2236
rect 37581 2130 37615 2164
rect 37581 2058 37615 2092
rect 37581 1986 37615 2020
rect 37581 1914 37615 1948
rect 37581 1842 37615 1876
rect 37581 1770 37615 1804
rect 37581 1698 37615 1732
rect 37581 1626 37615 1660
rect 37581 1554 37615 1588
rect 37581 1482 37615 1516
rect 37581 1410 37615 1444
rect 37581 1338 37615 1372
rect 37581 1266 37615 1300
rect 37581 1194 37615 1228
rect 37677 3066 37711 3100
rect 37677 2994 37711 3028
rect 37677 2922 37711 2956
rect 37677 2850 37711 2884
rect 37677 2778 37711 2812
rect 37677 2706 37711 2740
rect 37677 2634 37711 2668
rect 37677 2562 37711 2596
rect 37677 2490 37711 2524
rect 37677 2418 37711 2452
rect 37677 2346 37711 2380
rect 37677 2274 37711 2308
rect 37677 2202 37711 2236
rect 37677 2130 37711 2164
rect 37677 2058 37711 2092
rect 37677 1986 37711 2020
rect 37677 1914 37711 1948
rect 37677 1842 37711 1876
rect 37677 1770 37711 1804
rect 37677 1698 37711 1732
rect 37677 1626 37711 1660
rect 37677 1554 37711 1588
rect 37677 1482 37711 1516
rect 37677 1410 37711 1444
rect 37677 1338 37711 1372
rect 37677 1266 37711 1300
rect 37677 1194 37711 1228
rect 37773 3066 37807 3100
rect 37773 2994 37807 3028
rect 37773 2922 37807 2956
rect 37773 2850 37807 2884
rect 37773 2778 37807 2812
rect 37773 2706 37807 2740
rect 37773 2634 37807 2668
rect 37773 2562 37807 2596
rect 37773 2490 37807 2524
rect 37773 2418 37807 2452
rect 37773 2346 37807 2380
rect 37773 2274 37807 2308
rect 37773 2202 37807 2236
rect 37773 2130 37807 2164
rect 37773 2058 37807 2092
rect 37773 1986 37807 2020
rect 37773 1914 37807 1948
rect 37773 1842 37807 1876
rect 37773 1770 37807 1804
rect 37773 1698 37807 1732
rect 37773 1626 37807 1660
rect 37773 1554 37807 1588
rect 37773 1482 37807 1516
rect 37773 1410 37807 1444
rect 37773 1338 37807 1372
rect 37773 1266 37807 1300
rect 37773 1194 37807 1228
rect 37869 3066 37903 3100
rect 37869 2994 37903 3028
rect 37869 2922 37903 2956
rect 37869 2850 37903 2884
rect 37869 2778 37903 2812
rect 37869 2706 37903 2740
rect 37869 2634 37903 2668
rect 37869 2562 37903 2596
rect 37869 2490 37903 2524
rect 37869 2418 37903 2452
rect 37869 2346 37903 2380
rect 37869 2274 37903 2308
rect 37869 2202 37903 2236
rect 37869 2130 37903 2164
rect 37869 2058 37903 2092
rect 37869 1986 37903 2020
rect 37869 1914 37903 1948
rect 37869 1842 37903 1876
rect 37869 1770 37903 1804
rect 37869 1698 37903 1732
rect 37869 1626 37903 1660
rect 37869 1554 37903 1588
rect 37869 1482 37903 1516
rect 37869 1410 37903 1444
rect 37869 1338 37903 1372
rect 37869 1266 37903 1300
rect 37869 1194 37903 1228
rect 37965 3066 37999 3100
rect 37965 2994 37999 3028
rect 37965 2922 37999 2956
rect 37965 2850 37999 2884
rect 37965 2778 37999 2812
rect 37965 2706 37999 2740
rect 37965 2634 37999 2668
rect 37965 2562 37999 2596
rect 37965 2490 37999 2524
rect 37965 2418 37999 2452
rect 37965 2346 37999 2380
rect 37965 2274 37999 2308
rect 37965 2202 37999 2236
rect 37965 2130 37999 2164
rect 37965 2058 37999 2092
rect 37965 1986 37999 2020
rect 37965 1914 37999 1948
rect 37965 1842 37999 1876
rect 37965 1770 37999 1804
rect 37965 1698 37999 1732
rect 37965 1626 37999 1660
rect 37965 1554 37999 1588
rect 37965 1482 37999 1516
rect 37965 1410 37999 1444
rect 37965 1338 37999 1372
rect 37965 1266 37999 1300
rect 37965 1194 37999 1228
rect 38061 3066 38095 3100
rect 38061 2994 38095 3028
rect 38061 2922 38095 2956
rect 38061 2850 38095 2884
rect 38061 2778 38095 2812
rect 38061 2706 38095 2740
rect 38061 2634 38095 2668
rect 38061 2562 38095 2596
rect 38061 2490 38095 2524
rect 38061 2418 38095 2452
rect 38061 2346 38095 2380
rect 38061 2274 38095 2308
rect 38061 2202 38095 2236
rect 38061 2130 38095 2164
rect 38061 2058 38095 2092
rect 38061 1986 38095 2020
rect 38061 1914 38095 1948
rect 38061 1842 38095 1876
rect 38061 1770 38095 1804
rect 38061 1698 38095 1732
rect 38061 1626 38095 1660
rect 38061 1554 38095 1588
rect 38061 1482 38095 1516
rect 38061 1410 38095 1444
rect 38061 1338 38095 1372
rect 38061 1266 38095 1300
rect 38061 1194 38095 1228
rect 38157 3066 38191 3100
rect 38157 2994 38191 3028
rect 38157 2922 38191 2956
rect 38157 2850 38191 2884
rect 38157 2778 38191 2812
rect 38157 2706 38191 2740
rect 38157 2634 38191 2668
rect 38157 2562 38191 2596
rect 38157 2490 38191 2524
rect 38157 2418 38191 2452
rect 38157 2346 38191 2380
rect 38157 2274 38191 2308
rect 38157 2202 38191 2236
rect 38157 2130 38191 2164
rect 38157 2058 38191 2092
rect 38157 1986 38191 2020
rect 38157 1914 38191 1948
rect 38157 1842 38191 1876
rect 38157 1770 38191 1804
rect 38157 1698 38191 1732
rect 38157 1626 38191 1660
rect 38157 1554 38191 1588
rect 38157 1482 38191 1516
rect 38157 1410 38191 1444
rect 38157 1338 38191 1372
rect 38157 1266 38191 1300
rect 38157 1194 38191 1228
rect 38253 3066 38287 3100
rect 38253 2994 38287 3028
rect 38253 2922 38287 2956
rect 38253 2850 38287 2884
rect 38253 2778 38287 2812
rect 38253 2706 38287 2740
rect 38253 2634 38287 2668
rect 38253 2562 38287 2596
rect 38253 2490 38287 2524
rect 38253 2418 38287 2452
rect 38253 2346 38287 2380
rect 38253 2274 38287 2308
rect 38253 2202 38287 2236
rect 38253 2130 38287 2164
rect 38253 2058 38287 2092
rect 38253 1986 38287 2020
rect 38253 1914 38287 1948
rect 38253 1842 38287 1876
rect 38253 1770 38287 1804
rect 38253 1698 38287 1732
rect 38253 1626 38287 1660
rect 38253 1554 38287 1588
rect 38253 1482 38287 1516
rect 38253 1410 38287 1444
rect 38253 1338 38287 1372
rect 38253 1266 38287 1300
rect 38253 1194 38287 1228
rect 38349 3066 38383 3100
rect 38349 2994 38383 3028
rect 38349 2922 38383 2956
rect 38349 2850 38383 2884
rect 38349 2778 38383 2812
rect 38349 2706 38383 2740
rect 38349 2634 38383 2668
rect 38349 2562 38383 2596
rect 38349 2490 38383 2524
rect 38349 2418 38383 2452
rect 38349 2346 38383 2380
rect 38349 2274 38383 2308
rect 38349 2202 38383 2236
rect 38349 2130 38383 2164
rect 38349 2058 38383 2092
rect 38349 1986 38383 2020
rect 38349 1914 38383 1948
rect 38349 1842 38383 1876
rect 38349 1770 38383 1804
rect 38349 1698 38383 1732
rect 38349 1626 38383 1660
rect 38349 1554 38383 1588
rect 38349 1482 38383 1516
rect 38349 1410 38383 1444
rect 38349 1338 38383 1372
rect 38349 1266 38383 1300
rect 38349 1194 38383 1228
rect 38445 3066 38479 3100
rect 38445 2994 38479 3028
rect 38445 2922 38479 2956
rect 38445 2850 38479 2884
rect 38445 2778 38479 2812
rect 38445 2706 38479 2740
rect 38445 2634 38479 2668
rect 38445 2562 38479 2596
rect 38445 2490 38479 2524
rect 38445 2418 38479 2452
rect 38445 2346 38479 2380
rect 38445 2274 38479 2308
rect 38445 2202 38479 2236
rect 38445 2130 38479 2164
rect 38445 2058 38479 2092
rect 38445 1986 38479 2020
rect 38445 1914 38479 1948
rect 38445 1842 38479 1876
rect 38445 1770 38479 1804
rect 38445 1698 38479 1732
rect 38445 1626 38479 1660
rect 38445 1554 38479 1588
rect 38445 1482 38479 1516
rect 38445 1410 38479 1444
rect 38445 1338 38479 1372
rect 38445 1266 38479 1300
rect 38445 1194 38479 1228
rect 38541 3066 38575 3100
rect 38541 2994 38575 3028
rect 38541 2922 38575 2956
rect 38541 2850 38575 2884
rect 38541 2778 38575 2812
rect 38541 2706 38575 2740
rect 38541 2634 38575 2668
rect 38541 2562 38575 2596
rect 38541 2490 38575 2524
rect 38541 2418 38575 2452
rect 38541 2346 38575 2380
rect 38541 2274 38575 2308
rect 38541 2202 38575 2236
rect 38541 2130 38575 2164
rect 38541 2058 38575 2092
rect 38541 1986 38575 2020
rect 38541 1914 38575 1948
rect 38541 1842 38575 1876
rect 38541 1770 38575 1804
rect 38541 1698 38575 1732
rect 38541 1626 38575 1660
rect 38541 1554 38575 1588
rect 38541 1482 38575 1516
rect 38541 1410 38575 1444
rect 38541 1338 38575 1372
rect 38541 1266 38575 1300
rect 38541 1194 38575 1228
rect 38637 3065 38671 3099
rect 38637 2993 38671 3027
rect 38637 2921 38671 2955
rect 38637 2849 38671 2883
rect 38637 2777 38671 2811
rect 38637 2705 38671 2739
rect 38637 2633 38671 2667
rect 38637 2561 38671 2595
rect 38637 2489 38671 2523
rect 38637 2417 38671 2451
rect 38637 2345 38671 2379
rect 38637 2273 38671 2307
rect 38637 2201 38671 2235
rect 38637 2129 38671 2163
rect 38637 2057 38671 2091
rect 38637 1985 38671 2019
rect 38637 1913 38671 1947
rect 38637 1841 38671 1875
rect 38637 1769 38671 1803
rect 38637 1697 38671 1731
rect 38637 1625 38671 1659
rect 38637 1553 38671 1587
rect 38637 1481 38671 1515
rect 38637 1409 38671 1443
rect 38637 1337 38671 1371
rect 38637 1265 38671 1299
rect 38637 1193 38671 1227
rect 29100 1065 29134 1099
rect 29172 1065 29206 1099
rect 29244 1065 29278 1099
rect 29316 1065 29350 1099
rect 29388 1065 29422 1099
rect 29460 1065 29494 1099
rect 29532 1065 29566 1099
rect 29604 1065 29638 1099
rect 29676 1065 29710 1099
rect 29748 1065 29782 1099
rect 29820 1065 29854 1099
rect 29892 1065 29926 1099
rect 29964 1065 29998 1099
rect 30036 1065 30070 1099
rect 30108 1065 30142 1099
rect 30180 1065 30214 1099
rect 30252 1065 30286 1099
rect 30324 1065 30358 1099
rect 30396 1065 30430 1099
rect 30468 1065 30502 1099
rect 30540 1065 30574 1099
rect 30612 1065 30646 1099
rect 30684 1065 30718 1099
rect 30756 1065 30790 1099
rect 30828 1065 30862 1099
rect 30900 1065 30934 1099
rect 30972 1065 31006 1099
rect 31044 1065 31078 1099
rect 31116 1065 31150 1099
rect 31188 1065 31222 1099
rect 31260 1065 31294 1099
rect 31332 1065 31366 1099
rect 31404 1065 31438 1099
rect 31476 1065 31510 1099
rect 31548 1065 31582 1099
rect 31620 1065 31654 1099
rect 31692 1065 31726 1099
rect 31764 1065 31798 1099
rect 31836 1065 31870 1099
rect 31908 1065 31942 1099
rect 31980 1065 32014 1099
rect 32052 1065 32086 1099
rect 32124 1065 32158 1099
rect 32196 1065 32230 1099
rect 32268 1065 32302 1099
rect 32340 1065 32374 1099
rect 32412 1065 32446 1099
rect 32484 1065 32518 1099
rect 32556 1065 32590 1099
rect 32628 1065 32662 1099
rect 32700 1065 32734 1099
rect 32772 1065 32806 1099
rect 32844 1065 32878 1099
rect 32916 1065 32950 1099
rect 32988 1065 33022 1099
rect 33060 1065 33094 1099
rect 33132 1065 33166 1099
rect 33204 1065 33238 1099
rect 33276 1065 33310 1099
rect 33348 1065 33382 1099
rect 33420 1065 33454 1099
rect 33492 1065 33526 1099
rect 33564 1065 33598 1099
rect 33636 1065 33670 1099
rect 33708 1065 33742 1099
rect 33780 1065 33814 1099
rect 33852 1065 33886 1099
rect 33924 1065 33958 1099
rect 33996 1065 34030 1099
rect 34068 1065 34102 1099
rect 34140 1065 34174 1099
rect 34212 1065 34246 1099
rect 34284 1065 34318 1099
rect 34356 1065 34390 1099
rect 34428 1065 34462 1099
rect 34500 1065 34534 1099
rect 34572 1065 34606 1099
rect 34644 1065 34678 1099
rect 34716 1065 34750 1099
rect 34788 1065 34822 1099
rect 34860 1065 34894 1099
rect 34932 1065 34966 1099
rect 35004 1065 35038 1099
rect 35076 1065 35110 1099
rect 35148 1065 35182 1099
rect 35220 1065 35254 1099
rect 35292 1065 35326 1099
rect 35364 1065 35398 1099
rect 35436 1065 35470 1099
rect 35508 1065 35542 1099
rect 35580 1065 35614 1099
rect 35652 1065 35686 1099
rect 35724 1065 35758 1099
rect 35796 1065 35830 1099
rect 35868 1065 35902 1099
rect 35940 1065 35974 1099
rect 36012 1065 36046 1099
rect 36084 1065 36118 1099
rect 36156 1065 36190 1099
rect 36228 1065 36262 1099
rect 36300 1065 36334 1099
rect 36372 1065 36406 1099
rect 36444 1065 36478 1099
rect 36516 1065 36550 1099
rect 36588 1065 36622 1099
rect 36660 1065 36694 1099
rect 36732 1065 36766 1099
rect 36804 1065 36838 1099
rect 36876 1065 36910 1099
rect 36948 1065 36982 1099
rect 37020 1065 37054 1099
rect 37092 1065 37126 1099
rect 37164 1065 37198 1099
rect 37236 1065 37270 1099
rect 37308 1065 37342 1099
rect 37380 1065 37414 1099
rect 37452 1065 37486 1099
rect 37524 1065 37558 1099
rect 37596 1065 37630 1099
rect 37668 1065 37702 1099
rect 37740 1065 37774 1099
rect 37812 1065 37846 1099
rect 37884 1065 37918 1099
rect 37956 1065 37990 1099
rect 38028 1065 38062 1099
rect 38100 1065 38134 1099
rect 38172 1065 38206 1099
rect 38244 1065 38278 1099
rect 38316 1065 38350 1099
rect 38388 1065 38422 1099
rect 38460 1065 38494 1099
<< metal1 >>
rect 29140 3223 38986 3250
rect 29140 3189 29200 3223
rect 29234 3189 29272 3223
rect 29306 3189 29344 3223
rect 29378 3189 29416 3223
rect 29450 3189 29488 3223
rect 29522 3189 29560 3223
rect 29594 3189 29632 3223
rect 29666 3189 29704 3223
rect 29738 3189 29776 3223
rect 29810 3189 29848 3223
rect 29882 3189 29920 3223
rect 29954 3189 29992 3223
rect 30026 3189 30064 3223
rect 30098 3189 30136 3223
rect 30170 3189 30208 3223
rect 30242 3189 30280 3223
rect 30314 3189 30352 3223
rect 30386 3189 30424 3223
rect 30458 3189 30496 3223
rect 30530 3189 30568 3223
rect 30602 3189 30640 3223
rect 30674 3189 30712 3223
rect 30746 3189 30784 3223
rect 30818 3189 30856 3223
rect 30890 3189 30928 3223
rect 30962 3189 31000 3223
rect 31034 3189 31072 3223
rect 31106 3189 31144 3223
rect 31178 3189 31216 3223
rect 31250 3189 31288 3223
rect 31322 3189 31360 3223
rect 31394 3189 31432 3223
rect 31466 3189 31504 3223
rect 31538 3189 31576 3223
rect 31610 3189 31648 3223
rect 31682 3189 31720 3223
rect 31754 3189 31792 3223
rect 31826 3189 31864 3223
rect 31898 3189 31936 3223
rect 31970 3189 32008 3223
rect 32042 3189 32080 3223
rect 32114 3189 32152 3223
rect 32186 3189 32224 3223
rect 32258 3189 32296 3223
rect 32330 3189 32368 3223
rect 32402 3189 32440 3223
rect 32474 3189 32512 3223
rect 32546 3189 32584 3223
rect 32618 3189 32656 3223
rect 32690 3189 32728 3223
rect 32762 3189 32800 3223
rect 32834 3189 32872 3223
rect 32906 3189 32944 3223
rect 32978 3189 33016 3223
rect 33050 3189 33088 3223
rect 33122 3189 33160 3223
rect 33194 3189 33232 3223
rect 33266 3189 33304 3223
rect 33338 3189 33376 3223
rect 33410 3189 33448 3223
rect 33482 3189 33520 3223
rect 33554 3189 33592 3223
rect 33626 3189 33664 3223
rect 33698 3189 33736 3223
rect 33770 3189 33808 3223
rect 33842 3189 33880 3223
rect 33914 3189 33952 3223
rect 33986 3189 34024 3223
rect 34058 3189 34096 3223
rect 34130 3189 34168 3223
rect 34202 3189 34240 3223
rect 34274 3189 34312 3223
rect 34346 3189 34384 3223
rect 34418 3189 34456 3223
rect 34490 3189 34528 3223
rect 34562 3189 34600 3223
rect 34634 3189 34672 3223
rect 34706 3189 34744 3223
rect 34778 3189 34816 3223
rect 34850 3189 34888 3223
rect 34922 3189 34960 3223
rect 34994 3189 35032 3223
rect 35066 3189 35104 3223
rect 35138 3189 35176 3223
rect 35210 3189 35248 3223
rect 35282 3189 35320 3223
rect 35354 3189 35392 3223
rect 35426 3189 35464 3223
rect 35498 3189 35536 3223
rect 35570 3189 35608 3223
rect 35642 3189 35680 3223
rect 35714 3189 35752 3223
rect 35786 3189 35824 3223
rect 35858 3189 35896 3223
rect 35930 3189 35968 3223
rect 36002 3189 36040 3223
rect 36074 3189 36112 3223
rect 36146 3189 36184 3223
rect 36218 3189 36256 3223
rect 36290 3189 36328 3223
rect 36362 3189 36400 3223
rect 36434 3189 36472 3223
rect 36506 3189 36544 3223
rect 36578 3189 36616 3223
rect 36650 3189 36688 3223
rect 36722 3189 36760 3223
rect 36794 3189 36832 3223
rect 36866 3189 36904 3223
rect 36938 3189 36976 3223
rect 37010 3189 37048 3223
rect 37082 3189 37120 3223
rect 37154 3189 37192 3223
rect 37226 3189 37264 3223
rect 37298 3189 37336 3223
rect 37370 3189 37408 3223
rect 37442 3189 37480 3223
rect 37514 3189 37552 3223
rect 37586 3189 37624 3223
rect 37658 3189 37696 3223
rect 37730 3189 37768 3223
rect 37802 3189 37840 3223
rect 37874 3189 37912 3223
rect 37946 3189 37984 3223
rect 38018 3189 38056 3223
rect 38090 3189 38128 3223
rect 38162 3189 38200 3223
rect 38234 3189 38272 3223
rect 38306 3189 38344 3223
rect 38378 3189 38416 3223
rect 38450 3189 38488 3223
rect 38522 3189 38560 3223
rect 38594 3189 38986 3223
rect 29140 3180 38986 3189
rect 29140 3176 29186 3180
rect 29025 3133 29083 3147
rect 29025 3081 29028 3133
rect 29080 3081 29083 3133
rect 29025 3069 29037 3081
rect 29071 3069 29083 3081
rect 29025 3017 29028 3069
rect 29080 3017 29083 3069
rect 29025 3005 29037 3017
rect 29071 3005 29083 3017
rect 29025 2953 29028 3005
rect 29080 2953 29083 3005
rect 29025 2941 29037 2953
rect 29071 2941 29083 2953
rect 29025 2889 29028 2941
rect 29080 2889 29083 2941
rect 29025 2884 29083 2889
rect 29025 2877 29037 2884
rect 29071 2877 29083 2884
rect 29025 2825 29028 2877
rect 29080 2825 29083 2877
rect 29025 2813 29083 2825
rect 29025 2761 29028 2813
rect 29080 2761 29083 2813
rect 29025 2749 29083 2761
rect 29025 2697 29028 2749
rect 29080 2697 29083 2749
rect 29025 2685 29083 2697
rect 29025 2633 29028 2685
rect 29080 2633 29083 2685
rect 29025 2621 29083 2633
rect 29025 2569 29028 2621
rect 29080 2569 29083 2621
rect 29025 2562 29037 2569
rect 29071 2562 29083 2569
rect 29025 2557 29083 2562
rect 29025 2505 29028 2557
rect 29080 2505 29083 2557
rect 29025 2493 29037 2505
rect 29071 2493 29083 2505
rect 29025 2441 29028 2493
rect 29080 2441 29083 2493
rect 29025 2429 29037 2441
rect 29071 2429 29083 2441
rect 29025 2377 29028 2429
rect 29080 2377 29083 2429
rect 29025 2365 29037 2377
rect 29071 2365 29083 2377
rect 29025 2313 29028 2365
rect 29080 2313 29083 2365
rect 29025 2308 29083 2313
rect 29025 2301 29037 2308
rect 29071 2301 29083 2308
rect 29025 2249 29028 2301
rect 29080 2249 29083 2301
rect 29025 2237 29083 2249
rect 29025 2185 29028 2237
rect 29080 2185 29083 2237
rect 29025 2173 29083 2185
rect 29025 2121 29028 2173
rect 29080 2121 29083 2173
rect 29025 2109 29083 2121
rect 29025 2057 29028 2109
rect 29080 2057 29083 2109
rect 29025 2045 29083 2057
rect 29025 1993 29028 2045
rect 29080 1993 29083 2045
rect 29025 1986 29037 1993
rect 29071 1986 29083 1993
rect 29025 1981 29083 1986
rect 29025 1929 29028 1981
rect 29080 1929 29083 1981
rect 29025 1917 29037 1929
rect 29071 1917 29083 1929
rect 29025 1865 29028 1917
rect 29080 1865 29083 1917
rect 29025 1853 29037 1865
rect 29071 1853 29083 1865
rect 29025 1801 29028 1853
rect 29080 1801 29083 1853
rect 29025 1789 29037 1801
rect 29071 1789 29083 1801
rect 29025 1737 29028 1789
rect 29080 1737 29083 1789
rect 29025 1732 29083 1737
rect 29025 1725 29037 1732
rect 29071 1725 29083 1732
rect 29025 1673 29028 1725
rect 29080 1673 29083 1725
rect 29025 1661 29083 1673
rect 29025 1609 29028 1661
rect 29080 1609 29083 1661
rect 29025 1597 29083 1609
rect 29025 1545 29028 1597
rect 29080 1545 29083 1597
rect 29025 1533 29083 1545
rect 29025 1481 29028 1533
rect 29080 1481 29083 1533
rect 29025 1469 29083 1481
rect 29025 1417 29028 1469
rect 29080 1417 29083 1469
rect 29025 1410 29037 1417
rect 29071 1410 29083 1417
rect 29025 1405 29083 1410
rect 29025 1353 29028 1405
rect 29080 1353 29083 1405
rect 29025 1341 29037 1353
rect 29071 1341 29083 1353
rect 29025 1289 29028 1341
rect 29080 1289 29083 1341
rect 29025 1277 29037 1289
rect 29071 1277 29083 1289
rect 29025 1225 29028 1277
rect 29080 1225 29083 1277
rect 29025 1213 29037 1225
rect 29071 1213 29083 1225
rect 29025 1161 29028 1213
rect 29080 1161 29083 1213
rect 29025 1147 29083 1161
rect 29121 3133 29179 3147
rect 29121 3081 29124 3133
rect 29176 3081 29179 3133
rect 29121 3069 29133 3081
rect 29167 3069 29179 3081
rect 29121 3017 29124 3069
rect 29176 3017 29179 3069
rect 29121 3005 29133 3017
rect 29167 3005 29179 3017
rect 29121 2953 29124 3005
rect 29176 2953 29179 3005
rect 29121 2941 29133 2953
rect 29167 2941 29179 2953
rect 29121 2889 29124 2941
rect 29176 2889 29179 2941
rect 29121 2884 29179 2889
rect 29121 2877 29133 2884
rect 29167 2877 29179 2884
rect 29121 2825 29124 2877
rect 29176 2825 29179 2877
rect 29121 2813 29179 2825
rect 29121 2761 29124 2813
rect 29176 2761 29179 2813
rect 29121 2749 29179 2761
rect 29121 2697 29124 2749
rect 29176 2697 29179 2749
rect 29121 2685 29179 2697
rect 29121 2633 29124 2685
rect 29176 2633 29179 2685
rect 29121 2621 29179 2633
rect 29121 2569 29124 2621
rect 29176 2569 29179 2621
rect 29121 2562 29133 2569
rect 29167 2562 29179 2569
rect 29121 2557 29179 2562
rect 29121 2505 29124 2557
rect 29176 2505 29179 2557
rect 29121 2493 29133 2505
rect 29167 2493 29179 2505
rect 29121 2441 29124 2493
rect 29176 2441 29179 2493
rect 29121 2429 29133 2441
rect 29167 2429 29179 2441
rect 29121 2377 29124 2429
rect 29176 2377 29179 2429
rect 29121 2365 29133 2377
rect 29167 2365 29179 2377
rect 29121 2313 29124 2365
rect 29176 2313 29179 2365
rect 29121 2308 29179 2313
rect 29121 2301 29133 2308
rect 29167 2301 29179 2308
rect 29121 2249 29124 2301
rect 29176 2249 29179 2301
rect 29121 2237 29179 2249
rect 29121 2185 29124 2237
rect 29176 2185 29179 2237
rect 29121 2173 29179 2185
rect 29121 2121 29124 2173
rect 29176 2121 29179 2173
rect 29121 2109 29179 2121
rect 29121 2057 29124 2109
rect 29176 2057 29179 2109
rect 29121 2045 29179 2057
rect 29121 1993 29124 2045
rect 29176 1993 29179 2045
rect 29121 1986 29133 1993
rect 29167 1986 29179 1993
rect 29121 1981 29179 1986
rect 29121 1929 29124 1981
rect 29176 1929 29179 1981
rect 29121 1917 29133 1929
rect 29167 1917 29179 1929
rect 29121 1865 29124 1917
rect 29176 1865 29179 1917
rect 29121 1853 29133 1865
rect 29167 1853 29179 1865
rect 29121 1801 29124 1853
rect 29176 1801 29179 1853
rect 29121 1789 29133 1801
rect 29167 1789 29179 1801
rect 29121 1737 29124 1789
rect 29176 1737 29179 1789
rect 29121 1732 29179 1737
rect 29121 1725 29133 1732
rect 29167 1725 29179 1732
rect 29121 1673 29124 1725
rect 29176 1673 29179 1725
rect 29121 1661 29179 1673
rect 29121 1609 29124 1661
rect 29176 1609 29179 1661
rect 29121 1597 29179 1609
rect 29121 1545 29124 1597
rect 29176 1545 29179 1597
rect 29121 1533 29179 1545
rect 29121 1481 29124 1533
rect 29176 1481 29179 1533
rect 29121 1469 29179 1481
rect 29121 1417 29124 1469
rect 29176 1417 29179 1469
rect 29121 1410 29133 1417
rect 29167 1410 29179 1417
rect 29121 1405 29179 1410
rect 29121 1353 29124 1405
rect 29176 1353 29179 1405
rect 29121 1341 29133 1353
rect 29167 1341 29179 1353
rect 29121 1289 29124 1341
rect 29176 1289 29179 1341
rect 29121 1277 29133 1289
rect 29167 1277 29179 1289
rect 29121 1225 29124 1277
rect 29176 1225 29179 1277
rect 29121 1213 29133 1225
rect 29167 1213 29179 1225
rect 29121 1161 29124 1213
rect 29176 1161 29179 1213
rect 29121 1147 29179 1161
rect 29217 3133 29275 3147
rect 29217 3081 29220 3133
rect 29272 3081 29275 3133
rect 29217 3069 29229 3081
rect 29263 3069 29275 3081
rect 29217 3017 29220 3069
rect 29272 3017 29275 3069
rect 29217 3005 29229 3017
rect 29263 3005 29275 3017
rect 29217 2953 29220 3005
rect 29272 2953 29275 3005
rect 29217 2941 29229 2953
rect 29263 2941 29275 2953
rect 29217 2889 29220 2941
rect 29272 2889 29275 2941
rect 29217 2884 29275 2889
rect 29217 2877 29229 2884
rect 29263 2877 29275 2884
rect 29217 2825 29220 2877
rect 29272 2825 29275 2877
rect 29217 2813 29275 2825
rect 29217 2761 29220 2813
rect 29272 2761 29275 2813
rect 29217 2749 29275 2761
rect 29217 2697 29220 2749
rect 29272 2697 29275 2749
rect 29217 2685 29275 2697
rect 29217 2633 29220 2685
rect 29272 2633 29275 2685
rect 29217 2621 29275 2633
rect 29217 2569 29220 2621
rect 29272 2569 29275 2621
rect 29217 2562 29229 2569
rect 29263 2562 29275 2569
rect 29217 2557 29275 2562
rect 29217 2505 29220 2557
rect 29272 2505 29275 2557
rect 29217 2493 29229 2505
rect 29263 2493 29275 2505
rect 29217 2441 29220 2493
rect 29272 2441 29275 2493
rect 29217 2429 29229 2441
rect 29263 2429 29275 2441
rect 29217 2377 29220 2429
rect 29272 2377 29275 2429
rect 29217 2365 29229 2377
rect 29263 2365 29275 2377
rect 29217 2313 29220 2365
rect 29272 2313 29275 2365
rect 29217 2308 29275 2313
rect 29217 2301 29229 2308
rect 29263 2301 29275 2308
rect 29217 2249 29220 2301
rect 29272 2249 29275 2301
rect 29217 2237 29275 2249
rect 29217 2185 29220 2237
rect 29272 2185 29275 2237
rect 29217 2173 29275 2185
rect 29217 2121 29220 2173
rect 29272 2121 29275 2173
rect 29217 2109 29275 2121
rect 29217 2057 29220 2109
rect 29272 2057 29275 2109
rect 29217 2045 29275 2057
rect 29217 1993 29220 2045
rect 29272 1993 29275 2045
rect 29217 1986 29229 1993
rect 29263 1986 29275 1993
rect 29217 1981 29275 1986
rect 29217 1929 29220 1981
rect 29272 1929 29275 1981
rect 29217 1917 29229 1929
rect 29263 1917 29275 1929
rect 29217 1865 29220 1917
rect 29272 1865 29275 1917
rect 29217 1853 29229 1865
rect 29263 1853 29275 1865
rect 29217 1801 29220 1853
rect 29272 1801 29275 1853
rect 29217 1789 29229 1801
rect 29263 1789 29275 1801
rect 29217 1737 29220 1789
rect 29272 1737 29275 1789
rect 29217 1732 29275 1737
rect 29217 1725 29229 1732
rect 29263 1725 29275 1732
rect 29217 1673 29220 1725
rect 29272 1673 29275 1725
rect 29217 1661 29275 1673
rect 29217 1609 29220 1661
rect 29272 1609 29275 1661
rect 29217 1597 29275 1609
rect 29217 1545 29220 1597
rect 29272 1545 29275 1597
rect 29217 1533 29275 1545
rect 29217 1481 29220 1533
rect 29272 1481 29275 1533
rect 29217 1469 29275 1481
rect 29217 1417 29220 1469
rect 29272 1417 29275 1469
rect 29217 1410 29229 1417
rect 29263 1410 29275 1417
rect 29217 1405 29275 1410
rect 29217 1353 29220 1405
rect 29272 1353 29275 1405
rect 29217 1341 29229 1353
rect 29263 1341 29275 1353
rect 29217 1289 29220 1341
rect 29272 1289 29275 1341
rect 29217 1277 29229 1289
rect 29263 1277 29275 1289
rect 29217 1225 29220 1277
rect 29272 1225 29275 1277
rect 29217 1213 29229 1225
rect 29263 1213 29275 1225
rect 29217 1161 29220 1213
rect 29272 1161 29275 1213
rect 29217 1147 29275 1161
rect 29316 3133 29368 3147
rect 29316 3069 29325 3081
rect 29359 3069 29368 3081
rect 29316 3005 29325 3017
rect 29359 3005 29368 3017
rect 29316 2941 29325 2953
rect 29359 2941 29368 2953
rect 29316 2884 29368 2889
rect 29316 2877 29325 2884
rect 29359 2877 29368 2884
rect 29316 2813 29368 2825
rect 29316 2749 29368 2761
rect 29316 2685 29368 2697
rect 29316 2621 29368 2633
rect 29316 2562 29325 2569
rect 29359 2562 29368 2569
rect 29316 2557 29368 2562
rect 29316 2493 29325 2505
rect 29359 2493 29368 2505
rect 29316 2429 29325 2441
rect 29359 2429 29368 2441
rect 29316 2365 29325 2377
rect 29359 2365 29368 2377
rect 29316 2308 29368 2313
rect 29316 2301 29325 2308
rect 29359 2301 29368 2308
rect 29316 2237 29368 2249
rect 29316 2173 29368 2185
rect 29316 2109 29368 2121
rect 29316 2045 29368 2057
rect 29316 1986 29325 1993
rect 29359 1986 29368 1993
rect 29316 1981 29368 1986
rect 29316 1917 29325 1929
rect 29359 1917 29368 1929
rect 29316 1853 29325 1865
rect 29359 1853 29368 1865
rect 29316 1789 29325 1801
rect 29359 1789 29368 1801
rect 29316 1732 29368 1737
rect 29316 1725 29325 1732
rect 29359 1725 29368 1732
rect 29316 1661 29368 1673
rect 29316 1597 29368 1609
rect 29316 1533 29368 1545
rect 29316 1469 29368 1481
rect 29316 1410 29325 1417
rect 29359 1410 29368 1417
rect 29316 1405 29368 1410
rect 29316 1341 29325 1353
rect 29359 1341 29368 1353
rect 29316 1277 29325 1289
rect 29359 1277 29368 1289
rect 29316 1213 29325 1225
rect 29359 1213 29368 1225
rect 29316 1147 29368 1161
rect 29409 3133 29467 3147
rect 29409 3081 29412 3133
rect 29464 3081 29467 3133
rect 29409 3069 29421 3081
rect 29455 3069 29467 3081
rect 29409 3017 29412 3069
rect 29464 3017 29467 3069
rect 29409 3005 29421 3017
rect 29455 3005 29467 3017
rect 29409 2953 29412 3005
rect 29464 2953 29467 3005
rect 29409 2941 29421 2953
rect 29455 2941 29467 2953
rect 29409 2889 29412 2941
rect 29464 2889 29467 2941
rect 29409 2884 29467 2889
rect 29409 2877 29421 2884
rect 29455 2877 29467 2884
rect 29409 2825 29412 2877
rect 29464 2825 29467 2877
rect 29409 2813 29467 2825
rect 29409 2761 29412 2813
rect 29464 2761 29467 2813
rect 29409 2749 29467 2761
rect 29409 2697 29412 2749
rect 29464 2697 29467 2749
rect 29409 2685 29467 2697
rect 29409 2633 29412 2685
rect 29464 2633 29467 2685
rect 29409 2621 29467 2633
rect 29409 2569 29412 2621
rect 29464 2569 29467 2621
rect 29409 2562 29421 2569
rect 29455 2562 29467 2569
rect 29409 2557 29467 2562
rect 29409 2505 29412 2557
rect 29464 2505 29467 2557
rect 29409 2493 29421 2505
rect 29455 2493 29467 2505
rect 29409 2441 29412 2493
rect 29464 2441 29467 2493
rect 29409 2429 29421 2441
rect 29455 2429 29467 2441
rect 29409 2377 29412 2429
rect 29464 2377 29467 2429
rect 29409 2365 29421 2377
rect 29455 2365 29467 2377
rect 29409 2313 29412 2365
rect 29464 2313 29467 2365
rect 29409 2308 29467 2313
rect 29409 2301 29421 2308
rect 29455 2301 29467 2308
rect 29409 2249 29412 2301
rect 29464 2249 29467 2301
rect 29409 2237 29467 2249
rect 29409 2185 29412 2237
rect 29464 2185 29467 2237
rect 29409 2173 29467 2185
rect 29409 2121 29412 2173
rect 29464 2121 29467 2173
rect 29409 2109 29467 2121
rect 29409 2057 29412 2109
rect 29464 2057 29467 2109
rect 29409 2045 29467 2057
rect 29409 1993 29412 2045
rect 29464 1993 29467 2045
rect 29409 1986 29421 1993
rect 29455 1986 29467 1993
rect 29409 1981 29467 1986
rect 29409 1929 29412 1981
rect 29464 1929 29467 1981
rect 29409 1917 29421 1929
rect 29455 1917 29467 1929
rect 29409 1865 29412 1917
rect 29464 1865 29467 1917
rect 29409 1853 29421 1865
rect 29455 1853 29467 1865
rect 29409 1801 29412 1853
rect 29464 1801 29467 1853
rect 29409 1789 29421 1801
rect 29455 1789 29467 1801
rect 29409 1737 29412 1789
rect 29464 1737 29467 1789
rect 29409 1732 29467 1737
rect 29409 1725 29421 1732
rect 29455 1725 29467 1732
rect 29409 1673 29412 1725
rect 29464 1673 29467 1725
rect 29409 1661 29467 1673
rect 29409 1609 29412 1661
rect 29464 1609 29467 1661
rect 29409 1597 29467 1609
rect 29409 1545 29412 1597
rect 29464 1545 29467 1597
rect 29409 1533 29467 1545
rect 29409 1481 29412 1533
rect 29464 1481 29467 1533
rect 29409 1469 29467 1481
rect 29409 1417 29412 1469
rect 29464 1417 29467 1469
rect 29409 1410 29421 1417
rect 29455 1410 29467 1417
rect 29409 1405 29467 1410
rect 29409 1353 29412 1405
rect 29464 1353 29467 1405
rect 29409 1341 29421 1353
rect 29455 1341 29467 1353
rect 29409 1289 29412 1341
rect 29464 1289 29467 1341
rect 29409 1277 29421 1289
rect 29455 1277 29467 1289
rect 29409 1225 29412 1277
rect 29464 1225 29467 1277
rect 29409 1213 29421 1225
rect 29455 1213 29467 1225
rect 29409 1161 29412 1213
rect 29464 1161 29467 1213
rect 29409 1147 29467 1161
rect 29505 3133 29563 3147
rect 29505 3081 29508 3133
rect 29560 3081 29563 3133
rect 29505 3069 29517 3081
rect 29551 3069 29563 3081
rect 29505 3017 29508 3069
rect 29560 3017 29563 3069
rect 29505 3005 29517 3017
rect 29551 3005 29563 3017
rect 29505 2953 29508 3005
rect 29560 2953 29563 3005
rect 29505 2941 29517 2953
rect 29551 2941 29563 2953
rect 29505 2889 29508 2941
rect 29560 2889 29563 2941
rect 29505 2884 29563 2889
rect 29505 2877 29517 2884
rect 29551 2877 29563 2884
rect 29505 2825 29508 2877
rect 29560 2825 29563 2877
rect 29505 2813 29563 2825
rect 29505 2761 29508 2813
rect 29560 2761 29563 2813
rect 29505 2749 29563 2761
rect 29505 2697 29508 2749
rect 29560 2697 29563 2749
rect 29505 2685 29563 2697
rect 29505 2633 29508 2685
rect 29560 2633 29563 2685
rect 29505 2621 29563 2633
rect 29505 2569 29508 2621
rect 29560 2569 29563 2621
rect 29505 2562 29517 2569
rect 29551 2562 29563 2569
rect 29505 2557 29563 2562
rect 29505 2505 29508 2557
rect 29560 2505 29563 2557
rect 29505 2493 29517 2505
rect 29551 2493 29563 2505
rect 29505 2441 29508 2493
rect 29560 2441 29563 2493
rect 29505 2429 29517 2441
rect 29551 2429 29563 2441
rect 29505 2377 29508 2429
rect 29560 2377 29563 2429
rect 29505 2365 29517 2377
rect 29551 2365 29563 2377
rect 29505 2313 29508 2365
rect 29560 2313 29563 2365
rect 29505 2308 29563 2313
rect 29505 2301 29517 2308
rect 29551 2301 29563 2308
rect 29505 2249 29508 2301
rect 29560 2249 29563 2301
rect 29505 2237 29563 2249
rect 29505 2185 29508 2237
rect 29560 2185 29563 2237
rect 29505 2173 29563 2185
rect 29505 2121 29508 2173
rect 29560 2121 29563 2173
rect 29505 2109 29563 2121
rect 29505 2057 29508 2109
rect 29560 2057 29563 2109
rect 29505 2045 29563 2057
rect 29505 1993 29508 2045
rect 29560 1993 29563 2045
rect 29505 1986 29517 1993
rect 29551 1986 29563 1993
rect 29505 1981 29563 1986
rect 29505 1929 29508 1981
rect 29560 1929 29563 1981
rect 29505 1917 29517 1929
rect 29551 1917 29563 1929
rect 29505 1865 29508 1917
rect 29560 1865 29563 1917
rect 29505 1853 29517 1865
rect 29551 1853 29563 1865
rect 29505 1801 29508 1853
rect 29560 1801 29563 1853
rect 29505 1789 29517 1801
rect 29551 1789 29563 1801
rect 29505 1737 29508 1789
rect 29560 1737 29563 1789
rect 29505 1732 29563 1737
rect 29505 1725 29517 1732
rect 29551 1725 29563 1732
rect 29505 1673 29508 1725
rect 29560 1673 29563 1725
rect 29505 1661 29563 1673
rect 29505 1609 29508 1661
rect 29560 1609 29563 1661
rect 29505 1597 29563 1609
rect 29505 1545 29508 1597
rect 29560 1545 29563 1597
rect 29505 1533 29563 1545
rect 29505 1481 29508 1533
rect 29560 1481 29563 1533
rect 29505 1469 29563 1481
rect 29505 1417 29508 1469
rect 29560 1417 29563 1469
rect 29505 1410 29517 1417
rect 29551 1410 29563 1417
rect 29505 1405 29563 1410
rect 29505 1353 29508 1405
rect 29560 1353 29563 1405
rect 29505 1341 29517 1353
rect 29551 1341 29563 1353
rect 29505 1289 29508 1341
rect 29560 1289 29563 1341
rect 29505 1277 29517 1289
rect 29551 1277 29563 1289
rect 29505 1225 29508 1277
rect 29560 1225 29563 1277
rect 29505 1213 29517 1225
rect 29551 1213 29563 1225
rect 29505 1161 29508 1213
rect 29560 1161 29563 1213
rect 29505 1147 29563 1161
rect 29601 3133 29659 3147
rect 29601 3081 29604 3133
rect 29656 3081 29659 3133
rect 29601 3069 29613 3081
rect 29647 3069 29659 3081
rect 29601 3017 29604 3069
rect 29656 3017 29659 3069
rect 29601 3005 29613 3017
rect 29647 3005 29659 3017
rect 29601 2953 29604 3005
rect 29656 2953 29659 3005
rect 29601 2941 29613 2953
rect 29647 2941 29659 2953
rect 29601 2889 29604 2941
rect 29656 2889 29659 2941
rect 29601 2884 29659 2889
rect 29601 2877 29613 2884
rect 29647 2877 29659 2884
rect 29601 2825 29604 2877
rect 29656 2825 29659 2877
rect 29601 2813 29659 2825
rect 29601 2761 29604 2813
rect 29656 2761 29659 2813
rect 29601 2749 29659 2761
rect 29601 2697 29604 2749
rect 29656 2697 29659 2749
rect 29601 2685 29659 2697
rect 29601 2633 29604 2685
rect 29656 2633 29659 2685
rect 29601 2621 29659 2633
rect 29601 2569 29604 2621
rect 29656 2569 29659 2621
rect 29601 2562 29613 2569
rect 29647 2562 29659 2569
rect 29601 2557 29659 2562
rect 29601 2505 29604 2557
rect 29656 2505 29659 2557
rect 29601 2493 29613 2505
rect 29647 2493 29659 2505
rect 29601 2441 29604 2493
rect 29656 2441 29659 2493
rect 29601 2429 29613 2441
rect 29647 2429 29659 2441
rect 29601 2377 29604 2429
rect 29656 2377 29659 2429
rect 29601 2365 29613 2377
rect 29647 2365 29659 2377
rect 29601 2313 29604 2365
rect 29656 2313 29659 2365
rect 29601 2308 29659 2313
rect 29601 2301 29613 2308
rect 29647 2301 29659 2308
rect 29601 2249 29604 2301
rect 29656 2249 29659 2301
rect 29601 2237 29659 2249
rect 29601 2185 29604 2237
rect 29656 2185 29659 2237
rect 29601 2173 29659 2185
rect 29601 2121 29604 2173
rect 29656 2121 29659 2173
rect 29601 2109 29659 2121
rect 29601 2057 29604 2109
rect 29656 2057 29659 2109
rect 29601 2045 29659 2057
rect 29601 1993 29604 2045
rect 29656 1993 29659 2045
rect 29601 1986 29613 1993
rect 29647 1986 29659 1993
rect 29601 1981 29659 1986
rect 29601 1929 29604 1981
rect 29656 1929 29659 1981
rect 29601 1917 29613 1929
rect 29647 1917 29659 1929
rect 29601 1865 29604 1917
rect 29656 1865 29659 1917
rect 29601 1853 29613 1865
rect 29647 1853 29659 1865
rect 29601 1801 29604 1853
rect 29656 1801 29659 1853
rect 29601 1789 29613 1801
rect 29647 1789 29659 1801
rect 29601 1737 29604 1789
rect 29656 1737 29659 1789
rect 29601 1732 29659 1737
rect 29601 1725 29613 1732
rect 29647 1725 29659 1732
rect 29601 1673 29604 1725
rect 29656 1673 29659 1725
rect 29601 1661 29659 1673
rect 29601 1609 29604 1661
rect 29656 1609 29659 1661
rect 29601 1597 29659 1609
rect 29601 1545 29604 1597
rect 29656 1545 29659 1597
rect 29601 1533 29659 1545
rect 29601 1481 29604 1533
rect 29656 1481 29659 1533
rect 29601 1469 29659 1481
rect 29601 1417 29604 1469
rect 29656 1417 29659 1469
rect 29601 1410 29613 1417
rect 29647 1410 29659 1417
rect 29601 1405 29659 1410
rect 29601 1353 29604 1405
rect 29656 1353 29659 1405
rect 29601 1341 29613 1353
rect 29647 1341 29659 1353
rect 29601 1289 29604 1341
rect 29656 1289 29659 1341
rect 29601 1277 29613 1289
rect 29647 1277 29659 1289
rect 29601 1225 29604 1277
rect 29656 1225 29659 1277
rect 29601 1213 29613 1225
rect 29647 1213 29659 1225
rect 29601 1161 29604 1213
rect 29656 1161 29659 1213
rect 29601 1147 29659 1161
rect 29700 3133 29752 3147
rect 29700 3069 29709 3081
rect 29743 3069 29752 3081
rect 29700 3005 29709 3017
rect 29743 3005 29752 3017
rect 29700 2941 29709 2953
rect 29743 2941 29752 2953
rect 29700 2884 29752 2889
rect 29700 2877 29709 2884
rect 29743 2877 29752 2884
rect 29700 2813 29752 2825
rect 29700 2749 29752 2761
rect 29700 2685 29752 2697
rect 29700 2621 29752 2633
rect 29700 2562 29709 2569
rect 29743 2562 29752 2569
rect 29700 2557 29752 2562
rect 29700 2493 29709 2505
rect 29743 2493 29752 2505
rect 29700 2429 29709 2441
rect 29743 2429 29752 2441
rect 29700 2365 29709 2377
rect 29743 2365 29752 2377
rect 29700 2308 29752 2313
rect 29700 2301 29709 2308
rect 29743 2301 29752 2308
rect 29700 2237 29752 2249
rect 29700 2173 29752 2185
rect 29700 2109 29752 2121
rect 29700 2045 29752 2057
rect 29700 1986 29709 1993
rect 29743 1986 29752 1993
rect 29700 1981 29752 1986
rect 29700 1917 29709 1929
rect 29743 1917 29752 1929
rect 29700 1853 29709 1865
rect 29743 1853 29752 1865
rect 29700 1789 29709 1801
rect 29743 1789 29752 1801
rect 29700 1732 29752 1737
rect 29700 1725 29709 1732
rect 29743 1725 29752 1732
rect 29700 1661 29752 1673
rect 29700 1597 29752 1609
rect 29700 1533 29752 1545
rect 29700 1469 29752 1481
rect 29700 1410 29709 1417
rect 29743 1410 29752 1417
rect 29700 1405 29752 1410
rect 29700 1341 29709 1353
rect 29743 1341 29752 1353
rect 29700 1277 29709 1289
rect 29743 1277 29752 1289
rect 29700 1213 29709 1225
rect 29743 1213 29752 1225
rect 29700 1147 29752 1161
rect 29793 3133 29851 3147
rect 29793 3081 29796 3133
rect 29848 3081 29851 3133
rect 29793 3069 29805 3081
rect 29839 3069 29851 3081
rect 29793 3017 29796 3069
rect 29848 3017 29851 3069
rect 29793 3005 29805 3017
rect 29839 3005 29851 3017
rect 29793 2953 29796 3005
rect 29848 2953 29851 3005
rect 29793 2941 29805 2953
rect 29839 2941 29851 2953
rect 29793 2889 29796 2941
rect 29848 2889 29851 2941
rect 29793 2884 29851 2889
rect 29793 2877 29805 2884
rect 29839 2877 29851 2884
rect 29793 2825 29796 2877
rect 29848 2825 29851 2877
rect 29793 2813 29851 2825
rect 29793 2761 29796 2813
rect 29848 2761 29851 2813
rect 29793 2749 29851 2761
rect 29793 2697 29796 2749
rect 29848 2697 29851 2749
rect 29793 2685 29851 2697
rect 29793 2633 29796 2685
rect 29848 2633 29851 2685
rect 29793 2621 29851 2633
rect 29793 2569 29796 2621
rect 29848 2569 29851 2621
rect 29793 2562 29805 2569
rect 29839 2562 29851 2569
rect 29793 2557 29851 2562
rect 29793 2505 29796 2557
rect 29848 2505 29851 2557
rect 29793 2493 29805 2505
rect 29839 2493 29851 2505
rect 29793 2441 29796 2493
rect 29848 2441 29851 2493
rect 29793 2429 29805 2441
rect 29839 2429 29851 2441
rect 29793 2377 29796 2429
rect 29848 2377 29851 2429
rect 29793 2365 29805 2377
rect 29839 2365 29851 2377
rect 29793 2313 29796 2365
rect 29848 2313 29851 2365
rect 29793 2308 29851 2313
rect 29793 2301 29805 2308
rect 29839 2301 29851 2308
rect 29793 2249 29796 2301
rect 29848 2249 29851 2301
rect 29793 2237 29851 2249
rect 29793 2185 29796 2237
rect 29848 2185 29851 2237
rect 29793 2173 29851 2185
rect 29793 2121 29796 2173
rect 29848 2121 29851 2173
rect 29793 2109 29851 2121
rect 29793 2057 29796 2109
rect 29848 2057 29851 2109
rect 29793 2045 29851 2057
rect 29793 1993 29796 2045
rect 29848 1993 29851 2045
rect 29793 1986 29805 1993
rect 29839 1986 29851 1993
rect 29793 1981 29851 1986
rect 29793 1929 29796 1981
rect 29848 1929 29851 1981
rect 29793 1917 29805 1929
rect 29839 1917 29851 1929
rect 29793 1865 29796 1917
rect 29848 1865 29851 1917
rect 29793 1853 29805 1865
rect 29839 1853 29851 1865
rect 29793 1801 29796 1853
rect 29848 1801 29851 1853
rect 29793 1789 29805 1801
rect 29839 1789 29851 1801
rect 29793 1737 29796 1789
rect 29848 1737 29851 1789
rect 29793 1732 29851 1737
rect 29793 1725 29805 1732
rect 29839 1725 29851 1732
rect 29793 1673 29796 1725
rect 29848 1673 29851 1725
rect 29793 1661 29851 1673
rect 29793 1609 29796 1661
rect 29848 1609 29851 1661
rect 29793 1597 29851 1609
rect 29793 1545 29796 1597
rect 29848 1545 29851 1597
rect 29793 1533 29851 1545
rect 29793 1481 29796 1533
rect 29848 1481 29851 1533
rect 29793 1469 29851 1481
rect 29793 1417 29796 1469
rect 29848 1417 29851 1469
rect 29793 1410 29805 1417
rect 29839 1410 29851 1417
rect 29793 1405 29851 1410
rect 29793 1353 29796 1405
rect 29848 1353 29851 1405
rect 29793 1341 29805 1353
rect 29839 1341 29851 1353
rect 29793 1289 29796 1341
rect 29848 1289 29851 1341
rect 29793 1277 29805 1289
rect 29839 1277 29851 1289
rect 29793 1225 29796 1277
rect 29848 1225 29851 1277
rect 29793 1213 29805 1225
rect 29839 1213 29851 1225
rect 29793 1161 29796 1213
rect 29848 1161 29851 1213
rect 29793 1147 29851 1161
rect 29889 3133 29947 3147
rect 29889 3081 29892 3133
rect 29944 3081 29947 3133
rect 29889 3069 29901 3081
rect 29935 3069 29947 3081
rect 29889 3017 29892 3069
rect 29944 3017 29947 3069
rect 29889 3005 29901 3017
rect 29935 3005 29947 3017
rect 29889 2953 29892 3005
rect 29944 2953 29947 3005
rect 29889 2941 29901 2953
rect 29935 2941 29947 2953
rect 29889 2889 29892 2941
rect 29944 2889 29947 2941
rect 29889 2884 29947 2889
rect 29889 2877 29901 2884
rect 29935 2877 29947 2884
rect 29889 2825 29892 2877
rect 29944 2825 29947 2877
rect 29889 2813 29947 2825
rect 29889 2761 29892 2813
rect 29944 2761 29947 2813
rect 29889 2749 29947 2761
rect 29889 2697 29892 2749
rect 29944 2697 29947 2749
rect 29889 2685 29947 2697
rect 29889 2633 29892 2685
rect 29944 2633 29947 2685
rect 29889 2621 29947 2633
rect 29889 2569 29892 2621
rect 29944 2569 29947 2621
rect 29889 2562 29901 2569
rect 29935 2562 29947 2569
rect 29889 2557 29947 2562
rect 29889 2505 29892 2557
rect 29944 2505 29947 2557
rect 29889 2493 29901 2505
rect 29935 2493 29947 2505
rect 29889 2441 29892 2493
rect 29944 2441 29947 2493
rect 29889 2429 29901 2441
rect 29935 2429 29947 2441
rect 29889 2377 29892 2429
rect 29944 2377 29947 2429
rect 29889 2365 29901 2377
rect 29935 2365 29947 2377
rect 29889 2313 29892 2365
rect 29944 2313 29947 2365
rect 29889 2308 29947 2313
rect 29889 2301 29901 2308
rect 29935 2301 29947 2308
rect 29889 2249 29892 2301
rect 29944 2249 29947 2301
rect 29889 2237 29947 2249
rect 29889 2185 29892 2237
rect 29944 2185 29947 2237
rect 29889 2173 29947 2185
rect 29889 2121 29892 2173
rect 29944 2121 29947 2173
rect 29889 2109 29947 2121
rect 29889 2057 29892 2109
rect 29944 2057 29947 2109
rect 29889 2045 29947 2057
rect 29889 1993 29892 2045
rect 29944 1993 29947 2045
rect 29889 1986 29901 1993
rect 29935 1986 29947 1993
rect 29889 1981 29947 1986
rect 29889 1929 29892 1981
rect 29944 1929 29947 1981
rect 29889 1917 29901 1929
rect 29935 1917 29947 1929
rect 29889 1865 29892 1917
rect 29944 1865 29947 1917
rect 29889 1853 29901 1865
rect 29935 1853 29947 1865
rect 29889 1801 29892 1853
rect 29944 1801 29947 1853
rect 29889 1789 29901 1801
rect 29935 1789 29947 1801
rect 29889 1737 29892 1789
rect 29944 1737 29947 1789
rect 29889 1732 29947 1737
rect 29889 1725 29901 1732
rect 29935 1725 29947 1732
rect 29889 1673 29892 1725
rect 29944 1673 29947 1725
rect 29889 1661 29947 1673
rect 29889 1609 29892 1661
rect 29944 1609 29947 1661
rect 29889 1597 29947 1609
rect 29889 1545 29892 1597
rect 29944 1545 29947 1597
rect 29889 1533 29947 1545
rect 29889 1481 29892 1533
rect 29944 1481 29947 1533
rect 29889 1469 29947 1481
rect 29889 1417 29892 1469
rect 29944 1417 29947 1469
rect 29889 1410 29901 1417
rect 29935 1410 29947 1417
rect 29889 1405 29947 1410
rect 29889 1353 29892 1405
rect 29944 1353 29947 1405
rect 29889 1341 29901 1353
rect 29935 1341 29947 1353
rect 29889 1289 29892 1341
rect 29944 1289 29947 1341
rect 29889 1277 29901 1289
rect 29935 1277 29947 1289
rect 29889 1225 29892 1277
rect 29944 1225 29947 1277
rect 29889 1213 29901 1225
rect 29935 1213 29947 1225
rect 29889 1161 29892 1213
rect 29944 1161 29947 1213
rect 29889 1147 29947 1161
rect 29985 3133 30043 3147
rect 29985 3081 29988 3133
rect 30040 3081 30043 3133
rect 29985 3069 29997 3081
rect 30031 3069 30043 3081
rect 29985 3017 29988 3069
rect 30040 3017 30043 3069
rect 29985 3005 29997 3017
rect 30031 3005 30043 3017
rect 29985 2953 29988 3005
rect 30040 2953 30043 3005
rect 29985 2941 29997 2953
rect 30031 2941 30043 2953
rect 29985 2889 29988 2941
rect 30040 2889 30043 2941
rect 29985 2884 30043 2889
rect 29985 2877 29997 2884
rect 30031 2877 30043 2884
rect 29985 2825 29988 2877
rect 30040 2825 30043 2877
rect 29985 2813 30043 2825
rect 29985 2761 29988 2813
rect 30040 2761 30043 2813
rect 29985 2749 30043 2761
rect 29985 2697 29988 2749
rect 30040 2697 30043 2749
rect 29985 2685 30043 2697
rect 29985 2633 29988 2685
rect 30040 2633 30043 2685
rect 29985 2621 30043 2633
rect 29985 2569 29988 2621
rect 30040 2569 30043 2621
rect 29985 2562 29997 2569
rect 30031 2562 30043 2569
rect 29985 2557 30043 2562
rect 29985 2505 29988 2557
rect 30040 2505 30043 2557
rect 29985 2493 29997 2505
rect 30031 2493 30043 2505
rect 29985 2441 29988 2493
rect 30040 2441 30043 2493
rect 29985 2429 29997 2441
rect 30031 2429 30043 2441
rect 29985 2377 29988 2429
rect 30040 2377 30043 2429
rect 29985 2365 29997 2377
rect 30031 2365 30043 2377
rect 29985 2313 29988 2365
rect 30040 2313 30043 2365
rect 29985 2308 30043 2313
rect 29985 2301 29997 2308
rect 30031 2301 30043 2308
rect 29985 2249 29988 2301
rect 30040 2249 30043 2301
rect 29985 2237 30043 2249
rect 29985 2185 29988 2237
rect 30040 2185 30043 2237
rect 29985 2173 30043 2185
rect 29985 2121 29988 2173
rect 30040 2121 30043 2173
rect 29985 2109 30043 2121
rect 29985 2057 29988 2109
rect 30040 2057 30043 2109
rect 29985 2045 30043 2057
rect 29985 1993 29988 2045
rect 30040 1993 30043 2045
rect 29985 1986 29997 1993
rect 30031 1986 30043 1993
rect 29985 1981 30043 1986
rect 29985 1929 29988 1981
rect 30040 1929 30043 1981
rect 29985 1917 29997 1929
rect 30031 1917 30043 1929
rect 29985 1865 29988 1917
rect 30040 1865 30043 1917
rect 29985 1853 29997 1865
rect 30031 1853 30043 1865
rect 29985 1801 29988 1853
rect 30040 1801 30043 1853
rect 29985 1789 29997 1801
rect 30031 1789 30043 1801
rect 29985 1737 29988 1789
rect 30040 1737 30043 1789
rect 29985 1732 30043 1737
rect 29985 1725 29997 1732
rect 30031 1725 30043 1732
rect 29985 1673 29988 1725
rect 30040 1673 30043 1725
rect 29985 1661 30043 1673
rect 29985 1609 29988 1661
rect 30040 1609 30043 1661
rect 29985 1597 30043 1609
rect 29985 1545 29988 1597
rect 30040 1545 30043 1597
rect 29985 1533 30043 1545
rect 29985 1481 29988 1533
rect 30040 1481 30043 1533
rect 29985 1469 30043 1481
rect 29985 1417 29988 1469
rect 30040 1417 30043 1469
rect 29985 1410 29997 1417
rect 30031 1410 30043 1417
rect 29985 1405 30043 1410
rect 29985 1353 29988 1405
rect 30040 1353 30043 1405
rect 29985 1341 29997 1353
rect 30031 1341 30043 1353
rect 29985 1289 29988 1341
rect 30040 1289 30043 1341
rect 29985 1277 29997 1289
rect 30031 1277 30043 1289
rect 29985 1225 29988 1277
rect 30040 1225 30043 1277
rect 29985 1213 29997 1225
rect 30031 1213 30043 1225
rect 29985 1161 29988 1213
rect 30040 1161 30043 1213
rect 29985 1147 30043 1161
rect 30084 3133 30136 3147
rect 30084 3069 30093 3081
rect 30127 3069 30136 3081
rect 30084 3005 30093 3017
rect 30127 3005 30136 3017
rect 30084 2941 30093 2953
rect 30127 2941 30136 2953
rect 30084 2884 30136 2889
rect 30084 2877 30093 2884
rect 30127 2877 30136 2884
rect 30084 2813 30136 2825
rect 30084 2749 30136 2761
rect 30084 2685 30136 2697
rect 30084 2621 30136 2633
rect 30084 2562 30093 2569
rect 30127 2562 30136 2569
rect 30084 2557 30136 2562
rect 30084 2493 30093 2505
rect 30127 2493 30136 2505
rect 30084 2429 30093 2441
rect 30127 2429 30136 2441
rect 30084 2365 30093 2377
rect 30127 2365 30136 2377
rect 30084 2308 30136 2313
rect 30084 2301 30093 2308
rect 30127 2301 30136 2308
rect 30084 2237 30136 2249
rect 30084 2173 30136 2185
rect 30084 2109 30136 2121
rect 30084 2045 30136 2057
rect 30084 1986 30093 1993
rect 30127 1986 30136 1993
rect 30084 1981 30136 1986
rect 30084 1917 30093 1929
rect 30127 1917 30136 1929
rect 30084 1853 30093 1865
rect 30127 1853 30136 1865
rect 30084 1789 30093 1801
rect 30127 1789 30136 1801
rect 30084 1732 30136 1737
rect 30084 1725 30093 1732
rect 30127 1725 30136 1732
rect 30084 1661 30136 1673
rect 30084 1597 30136 1609
rect 30084 1533 30136 1545
rect 30084 1469 30136 1481
rect 30084 1410 30093 1417
rect 30127 1410 30136 1417
rect 30084 1405 30136 1410
rect 30084 1341 30093 1353
rect 30127 1341 30136 1353
rect 30084 1277 30093 1289
rect 30127 1277 30136 1289
rect 30084 1213 30093 1225
rect 30127 1213 30136 1225
rect 30084 1147 30136 1161
rect 30177 3133 30235 3147
rect 30177 3081 30180 3133
rect 30232 3081 30235 3133
rect 30177 3069 30189 3081
rect 30223 3069 30235 3081
rect 30177 3017 30180 3069
rect 30232 3017 30235 3069
rect 30177 3005 30189 3017
rect 30223 3005 30235 3017
rect 30177 2953 30180 3005
rect 30232 2953 30235 3005
rect 30177 2941 30189 2953
rect 30223 2941 30235 2953
rect 30177 2889 30180 2941
rect 30232 2889 30235 2941
rect 30177 2884 30235 2889
rect 30177 2877 30189 2884
rect 30223 2877 30235 2884
rect 30177 2825 30180 2877
rect 30232 2825 30235 2877
rect 30177 2813 30235 2825
rect 30177 2761 30180 2813
rect 30232 2761 30235 2813
rect 30177 2749 30235 2761
rect 30177 2697 30180 2749
rect 30232 2697 30235 2749
rect 30177 2685 30235 2697
rect 30177 2633 30180 2685
rect 30232 2633 30235 2685
rect 30177 2621 30235 2633
rect 30177 2569 30180 2621
rect 30232 2569 30235 2621
rect 30177 2562 30189 2569
rect 30223 2562 30235 2569
rect 30177 2557 30235 2562
rect 30177 2505 30180 2557
rect 30232 2505 30235 2557
rect 30177 2493 30189 2505
rect 30223 2493 30235 2505
rect 30177 2441 30180 2493
rect 30232 2441 30235 2493
rect 30177 2429 30189 2441
rect 30223 2429 30235 2441
rect 30177 2377 30180 2429
rect 30232 2377 30235 2429
rect 30177 2365 30189 2377
rect 30223 2365 30235 2377
rect 30177 2313 30180 2365
rect 30232 2313 30235 2365
rect 30177 2308 30235 2313
rect 30177 2301 30189 2308
rect 30223 2301 30235 2308
rect 30177 2249 30180 2301
rect 30232 2249 30235 2301
rect 30177 2237 30235 2249
rect 30177 2185 30180 2237
rect 30232 2185 30235 2237
rect 30177 2173 30235 2185
rect 30177 2121 30180 2173
rect 30232 2121 30235 2173
rect 30177 2109 30235 2121
rect 30177 2057 30180 2109
rect 30232 2057 30235 2109
rect 30177 2045 30235 2057
rect 30177 1993 30180 2045
rect 30232 1993 30235 2045
rect 30177 1986 30189 1993
rect 30223 1986 30235 1993
rect 30177 1981 30235 1986
rect 30177 1929 30180 1981
rect 30232 1929 30235 1981
rect 30177 1917 30189 1929
rect 30223 1917 30235 1929
rect 30177 1865 30180 1917
rect 30232 1865 30235 1917
rect 30177 1853 30189 1865
rect 30223 1853 30235 1865
rect 30177 1801 30180 1853
rect 30232 1801 30235 1853
rect 30177 1789 30189 1801
rect 30223 1789 30235 1801
rect 30177 1737 30180 1789
rect 30232 1737 30235 1789
rect 30177 1732 30235 1737
rect 30177 1725 30189 1732
rect 30223 1725 30235 1732
rect 30177 1673 30180 1725
rect 30232 1673 30235 1725
rect 30177 1661 30235 1673
rect 30177 1609 30180 1661
rect 30232 1609 30235 1661
rect 30177 1597 30235 1609
rect 30177 1545 30180 1597
rect 30232 1545 30235 1597
rect 30177 1533 30235 1545
rect 30177 1481 30180 1533
rect 30232 1481 30235 1533
rect 30177 1469 30235 1481
rect 30177 1417 30180 1469
rect 30232 1417 30235 1469
rect 30177 1410 30189 1417
rect 30223 1410 30235 1417
rect 30177 1405 30235 1410
rect 30177 1353 30180 1405
rect 30232 1353 30235 1405
rect 30177 1341 30189 1353
rect 30223 1341 30235 1353
rect 30177 1289 30180 1341
rect 30232 1289 30235 1341
rect 30177 1277 30189 1289
rect 30223 1277 30235 1289
rect 30177 1225 30180 1277
rect 30232 1225 30235 1277
rect 30177 1213 30189 1225
rect 30223 1213 30235 1225
rect 30177 1161 30180 1213
rect 30232 1161 30235 1213
rect 30177 1147 30235 1161
rect 30273 3133 30331 3147
rect 30273 3081 30276 3133
rect 30328 3081 30331 3133
rect 30273 3069 30285 3081
rect 30319 3069 30331 3081
rect 30273 3017 30276 3069
rect 30328 3017 30331 3069
rect 30273 3005 30285 3017
rect 30319 3005 30331 3017
rect 30273 2953 30276 3005
rect 30328 2953 30331 3005
rect 30273 2941 30285 2953
rect 30319 2941 30331 2953
rect 30273 2889 30276 2941
rect 30328 2889 30331 2941
rect 30273 2884 30331 2889
rect 30273 2877 30285 2884
rect 30319 2877 30331 2884
rect 30273 2825 30276 2877
rect 30328 2825 30331 2877
rect 30273 2813 30331 2825
rect 30273 2761 30276 2813
rect 30328 2761 30331 2813
rect 30273 2749 30331 2761
rect 30273 2697 30276 2749
rect 30328 2697 30331 2749
rect 30273 2685 30331 2697
rect 30273 2633 30276 2685
rect 30328 2633 30331 2685
rect 30273 2621 30331 2633
rect 30273 2569 30276 2621
rect 30328 2569 30331 2621
rect 30273 2562 30285 2569
rect 30319 2562 30331 2569
rect 30273 2557 30331 2562
rect 30273 2505 30276 2557
rect 30328 2505 30331 2557
rect 30273 2493 30285 2505
rect 30319 2493 30331 2505
rect 30273 2441 30276 2493
rect 30328 2441 30331 2493
rect 30273 2429 30285 2441
rect 30319 2429 30331 2441
rect 30273 2377 30276 2429
rect 30328 2377 30331 2429
rect 30273 2365 30285 2377
rect 30319 2365 30331 2377
rect 30273 2313 30276 2365
rect 30328 2313 30331 2365
rect 30273 2308 30331 2313
rect 30273 2301 30285 2308
rect 30319 2301 30331 2308
rect 30273 2249 30276 2301
rect 30328 2249 30331 2301
rect 30273 2237 30331 2249
rect 30273 2185 30276 2237
rect 30328 2185 30331 2237
rect 30273 2173 30331 2185
rect 30273 2121 30276 2173
rect 30328 2121 30331 2173
rect 30273 2109 30331 2121
rect 30273 2057 30276 2109
rect 30328 2057 30331 2109
rect 30273 2045 30331 2057
rect 30273 1993 30276 2045
rect 30328 1993 30331 2045
rect 30273 1986 30285 1993
rect 30319 1986 30331 1993
rect 30273 1981 30331 1986
rect 30273 1929 30276 1981
rect 30328 1929 30331 1981
rect 30273 1917 30285 1929
rect 30319 1917 30331 1929
rect 30273 1865 30276 1917
rect 30328 1865 30331 1917
rect 30273 1853 30285 1865
rect 30319 1853 30331 1865
rect 30273 1801 30276 1853
rect 30328 1801 30331 1853
rect 30273 1789 30285 1801
rect 30319 1789 30331 1801
rect 30273 1737 30276 1789
rect 30328 1737 30331 1789
rect 30273 1732 30331 1737
rect 30273 1725 30285 1732
rect 30319 1725 30331 1732
rect 30273 1673 30276 1725
rect 30328 1673 30331 1725
rect 30273 1661 30331 1673
rect 30273 1609 30276 1661
rect 30328 1609 30331 1661
rect 30273 1597 30331 1609
rect 30273 1545 30276 1597
rect 30328 1545 30331 1597
rect 30273 1533 30331 1545
rect 30273 1481 30276 1533
rect 30328 1481 30331 1533
rect 30273 1469 30331 1481
rect 30273 1417 30276 1469
rect 30328 1417 30331 1469
rect 30273 1410 30285 1417
rect 30319 1410 30331 1417
rect 30273 1405 30331 1410
rect 30273 1353 30276 1405
rect 30328 1353 30331 1405
rect 30273 1341 30285 1353
rect 30319 1341 30331 1353
rect 30273 1289 30276 1341
rect 30328 1289 30331 1341
rect 30273 1277 30285 1289
rect 30319 1277 30331 1289
rect 30273 1225 30276 1277
rect 30328 1225 30331 1277
rect 30273 1213 30285 1225
rect 30319 1213 30331 1225
rect 30273 1161 30276 1213
rect 30328 1161 30331 1213
rect 30273 1147 30331 1161
rect 30369 3133 30427 3147
rect 30369 3081 30372 3133
rect 30424 3081 30427 3133
rect 30369 3069 30381 3081
rect 30415 3069 30427 3081
rect 30369 3017 30372 3069
rect 30424 3017 30427 3069
rect 30369 3005 30381 3017
rect 30415 3005 30427 3017
rect 30369 2953 30372 3005
rect 30424 2953 30427 3005
rect 30369 2941 30381 2953
rect 30415 2941 30427 2953
rect 30369 2889 30372 2941
rect 30424 2889 30427 2941
rect 30369 2884 30427 2889
rect 30369 2877 30381 2884
rect 30415 2877 30427 2884
rect 30369 2825 30372 2877
rect 30424 2825 30427 2877
rect 30369 2813 30427 2825
rect 30369 2761 30372 2813
rect 30424 2761 30427 2813
rect 30369 2749 30427 2761
rect 30369 2697 30372 2749
rect 30424 2697 30427 2749
rect 30369 2685 30427 2697
rect 30369 2633 30372 2685
rect 30424 2633 30427 2685
rect 30369 2621 30427 2633
rect 30369 2569 30372 2621
rect 30424 2569 30427 2621
rect 30369 2562 30381 2569
rect 30415 2562 30427 2569
rect 30369 2557 30427 2562
rect 30369 2505 30372 2557
rect 30424 2505 30427 2557
rect 30369 2493 30381 2505
rect 30415 2493 30427 2505
rect 30369 2441 30372 2493
rect 30424 2441 30427 2493
rect 30369 2429 30381 2441
rect 30415 2429 30427 2441
rect 30369 2377 30372 2429
rect 30424 2377 30427 2429
rect 30369 2365 30381 2377
rect 30415 2365 30427 2377
rect 30369 2313 30372 2365
rect 30424 2313 30427 2365
rect 30369 2308 30427 2313
rect 30369 2301 30381 2308
rect 30415 2301 30427 2308
rect 30369 2249 30372 2301
rect 30424 2249 30427 2301
rect 30369 2237 30427 2249
rect 30369 2185 30372 2237
rect 30424 2185 30427 2237
rect 30369 2173 30427 2185
rect 30369 2121 30372 2173
rect 30424 2121 30427 2173
rect 30369 2109 30427 2121
rect 30369 2057 30372 2109
rect 30424 2057 30427 2109
rect 30369 2045 30427 2057
rect 30369 1993 30372 2045
rect 30424 1993 30427 2045
rect 30369 1986 30381 1993
rect 30415 1986 30427 1993
rect 30369 1981 30427 1986
rect 30369 1929 30372 1981
rect 30424 1929 30427 1981
rect 30369 1917 30381 1929
rect 30415 1917 30427 1929
rect 30369 1865 30372 1917
rect 30424 1865 30427 1917
rect 30369 1853 30381 1865
rect 30415 1853 30427 1865
rect 30369 1801 30372 1853
rect 30424 1801 30427 1853
rect 30369 1789 30381 1801
rect 30415 1789 30427 1801
rect 30369 1737 30372 1789
rect 30424 1737 30427 1789
rect 30369 1732 30427 1737
rect 30369 1725 30381 1732
rect 30415 1725 30427 1732
rect 30369 1673 30372 1725
rect 30424 1673 30427 1725
rect 30369 1661 30427 1673
rect 30369 1609 30372 1661
rect 30424 1609 30427 1661
rect 30369 1597 30427 1609
rect 30369 1545 30372 1597
rect 30424 1545 30427 1597
rect 30369 1533 30427 1545
rect 30369 1481 30372 1533
rect 30424 1481 30427 1533
rect 30369 1469 30427 1481
rect 30369 1417 30372 1469
rect 30424 1417 30427 1469
rect 30369 1410 30381 1417
rect 30415 1410 30427 1417
rect 30369 1405 30427 1410
rect 30369 1353 30372 1405
rect 30424 1353 30427 1405
rect 30369 1341 30381 1353
rect 30415 1341 30427 1353
rect 30369 1289 30372 1341
rect 30424 1289 30427 1341
rect 30369 1277 30381 1289
rect 30415 1277 30427 1289
rect 30369 1225 30372 1277
rect 30424 1225 30427 1277
rect 30369 1213 30381 1225
rect 30415 1213 30427 1225
rect 30369 1161 30372 1213
rect 30424 1161 30427 1213
rect 30369 1147 30427 1161
rect 30468 3133 30520 3147
rect 30468 3069 30477 3081
rect 30511 3069 30520 3081
rect 30468 3005 30477 3017
rect 30511 3005 30520 3017
rect 30468 2941 30477 2953
rect 30511 2941 30520 2953
rect 30468 2884 30520 2889
rect 30468 2877 30477 2884
rect 30511 2877 30520 2884
rect 30468 2813 30520 2825
rect 30468 2749 30520 2761
rect 30468 2685 30520 2697
rect 30468 2621 30520 2633
rect 30468 2562 30477 2569
rect 30511 2562 30520 2569
rect 30468 2557 30520 2562
rect 30468 2493 30477 2505
rect 30511 2493 30520 2505
rect 30468 2429 30477 2441
rect 30511 2429 30520 2441
rect 30468 2365 30477 2377
rect 30511 2365 30520 2377
rect 30468 2308 30520 2313
rect 30468 2301 30477 2308
rect 30511 2301 30520 2308
rect 30468 2237 30520 2249
rect 30468 2173 30520 2185
rect 30468 2109 30520 2121
rect 30468 2045 30520 2057
rect 30468 1986 30477 1993
rect 30511 1986 30520 1993
rect 30468 1981 30520 1986
rect 30468 1917 30477 1929
rect 30511 1917 30520 1929
rect 30468 1853 30477 1865
rect 30511 1853 30520 1865
rect 30468 1789 30477 1801
rect 30511 1789 30520 1801
rect 30468 1732 30520 1737
rect 30468 1725 30477 1732
rect 30511 1725 30520 1732
rect 30468 1661 30520 1673
rect 30468 1597 30520 1609
rect 30468 1533 30520 1545
rect 30468 1469 30520 1481
rect 30468 1410 30477 1417
rect 30511 1410 30520 1417
rect 30468 1405 30520 1410
rect 30468 1341 30477 1353
rect 30511 1341 30520 1353
rect 30468 1277 30477 1289
rect 30511 1277 30520 1289
rect 30468 1213 30477 1225
rect 30511 1213 30520 1225
rect 30468 1147 30520 1161
rect 30561 3133 30619 3147
rect 30561 3081 30564 3133
rect 30616 3081 30619 3133
rect 30561 3069 30573 3081
rect 30607 3069 30619 3081
rect 30561 3017 30564 3069
rect 30616 3017 30619 3069
rect 30561 3005 30573 3017
rect 30607 3005 30619 3017
rect 30561 2953 30564 3005
rect 30616 2953 30619 3005
rect 30561 2941 30573 2953
rect 30607 2941 30619 2953
rect 30561 2889 30564 2941
rect 30616 2889 30619 2941
rect 30561 2884 30619 2889
rect 30561 2877 30573 2884
rect 30607 2877 30619 2884
rect 30561 2825 30564 2877
rect 30616 2825 30619 2877
rect 30561 2813 30619 2825
rect 30561 2761 30564 2813
rect 30616 2761 30619 2813
rect 30561 2749 30619 2761
rect 30561 2697 30564 2749
rect 30616 2697 30619 2749
rect 30561 2685 30619 2697
rect 30561 2633 30564 2685
rect 30616 2633 30619 2685
rect 30561 2621 30619 2633
rect 30561 2569 30564 2621
rect 30616 2569 30619 2621
rect 30561 2562 30573 2569
rect 30607 2562 30619 2569
rect 30561 2557 30619 2562
rect 30561 2505 30564 2557
rect 30616 2505 30619 2557
rect 30561 2493 30573 2505
rect 30607 2493 30619 2505
rect 30561 2441 30564 2493
rect 30616 2441 30619 2493
rect 30561 2429 30573 2441
rect 30607 2429 30619 2441
rect 30561 2377 30564 2429
rect 30616 2377 30619 2429
rect 30561 2365 30573 2377
rect 30607 2365 30619 2377
rect 30561 2313 30564 2365
rect 30616 2313 30619 2365
rect 30561 2308 30619 2313
rect 30561 2301 30573 2308
rect 30607 2301 30619 2308
rect 30561 2249 30564 2301
rect 30616 2249 30619 2301
rect 30561 2237 30619 2249
rect 30561 2185 30564 2237
rect 30616 2185 30619 2237
rect 30561 2173 30619 2185
rect 30561 2121 30564 2173
rect 30616 2121 30619 2173
rect 30561 2109 30619 2121
rect 30561 2057 30564 2109
rect 30616 2057 30619 2109
rect 30561 2045 30619 2057
rect 30561 1993 30564 2045
rect 30616 1993 30619 2045
rect 30561 1986 30573 1993
rect 30607 1986 30619 1993
rect 30561 1981 30619 1986
rect 30561 1929 30564 1981
rect 30616 1929 30619 1981
rect 30561 1917 30573 1929
rect 30607 1917 30619 1929
rect 30561 1865 30564 1917
rect 30616 1865 30619 1917
rect 30561 1853 30573 1865
rect 30607 1853 30619 1865
rect 30561 1801 30564 1853
rect 30616 1801 30619 1853
rect 30561 1789 30573 1801
rect 30607 1789 30619 1801
rect 30561 1737 30564 1789
rect 30616 1737 30619 1789
rect 30561 1732 30619 1737
rect 30561 1725 30573 1732
rect 30607 1725 30619 1732
rect 30561 1673 30564 1725
rect 30616 1673 30619 1725
rect 30561 1661 30619 1673
rect 30561 1609 30564 1661
rect 30616 1609 30619 1661
rect 30561 1597 30619 1609
rect 30561 1545 30564 1597
rect 30616 1545 30619 1597
rect 30561 1533 30619 1545
rect 30561 1481 30564 1533
rect 30616 1481 30619 1533
rect 30561 1469 30619 1481
rect 30561 1417 30564 1469
rect 30616 1417 30619 1469
rect 30561 1410 30573 1417
rect 30607 1410 30619 1417
rect 30561 1405 30619 1410
rect 30561 1353 30564 1405
rect 30616 1353 30619 1405
rect 30561 1341 30573 1353
rect 30607 1341 30619 1353
rect 30561 1289 30564 1341
rect 30616 1289 30619 1341
rect 30561 1277 30573 1289
rect 30607 1277 30619 1289
rect 30561 1225 30564 1277
rect 30616 1225 30619 1277
rect 30561 1213 30573 1225
rect 30607 1213 30619 1225
rect 30561 1161 30564 1213
rect 30616 1161 30619 1213
rect 30561 1147 30619 1161
rect 30657 3133 30715 3147
rect 30657 3081 30660 3133
rect 30712 3081 30715 3133
rect 30657 3069 30669 3081
rect 30703 3069 30715 3081
rect 30657 3017 30660 3069
rect 30712 3017 30715 3069
rect 30657 3005 30669 3017
rect 30703 3005 30715 3017
rect 30657 2953 30660 3005
rect 30712 2953 30715 3005
rect 30657 2941 30669 2953
rect 30703 2941 30715 2953
rect 30657 2889 30660 2941
rect 30712 2889 30715 2941
rect 30657 2884 30715 2889
rect 30657 2877 30669 2884
rect 30703 2877 30715 2884
rect 30657 2825 30660 2877
rect 30712 2825 30715 2877
rect 30657 2813 30715 2825
rect 30657 2761 30660 2813
rect 30712 2761 30715 2813
rect 30657 2749 30715 2761
rect 30657 2697 30660 2749
rect 30712 2697 30715 2749
rect 30657 2685 30715 2697
rect 30657 2633 30660 2685
rect 30712 2633 30715 2685
rect 30657 2621 30715 2633
rect 30657 2569 30660 2621
rect 30712 2569 30715 2621
rect 30657 2562 30669 2569
rect 30703 2562 30715 2569
rect 30657 2557 30715 2562
rect 30657 2505 30660 2557
rect 30712 2505 30715 2557
rect 30657 2493 30669 2505
rect 30703 2493 30715 2505
rect 30657 2441 30660 2493
rect 30712 2441 30715 2493
rect 30657 2429 30669 2441
rect 30703 2429 30715 2441
rect 30657 2377 30660 2429
rect 30712 2377 30715 2429
rect 30657 2365 30669 2377
rect 30703 2365 30715 2377
rect 30657 2313 30660 2365
rect 30712 2313 30715 2365
rect 30657 2308 30715 2313
rect 30657 2301 30669 2308
rect 30703 2301 30715 2308
rect 30657 2249 30660 2301
rect 30712 2249 30715 2301
rect 30657 2237 30715 2249
rect 30657 2185 30660 2237
rect 30712 2185 30715 2237
rect 30657 2173 30715 2185
rect 30657 2121 30660 2173
rect 30712 2121 30715 2173
rect 30657 2109 30715 2121
rect 30657 2057 30660 2109
rect 30712 2057 30715 2109
rect 30657 2045 30715 2057
rect 30657 1993 30660 2045
rect 30712 1993 30715 2045
rect 30657 1986 30669 1993
rect 30703 1986 30715 1993
rect 30657 1981 30715 1986
rect 30657 1929 30660 1981
rect 30712 1929 30715 1981
rect 30657 1917 30669 1929
rect 30703 1917 30715 1929
rect 30657 1865 30660 1917
rect 30712 1865 30715 1917
rect 30657 1853 30669 1865
rect 30703 1853 30715 1865
rect 30657 1801 30660 1853
rect 30712 1801 30715 1853
rect 30657 1789 30669 1801
rect 30703 1789 30715 1801
rect 30657 1737 30660 1789
rect 30712 1737 30715 1789
rect 30657 1732 30715 1737
rect 30657 1725 30669 1732
rect 30703 1725 30715 1732
rect 30657 1673 30660 1725
rect 30712 1673 30715 1725
rect 30657 1661 30715 1673
rect 30657 1609 30660 1661
rect 30712 1609 30715 1661
rect 30657 1597 30715 1609
rect 30657 1545 30660 1597
rect 30712 1545 30715 1597
rect 30657 1533 30715 1545
rect 30657 1481 30660 1533
rect 30712 1481 30715 1533
rect 30657 1469 30715 1481
rect 30657 1417 30660 1469
rect 30712 1417 30715 1469
rect 30657 1410 30669 1417
rect 30703 1410 30715 1417
rect 30657 1405 30715 1410
rect 30657 1353 30660 1405
rect 30712 1353 30715 1405
rect 30657 1341 30669 1353
rect 30703 1341 30715 1353
rect 30657 1289 30660 1341
rect 30712 1289 30715 1341
rect 30657 1277 30669 1289
rect 30703 1277 30715 1289
rect 30657 1225 30660 1277
rect 30712 1225 30715 1277
rect 30657 1213 30669 1225
rect 30703 1213 30715 1225
rect 30657 1161 30660 1213
rect 30712 1161 30715 1213
rect 30657 1147 30715 1161
rect 30753 3133 30811 3147
rect 30753 3081 30756 3133
rect 30808 3081 30811 3133
rect 30753 3069 30765 3081
rect 30799 3069 30811 3081
rect 30753 3017 30756 3069
rect 30808 3017 30811 3069
rect 30753 3005 30765 3017
rect 30799 3005 30811 3017
rect 30753 2953 30756 3005
rect 30808 2953 30811 3005
rect 30753 2941 30765 2953
rect 30799 2941 30811 2953
rect 30753 2889 30756 2941
rect 30808 2889 30811 2941
rect 30753 2884 30811 2889
rect 30753 2877 30765 2884
rect 30799 2877 30811 2884
rect 30753 2825 30756 2877
rect 30808 2825 30811 2877
rect 30753 2813 30811 2825
rect 30753 2761 30756 2813
rect 30808 2761 30811 2813
rect 30753 2749 30811 2761
rect 30753 2697 30756 2749
rect 30808 2697 30811 2749
rect 30753 2685 30811 2697
rect 30753 2633 30756 2685
rect 30808 2633 30811 2685
rect 30753 2621 30811 2633
rect 30753 2569 30756 2621
rect 30808 2569 30811 2621
rect 30753 2562 30765 2569
rect 30799 2562 30811 2569
rect 30753 2557 30811 2562
rect 30753 2505 30756 2557
rect 30808 2505 30811 2557
rect 30753 2493 30765 2505
rect 30799 2493 30811 2505
rect 30753 2441 30756 2493
rect 30808 2441 30811 2493
rect 30753 2429 30765 2441
rect 30799 2429 30811 2441
rect 30753 2377 30756 2429
rect 30808 2377 30811 2429
rect 30753 2365 30765 2377
rect 30799 2365 30811 2377
rect 30753 2313 30756 2365
rect 30808 2313 30811 2365
rect 30753 2308 30811 2313
rect 30753 2301 30765 2308
rect 30799 2301 30811 2308
rect 30753 2249 30756 2301
rect 30808 2249 30811 2301
rect 30753 2237 30811 2249
rect 30753 2185 30756 2237
rect 30808 2185 30811 2237
rect 30753 2173 30811 2185
rect 30753 2121 30756 2173
rect 30808 2121 30811 2173
rect 30753 2109 30811 2121
rect 30753 2057 30756 2109
rect 30808 2057 30811 2109
rect 30753 2045 30811 2057
rect 30753 1993 30756 2045
rect 30808 1993 30811 2045
rect 30753 1986 30765 1993
rect 30799 1986 30811 1993
rect 30753 1981 30811 1986
rect 30753 1929 30756 1981
rect 30808 1929 30811 1981
rect 30753 1917 30765 1929
rect 30799 1917 30811 1929
rect 30753 1865 30756 1917
rect 30808 1865 30811 1917
rect 30753 1853 30765 1865
rect 30799 1853 30811 1865
rect 30753 1801 30756 1853
rect 30808 1801 30811 1853
rect 30753 1789 30765 1801
rect 30799 1789 30811 1801
rect 30753 1737 30756 1789
rect 30808 1737 30811 1789
rect 30753 1732 30811 1737
rect 30753 1725 30765 1732
rect 30799 1725 30811 1732
rect 30753 1673 30756 1725
rect 30808 1673 30811 1725
rect 30753 1661 30811 1673
rect 30753 1609 30756 1661
rect 30808 1609 30811 1661
rect 30753 1597 30811 1609
rect 30753 1545 30756 1597
rect 30808 1545 30811 1597
rect 30753 1533 30811 1545
rect 30753 1481 30756 1533
rect 30808 1481 30811 1533
rect 30753 1469 30811 1481
rect 30753 1417 30756 1469
rect 30808 1417 30811 1469
rect 30753 1410 30765 1417
rect 30799 1410 30811 1417
rect 30753 1405 30811 1410
rect 30753 1353 30756 1405
rect 30808 1353 30811 1405
rect 30753 1341 30765 1353
rect 30799 1341 30811 1353
rect 30753 1289 30756 1341
rect 30808 1289 30811 1341
rect 30753 1277 30765 1289
rect 30799 1277 30811 1289
rect 30753 1225 30756 1277
rect 30808 1225 30811 1277
rect 30753 1213 30765 1225
rect 30799 1213 30811 1225
rect 30753 1161 30756 1213
rect 30808 1161 30811 1213
rect 30753 1147 30811 1161
rect 30852 3133 30904 3147
rect 30852 3069 30861 3081
rect 30895 3069 30904 3081
rect 30852 3005 30861 3017
rect 30895 3005 30904 3017
rect 30852 2941 30861 2953
rect 30895 2941 30904 2953
rect 30852 2884 30904 2889
rect 30852 2877 30861 2884
rect 30895 2877 30904 2884
rect 30852 2813 30904 2825
rect 30852 2749 30904 2761
rect 30852 2685 30904 2697
rect 30852 2621 30904 2633
rect 30852 2562 30861 2569
rect 30895 2562 30904 2569
rect 30852 2557 30904 2562
rect 30852 2493 30861 2505
rect 30895 2493 30904 2505
rect 30852 2429 30861 2441
rect 30895 2429 30904 2441
rect 30852 2365 30861 2377
rect 30895 2365 30904 2377
rect 30852 2308 30904 2313
rect 30852 2301 30861 2308
rect 30895 2301 30904 2308
rect 30852 2237 30904 2249
rect 30852 2173 30904 2185
rect 30852 2109 30904 2121
rect 30852 2045 30904 2057
rect 30852 1986 30861 1993
rect 30895 1986 30904 1993
rect 30852 1981 30904 1986
rect 30852 1917 30861 1929
rect 30895 1917 30904 1929
rect 30852 1853 30861 1865
rect 30895 1853 30904 1865
rect 30852 1789 30861 1801
rect 30895 1789 30904 1801
rect 30852 1732 30904 1737
rect 30852 1725 30861 1732
rect 30895 1725 30904 1732
rect 30852 1661 30904 1673
rect 30852 1597 30904 1609
rect 30852 1533 30904 1545
rect 30852 1469 30904 1481
rect 30852 1410 30861 1417
rect 30895 1410 30904 1417
rect 30852 1405 30904 1410
rect 30852 1341 30861 1353
rect 30895 1341 30904 1353
rect 30852 1277 30861 1289
rect 30895 1277 30904 1289
rect 30852 1213 30861 1225
rect 30895 1213 30904 1225
rect 30852 1147 30904 1161
rect 30945 3133 31003 3147
rect 30945 3081 30948 3133
rect 31000 3081 31003 3133
rect 30945 3069 30957 3081
rect 30991 3069 31003 3081
rect 30945 3017 30948 3069
rect 31000 3017 31003 3069
rect 30945 3005 30957 3017
rect 30991 3005 31003 3017
rect 30945 2953 30948 3005
rect 31000 2953 31003 3005
rect 30945 2941 30957 2953
rect 30991 2941 31003 2953
rect 30945 2889 30948 2941
rect 31000 2889 31003 2941
rect 30945 2884 31003 2889
rect 30945 2877 30957 2884
rect 30991 2877 31003 2884
rect 30945 2825 30948 2877
rect 31000 2825 31003 2877
rect 30945 2813 31003 2825
rect 30945 2761 30948 2813
rect 31000 2761 31003 2813
rect 30945 2749 31003 2761
rect 30945 2697 30948 2749
rect 31000 2697 31003 2749
rect 30945 2685 31003 2697
rect 30945 2633 30948 2685
rect 31000 2633 31003 2685
rect 30945 2621 31003 2633
rect 30945 2569 30948 2621
rect 31000 2569 31003 2621
rect 30945 2562 30957 2569
rect 30991 2562 31003 2569
rect 30945 2557 31003 2562
rect 30945 2505 30948 2557
rect 31000 2505 31003 2557
rect 30945 2493 30957 2505
rect 30991 2493 31003 2505
rect 30945 2441 30948 2493
rect 31000 2441 31003 2493
rect 30945 2429 30957 2441
rect 30991 2429 31003 2441
rect 30945 2377 30948 2429
rect 31000 2377 31003 2429
rect 30945 2365 30957 2377
rect 30991 2365 31003 2377
rect 30945 2313 30948 2365
rect 31000 2313 31003 2365
rect 30945 2308 31003 2313
rect 30945 2301 30957 2308
rect 30991 2301 31003 2308
rect 30945 2249 30948 2301
rect 31000 2249 31003 2301
rect 30945 2237 31003 2249
rect 30945 2185 30948 2237
rect 31000 2185 31003 2237
rect 30945 2173 31003 2185
rect 30945 2121 30948 2173
rect 31000 2121 31003 2173
rect 30945 2109 31003 2121
rect 30945 2057 30948 2109
rect 31000 2057 31003 2109
rect 30945 2045 31003 2057
rect 30945 1993 30948 2045
rect 31000 1993 31003 2045
rect 30945 1986 30957 1993
rect 30991 1986 31003 1993
rect 30945 1981 31003 1986
rect 30945 1929 30948 1981
rect 31000 1929 31003 1981
rect 30945 1917 30957 1929
rect 30991 1917 31003 1929
rect 30945 1865 30948 1917
rect 31000 1865 31003 1917
rect 30945 1853 30957 1865
rect 30991 1853 31003 1865
rect 30945 1801 30948 1853
rect 31000 1801 31003 1853
rect 30945 1789 30957 1801
rect 30991 1789 31003 1801
rect 30945 1737 30948 1789
rect 31000 1737 31003 1789
rect 30945 1732 31003 1737
rect 30945 1725 30957 1732
rect 30991 1725 31003 1732
rect 30945 1673 30948 1725
rect 31000 1673 31003 1725
rect 30945 1661 31003 1673
rect 30945 1609 30948 1661
rect 31000 1609 31003 1661
rect 30945 1597 31003 1609
rect 30945 1545 30948 1597
rect 31000 1545 31003 1597
rect 30945 1533 31003 1545
rect 30945 1481 30948 1533
rect 31000 1481 31003 1533
rect 30945 1469 31003 1481
rect 30945 1417 30948 1469
rect 31000 1417 31003 1469
rect 30945 1410 30957 1417
rect 30991 1410 31003 1417
rect 30945 1405 31003 1410
rect 30945 1353 30948 1405
rect 31000 1353 31003 1405
rect 30945 1341 30957 1353
rect 30991 1341 31003 1353
rect 30945 1289 30948 1341
rect 31000 1289 31003 1341
rect 30945 1277 30957 1289
rect 30991 1277 31003 1289
rect 30945 1225 30948 1277
rect 31000 1225 31003 1277
rect 30945 1213 30957 1225
rect 30991 1213 31003 1225
rect 30945 1161 30948 1213
rect 31000 1161 31003 1213
rect 30945 1147 31003 1161
rect 31041 3133 31099 3147
rect 31041 3081 31044 3133
rect 31096 3081 31099 3133
rect 31041 3069 31053 3081
rect 31087 3069 31099 3081
rect 31041 3017 31044 3069
rect 31096 3017 31099 3069
rect 31041 3005 31053 3017
rect 31087 3005 31099 3017
rect 31041 2953 31044 3005
rect 31096 2953 31099 3005
rect 31041 2941 31053 2953
rect 31087 2941 31099 2953
rect 31041 2889 31044 2941
rect 31096 2889 31099 2941
rect 31041 2884 31099 2889
rect 31041 2877 31053 2884
rect 31087 2877 31099 2884
rect 31041 2825 31044 2877
rect 31096 2825 31099 2877
rect 31041 2813 31099 2825
rect 31041 2761 31044 2813
rect 31096 2761 31099 2813
rect 31041 2749 31099 2761
rect 31041 2697 31044 2749
rect 31096 2697 31099 2749
rect 31041 2685 31099 2697
rect 31041 2633 31044 2685
rect 31096 2633 31099 2685
rect 31041 2621 31099 2633
rect 31041 2569 31044 2621
rect 31096 2569 31099 2621
rect 31041 2562 31053 2569
rect 31087 2562 31099 2569
rect 31041 2557 31099 2562
rect 31041 2505 31044 2557
rect 31096 2505 31099 2557
rect 31041 2493 31053 2505
rect 31087 2493 31099 2505
rect 31041 2441 31044 2493
rect 31096 2441 31099 2493
rect 31041 2429 31053 2441
rect 31087 2429 31099 2441
rect 31041 2377 31044 2429
rect 31096 2377 31099 2429
rect 31041 2365 31053 2377
rect 31087 2365 31099 2377
rect 31041 2313 31044 2365
rect 31096 2313 31099 2365
rect 31041 2308 31099 2313
rect 31041 2301 31053 2308
rect 31087 2301 31099 2308
rect 31041 2249 31044 2301
rect 31096 2249 31099 2301
rect 31041 2237 31099 2249
rect 31041 2185 31044 2237
rect 31096 2185 31099 2237
rect 31041 2173 31099 2185
rect 31041 2121 31044 2173
rect 31096 2121 31099 2173
rect 31041 2109 31099 2121
rect 31041 2057 31044 2109
rect 31096 2057 31099 2109
rect 31041 2045 31099 2057
rect 31041 1993 31044 2045
rect 31096 1993 31099 2045
rect 31041 1986 31053 1993
rect 31087 1986 31099 1993
rect 31041 1981 31099 1986
rect 31041 1929 31044 1981
rect 31096 1929 31099 1981
rect 31041 1917 31053 1929
rect 31087 1917 31099 1929
rect 31041 1865 31044 1917
rect 31096 1865 31099 1917
rect 31041 1853 31053 1865
rect 31087 1853 31099 1865
rect 31041 1801 31044 1853
rect 31096 1801 31099 1853
rect 31041 1789 31053 1801
rect 31087 1789 31099 1801
rect 31041 1737 31044 1789
rect 31096 1737 31099 1789
rect 31041 1732 31099 1737
rect 31041 1725 31053 1732
rect 31087 1725 31099 1732
rect 31041 1673 31044 1725
rect 31096 1673 31099 1725
rect 31041 1661 31099 1673
rect 31041 1609 31044 1661
rect 31096 1609 31099 1661
rect 31041 1597 31099 1609
rect 31041 1545 31044 1597
rect 31096 1545 31099 1597
rect 31041 1533 31099 1545
rect 31041 1481 31044 1533
rect 31096 1481 31099 1533
rect 31041 1469 31099 1481
rect 31041 1417 31044 1469
rect 31096 1417 31099 1469
rect 31041 1410 31053 1417
rect 31087 1410 31099 1417
rect 31041 1405 31099 1410
rect 31041 1353 31044 1405
rect 31096 1353 31099 1405
rect 31041 1341 31053 1353
rect 31087 1341 31099 1353
rect 31041 1289 31044 1341
rect 31096 1289 31099 1341
rect 31041 1277 31053 1289
rect 31087 1277 31099 1289
rect 31041 1225 31044 1277
rect 31096 1225 31099 1277
rect 31041 1213 31053 1225
rect 31087 1213 31099 1225
rect 31041 1161 31044 1213
rect 31096 1161 31099 1213
rect 31041 1147 31099 1161
rect 31137 3133 31195 3147
rect 31137 3081 31140 3133
rect 31192 3081 31195 3133
rect 31137 3069 31149 3081
rect 31183 3069 31195 3081
rect 31137 3017 31140 3069
rect 31192 3017 31195 3069
rect 31137 3005 31149 3017
rect 31183 3005 31195 3017
rect 31137 2953 31140 3005
rect 31192 2953 31195 3005
rect 31137 2941 31149 2953
rect 31183 2941 31195 2953
rect 31137 2889 31140 2941
rect 31192 2889 31195 2941
rect 31137 2884 31195 2889
rect 31137 2877 31149 2884
rect 31183 2877 31195 2884
rect 31137 2825 31140 2877
rect 31192 2825 31195 2877
rect 31137 2813 31195 2825
rect 31137 2761 31140 2813
rect 31192 2761 31195 2813
rect 31137 2749 31195 2761
rect 31137 2697 31140 2749
rect 31192 2697 31195 2749
rect 31137 2685 31195 2697
rect 31137 2633 31140 2685
rect 31192 2633 31195 2685
rect 31137 2621 31195 2633
rect 31137 2569 31140 2621
rect 31192 2569 31195 2621
rect 31137 2562 31149 2569
rect 31183 2562 31195 2569
rect 31137 2557 31195 2562
rect 31137 2505 31140 2557
rect 31192 2505 31195 2557
rect 31137 2493 31149 2505
rect 31183 2493 31195 2505
rect 31137 2441 31140 2493
rect 31192 2441 31195 2493
rect 31137 2429 31149 2441
rect 31183 2429 31195 2441
rect 31137 2377 31140 2429
rect 31192 2377 31195 2429
rect 31137 2365 31149 2377
rect 31183 2365 31195 2377
rect 31137 2313 31140 2365
rect 31192 2313 31195 2365
rect 31137 2308 31195 2313
rect 31137 2301 31149 2308
rect 31183 2301 31195 2308
rect 31137 2249 31140 2301
rect 31192 2249 31195 2301
rect 31137 2237 31195 2249
rect 31137 2185 31140 2237
rect 31192 2185 31195 2237
rect 31137 2173 31195 2185
rect 31137 2121 31140 2173
rect 31192 2121 31195 2173
rect 31137 2109 31195 2121
rect 31137 2057 31140 2109
rect 31192 2057 31195 2109
rect 31137 2045 31195 2057
rect 31137 1993 31140 2045
rect 31192 1993 31195 2045
rect 31137 1986 31149 1993
rect 31183 1986 31195 1993
rect 31137 1981 31195 1986
rect 31137 1929 31140 1981
rect 31192 1929 31195 1981
rect 31137 1917 31149 1929
rect 31183 1917 31195 1929
rect 31137 1865 31140 1917
rect 31192 1865 31195 1917
rect 31137 1853 31149 1865
rect 31183 1853 31195 1865
rect 31137 1801 31140 1853
rect 31192 1801 31195 1853
rect 31137 1789 31149 1801
rect 31183 1789 31195 1801
rect 31137 1737 31140 1789
rect 31192 1737 31195 1789
rect 31137 1732 31195 1737
rect 31137 1725 31149 1732
rect 31183 1725 31195 1732
rect 31137 1673 31140 1725
rect 31192 1673 31195 1725
rect 31137 1661 31195 1673
rect 31137 1609 31140 1661
rect 31192 1609 31195 1661
rect 31137 1597 31195 1609
rect 31137 1545 31140 1597
rect 31192 1545 31195 1597
rect 31137 1533 31195 1545
rect 31137 1481 31140 1533
rect 31192 1481 31195 1533
rect 31137 1469 31195 1481
rect 31137 1417 31140 1469
rect 31192 1417 31195 1469
rect 31137 1410 31149 1417
rect 31183 1410 31195 1417
rect 31137 1405 31195 1410
rect 31137 1353 31140 1405
rect 31192 1353 31195 1405
rect 31137 1341 31149 1353
rect 31183 1341 31195 1353
rect 31137 1289 31140 1341
rect 31192 1289 31195 1341
rect 31137 1277 31149 1289
rect 31183 1277 31195 1289
rect 31137 1225 31140 1277
rect 31192 1225 31195 1277
rect 31137 1213 31149 1225
rect 31183 1213 31195 1225
rect 31137 1161 31140 1213
rect 31192 1161 31195 1213
rect 31137 1147 31195 1161
rect 31236 3133 31288 3147
rect 31236 3069 31245 3081
rect 31279 3069 31288 3081
rect 31236 3005 31245 3017
rect 31279 3005 31288 3017
rect 31236 2941 31245 2953
rect 31279 2941 31288 2953
rect 31236 2884 31288 2889
rect 31236 2877 31245 2884
rect 31279 2877 31288 2884
rect 31236 2813 31288 2825
rect 31236 2749 31288 2761
rect 31236 2685 31288 2697
rect 31236 2621 31288 2633
rect 31236 2562 31245 2569
rect 31279 2562 31288 2569
rect 31236 2557 31288 2562
rect 31236 2493 31245 2505
rect 31279 2493 31288 2505
rect 31236 2429 31245 2441
rect 31279 2429 31288 2441
rect 31236 2365 31245 2377
rect 31279 2365 31288 2377
rect 31236 2308 31288 2313
rect 31236 2301 31245 2308
rect 31279 2301 31288 2308
rect 31236 2237 31288 2249
rect 31236 2173 31288 2185
rect 31236 2109 31288 2121
rect 31236 2045 31288 2057
rect 31236 1986 31245 1993
rect 31279 1986 31288 1993
rect 31236 1981 31288 1986
rect 31236 1917 31245 1929
rect 31279 1917 31288 1929
rect 31236 1853 31245 1865
rect 31279 1853 31288 1865
rect 31236 1789 31245 1801
rect 31279 1789 31288 1801
rect 31236 1732 31288 1737
rect 31236 1725 31245 1732
rect 31279 1725 31288 1732
rect 31236 1661 31288 1673
rect 31236 1597 31288 1609
rect 31236 1533 31288 1545
rect 31236 1469 31288 1481
rect 31236 1410 31245 1417
rect 31279 1410 31288 1417
rect 31236 1405 31288 1410
rect 31236 1341 31245 1353
rect 31279 1341 31288 1353
rect 31236 1277 31245 1289
rect 31279 1277 31288 1289
rect 31236 1213 31245 1225
rect 31279 1213 31288 1225
rect 31236 1147 31288 1161
rect 31329 3133 31387 3147
rect 31329 3081 31332 3133
rect 31384 3081 31387 3133
rect 31329 3069 31341 3081
rect 31375 3069 31387 3081
rect 31329 3017 31332 3069
rect 31384 3017 31387 3069
rect 31329 3005 31341 3017
rect 31375 3005 31387 3017
rect 31329 2953 31332 3005
rect 31384 2953 31387 3005
rect 31329 2941 31341 2953
rect 31375 2941 31387 2953
rect 31329 2889 31332 2941
rect 31384 2889 31387 2941
rect 31329 2884 31387 2889
rect 31329 2877 31341 2884
rect 31375 2877 31387 2884
rect 31329 2825 31332 2877
rect 31384 2825 31387 2877
rect 31329 2813 31387 2825
rect 31329 2761 31332 2813
rect 31384 2761 31387 2813
rect 31329 2749 31387 2761
rect 31329 2697 31332 2749
rect 31384 2697 31387 2749
rect 31329 2685 31387 2697
rect 31329 2633 31332 2685
rect 31384 2633 31387 2685
rect 31329 2621 31387 2633
rect 31329 2569 31332 2621
rect 31384 2569 31387 2621
rect 31329 2562 31341 2569
rect 31375 2562 31387 2569
rect 31329 2557 31387 2562
rect 31329 2505 31332 2557
rect 31384 2505 31387 2557
rect 31329 2493 31341 2505
rect 31375 2493 31387 2505
rect 31329 2441 31332 2493
rect 31384 2441 31387 2493
rect 31329 2429 31341 2441
rect 31375 2429 31387 2441
rect 31329 2377 31332 2429
rect 31384 2377 31387 2429
rect 31329 2365 31341 2377
rect 31375 2365 31387 2377
rect 31329 2313 31332 2365
rect 31384 2313 31387 2365
rect 31329 2308 31387 2313
rect 31329 2301 31341 2308
rect 31375 2301 31387 2308
rect 31329 2249 31332 2301
rect 31384 2249 31387 2301
rect 31329 2237 31387 2249
rect 31329 2185 31332 2237
rect 31384 2185 31387 2237
rect 31329 2173 31387 2185
rect 31329 2121 31332 2173
rect 31384 2121 31387 2173
rect 31329 2109 31387 2121
rect 31329 2057 31332 2109
rect 31384 2057 31387 2109
rect 31329 2045 31387 2057
rect 31329 1993 31332 2045
rect 31384 1993 31387 2045
rect 31329 1986 31341 1993
rect 31375 1986 31387 1993
rect 31329 1981 31387 1986
rect 31329 1929 31332 1981
rect 31384 1929 31387 1981
rect 31329 1917 31341 1929
rect 31375 1917 31387 1929
rect 31329 1865 31332 1917
rect 31384 1865 31387 1917
rect 31329 1853 31341 1865
rect 31375 1853 31387 1865
rect 31329 1801 31332 1853
rect 31384 1801 31387 1853
rect 31329 1789 31341 1801
rect 31375 1789 31387 1801
rect 31329 1737 31332 1789
rect 31384 1737 31387 1789
rect 31329 1732 31387 1737
rect 31329 1725 31341 1732
rect 31375 1725 31387 1732
rect 31329 1673 31332 1725
rect 31384 1673 31387 1725
rect 31329 1661 31387 1673
rect 31329 1609 31332 1661
rect 31384 1609 31387 1661
rect 31329 1597 31387 1609
rect 31329 1545 31332 1597
rect 31384 1545 31387 1597
rect 31329 1533 31387 1545
rect 31329 1481 31332 1533
rect 31384 1481 31387 1533
rect 31329 1469 31387 1481
rect 31329 1417 31332 1469
rect 31384 1417 31387 1469
rect 31329 1410 31341 1417
rect 31375 1410 31387 1417
rect 31329 1405 31387 1410
rect 31329 1353 31332 1405
rect 31384 1353 31387 1405
rect 31329 1341 31341 1353
rect 31375 1341 31387 1353
rect 31329 1289 31332 1341
rect 31384 1289 31387 1341
rect 31329 1277 31341 1289
rect 31375 1277 31387 1289
rect 31329 1225 31332 1277
rect 31384 1225 31387 1277
rect 31329 1213 31341 1225
rect 31375 1213 31387 1225
rect 31329 1161 31332 1213
rect 31384 1161 31387 1213
rect 31329 1147 31387 1161
rect 31425 3133 31483 3147
rect 31425 3081 31428 3133
rect 31480 3081 31483 3133
rect 31425 3069 31437 3081
rect 31471 3069 31483 3081
rect 31425 3017 31428 3069
rect 31480 3017 31483 3069
rect 31425 3005 31437 3017
rect 31471 3005 31483 3017
rect 31425 2953 31428 3005
rect 31480 2953 31483 3005
rect 31425 2941 31437 2953
rect 31471 2941 31483 2953
rect 31425 2889 31428 2941
rect 31480 2889 31483 2941
rect 31425 2884 31483 2889
rect 31425 2877 31437 2884
rect 31471 2877 31483 2884
rect 31425 2825 31428 2877
rect 31480 2825 31483 2877
rect 31425 2813 31483 2825
rect 31425 2761 31428 2813
rect 31480 2761 31483 2813
rect 31425 2749 31483 2761
rect 31425 2697 31428 2749
rect 31480 2697 31483 2749
rect 31425 2685 31483 2697
rect 31425 2633 31428 2685
rect 31480 2633 31483 2685
rect 31425 2621 31483 2633
rect 31425 2569 31428 2621
rect 31480 2569 31483 2621
rect 31425 2562 31437 2569
rect 31471 2562 31483 2569
rect 31425 2557 31483 2562
rect 31425 2505 31428 2557
rect 31480 2505 31483 2557
rect 31425 2493 31437 2505
rect 31471 2493 31483 2505
rect 31425 2441 31428 2493
rect 31480 2441 31483 2493
rect 31425 2429 31437 2441
rect 31471 2429 31483 2441
rect 31425 2377 31428 2429
rect 31480 2377 31483 2429
rect 31425 2365 31437 2377
rect 31471 2365 31483 2377
rect 31425 2313 31428 2365
rect 31480 2313 31483 2365
rect 31425 2308 31483 2313
rect 31425 2301 31437 2308
rect 31471 2301 31483 2308
rect 31425 2249 31428 2301
rect 31480 2249 31483 2301
rect 31425 2237 31483 2249
rect 31425 2185 31428 2237
rect 31480 2185 31483 2237
rect 31425 2173 31483 2185
rect 31425 2121 31428 2173
rect 31480 2121 31483 2173
rect 31425 2109 31483 2121
rect 31425 2057 31428 2109
rect 31480 2057 31483 2109
rect 31425 2045 31483 2057
rect 31425 1993 31428 2045
rect 31480 1993 31483 2045
rect 31425 1986 31437 1993
rect 31471 1986 31483 1993
rect 31425 1981 31483 1986
rect 31425 1929 31428 1981
rect 31480 1929 31483 1981
rect 31425 1917 31437 1929
rect 31471 1917 31483 1929
rect 31425 1865 31428 1917
rect 31480 1865 31483 1917
rect 31425 1853 31437 1865
rect 31471 1853 31483 1865
rect 31425 1801 31428 1853
rect 31480 1801 31483 1853
rect 31425 1789 31437 1801
rect 31471 1789 31483 1801
rect 31425 1737 31428 1789
rect 31480 1737 31483 1789
rect 31425 1732 31483 1737
rect 31425 1725 31437 1732
rect 31471 1725 31483 1732
rect 31425 1673 31428 1725
rect 31480 1673 31483 1725
rect 31425 1661 31483 1673
rect 31425 1609 31428 1661
rect 31480 1609 31483 1661
rect 31425 1597 31483 1609
rect 31425 1545 31428 1597
rect 31480 1545 31483 1597
rect 31425 1533 31483 1545
rect 31425 1481 31428 1533
rect 31480 1481 31483 1533
rect 31425 1469 31483 1481
rect 31425 1417 31428 1469
rect 31480 1417 31483 1469
rect 31425 1410 31437 1417
rect 31471 1410 31483 1417
rect 31425 1405 31483 1410
rect 31425 1353 31428 1405
rect 31480 1353 31483 1405
rect 31425 1341 31437 1353
rect 31471 1341 31483 1353
rect 31425 1289 31428 1341
rect 31480 1289 31483 1341
rect 31425 1277 31437 1289
rect 31471 1277 31483 1289
rect 31425 1225 31428 1277
rect 31480 1225 31483 1277
rect 31425 1213 31437 1225
rect 31471 1213 31483 1225
rect 31425 1161 31428 1213
rect 31480 1161 31483 1213
rect 31425 1147 31483 1161
rect 31521 3133 31579 3147
rect 31521 3081 31524 3133
rect 31576 3081 31579 3133
rect 31521 3069 31533 3081
rect 31567 3069 31579 3081
rect 31521 3017 31524 3069
rect 31576 3017 31579 3069
rect 31521 3005 31533 3017
rect 31567 3005 31579 3017
rect 31521 2953 31524 3005
rect 31576 2953 31579 3005
rect 31521 2941 31533 2953
rect 31567 2941 31579 2953
rect 31521 2889 31524 2941
rect 31576 2889 31579 2941
rect 31521 2884 31579 2889
rect 31521 2877 31533 2884
rect 31567 2877 31579 2884
rect 31521 2825 31524 2877
rect 31576 2825 31579 2877
rect 31521 2813 31579 2825
rect 31521 2761 31524 2813
rect 31576 2761 31579 2813
rect 31521 2749 31579 2761
rect 31521 2697 31524 2749
rect 31576 2697 31579 2749
rect 31521 2685 31579 2697
rect 31521 2633 31524 2685
rect 31576 2633 31579 2685
rect 31521 2621 31579 2633
rect 31521 2569 31524 2621
rect 31576 2569 31579 2621
rect 31521 2562 31533 2569
rect 31567 2562 31579 2569
rect 31521 2557 31579 2562
rect 31521 2505 31524 2557
rect 31576 2505 31579 2557
rect 31521 2493 31533 2505
rect 31567 2493 31579 2505
rect 31521 2441 31524 2493
rect 31576 2441 31579 2493
rect 31521 2429 31533 2441
rect 31567 2429 31579 2441
rect 31521 2377 31524 2429
rect 31576 2377 31579 2429
rect 31521 2365 31533 2377
rect 31567 2365 31579 2377
rect 31521 2313 31524 2365
rect 31576 2313 31579 2365
rect 31521 2308 31579 2313
rect 31521 2301 31533 2308
rect 31567 2301 31579 2308
rect 31521 2249 31524 2301
rect 31576 2249 31579 2301
rect 31521 2237 31579 2249
rect 31521 2185 31524 2237
rect 31576 2185 31579 2237
rect 31521 2173 31579 2185
rect 31521 2121 31524 2173
rect 31576 2121 31579 2173
rect 31521 2109 31579 2121
rect 31521 2057 31524 2109
rect 31576 2057 31579 2109
rect 31521 2045 31579 2057
rect 31521 1993 31524 2045
rect 31576 1993 31579 2045
rect 31521 1986 31533 1993
rect 31567 1986 31579 1993
rect 31521 1981 31579 1986
rect 31521 1929 31524 1981
rect 31576 1929 31579 1981
rect 31521 1917 31533 1929
rect 31567 1917 31579 1929
rect 31521 1865 31524 1917
rect 31576 1865 31579 1917
rect 31521 1853 31533 1865
rect 31567 1853 31579 1865
rect 31521 1801 31524 1853
rect 31576 1801 31579 1853
rect 31521 1789 31533 1801
rect 31567 1789 31579 1801
rect 31521 1737 31524 1789
rect 31576 1737 31579 1789
rect 31521 1732 31579 1737
rect 31521 1725 31533 1732
rect 31567 1725 31579 1732
rect 31521 1673 31524 1725
rect 31576 1673 31579 1725
rect 31521 1661 31579 1673
rect 31521 1609 31524 1661
rect 31576 1609 31579 1661
rect 31521 1597 31579 1609
rect 31521 1545 31524 1597
rect 31576 1545 31579 1597
rect 31521 1533 31579 1545
rect 31521 1481 31524 1533
rect 31576 1481 31579 1533
rect 31521 1469 31579 1481
rect 31521 1417 31524 1469
rect 31576 1417 31579 1469
rect 31521 1410 31533 1417
rect 31567 1410 31579 1417
rect 31521 1405 31579 1410
rect 31521 1353 31524 1405
rect 31576 1353 31579 1405
rect 31521 1341 31533 1353
rect 31567 1341 31579 1353
rect 31521 1289 31524 1341
rect 31576 1289 31579 1341
rect 31521 1277 31533 1289
rect 31567 1277 31579 1289
rect 31521 1225 31524 1277
rect 31576 1225 31579 1277
rect 31521 1213 31533 1225
rect 31567 1213 31579 1225
rect 31521 1161 31524 1213
rect 31576 1161 31579 1213
rect 31521 1147 31579 1161
rect 31620 3133 31672 3147
rect 31620 3069 31629 3081
rect 31663 3069 31672 3081
rect 31620 3005 31629 3017
rect 31663 3005 31672 3017
rect 31620 2941 31629 2953
rect 31663 2941 31672 2953
rect 31620 2884 31672 2889
rect 31620 2877 31629 2884
rect 31663 2877 31672 2884
rect 31620 2813 31672 2825
rect 31620 2749 31672 2761
rect 31620 2685 31672 2697
rect 31620 2621 31672 2633
rect 31620 2562 31629 2569
rect 31663 2562 31672 2569
rect 31620 2557 31672 2562
rect 31620 2493 31629 2505
rect 31663 2493 31672 2505
rect 31620 2429 31629 2441
rect 31663 2429 31672 2441
rect 31620 2365 31629 2377
rect 31663 2365 31672 2377
rect 31620 2308 31672 2313
rect 31620 2301 31629 2308
rect 31663 2301 31672 2308
rect 31620 2237 31672 2249
rect 31620 2173 31672 2185
rect 31620 2109 31672 2121
rect 31620 2045 31672 2057
rect 31620 1986 31629 1993
rect 31663 1986 31672 1993
rect 31620 1981 31672 1986
rect 31620 1917 31629 1929
rect 31663 1917 31672 1929
rect 31620 1853 31629 1865
rect 31663 1853 31672 1865
rect 31620 1789 31629 1801
rect 31663 1789 31672 1801
rect 31620 1732 31672 1737
rect 31620 1725 31629 1732
rect 31663 1725 31672 1732
rect 31620 1661 31672 1673
rect 31620 1597 31672 1609
rect 31620 1533 31672 1545
rect 31620 1469 31672 1481
rect 31620 1410 31629 1417
rect 31663 1410 31672 1417
rect 31620 1405 31672 1410
rect 31620 1341 31629 1353
rect 31663 1341 31672 1353
rect 31620 1277 31629 1289
rect 31663 1277 31672 1289
rect 31620 1213 31629 1225
rect 31663 1213 31672 1225
rect 31620 1147 31672 1161
rect 31713 3133 31771 3147
rect 31713 3081 31716 3133
rect 31768 3081 31771 3133
rect 31713 3069 31725 3081
rect 31759 3069 31771 3081
rect 31713 3017 31716 3069
rect 31768 3017 31771 3069
rect 31713 3005 31725 3017
rect 31759 3005 31771 3017
rect 31713 2953 31716 3005
rect 31768 2953 31771 3005
rect 31713 2941 31725 2953
rect 31759 2941 31771 2953
rect 31713 2889 31716 2941
rect 31768 2889 31771 2941
rect 31713 2884 31771 2889
rect 31713 2877 31725 2884
rect 31759 2877 31771 2884
rect 31713 2825 31716 2877
rect 31768 2825 31771 2877
rect 31713 2813 31771 2825
rect 31713 2761 31716 2813
rect 31768 2761 31771 2813
rect 31713 2749 31771 2761
rect 31713 2697 31716 2749
rect 31768 2697 31771 2749
rect 31713 2685 31771 2697
rect 31713 2633 31716 2685
rect 31768 2633 31771 2685
rect 31713 2621 31771 2633
rect 31713 2569 31716 2621
rect 31768 2569 31771 2621
rect 31713 2562 31725 2569
rect 31759 2562 31771 2569
rect 31713 2557 31771 2562
rect 31713 2505 31716 2557
rect 31768 2505 31771 2557
rect 31713 2493 31725 2505
rect 31759 2493 31771 2505
rect 31713 2441 31716 2493
rect 31768 2441 31771 2493
rect 31713 2429 31725 2441
rect 31759 2429 31771 2441
rect 31713 2377 31716 2429
rect 31768 2377 31771 2429
rect 31713 2365 31725 2377
rect 31759 2365 31771 2377
rect 31713 2313 31716 2365
rect 31768 2313 31771 2365
rect 31713 2308 31771 2313
rect 31713 2301 31725 2308
rect 31759 2301 31771 2308
rect 31713 2249 31716 2301
rect 31768 2249 31771 2301
rect 31713 2237 31771 2249
rect 31713 2185 31716 2237
rect 31768 2185 31771 2237
rect 31713 2173 31771 2185
rect 31713 2121 31716 2173
rect 31768 2121 31771 2173
rect 31713 2109 31771 2121
rect 31713 2057 31716 2109
rect 31768 2057 31771 2109
rect 31713 2045 31771 2057
rect 31713 1993 31716 2045
rect 31768 1993 31771 2045
rect 31713 1986 31725 1993
rect 31759 1986 31771 1993
rect 31713 1981 31771 1986
rect 31713 1929 31716 1981
rect 31768 1929 31771 1981
rect 31713 1917 31725 1929
rect 31759 1917 31771 1929
rect 31713 1865 31716 1917
rect 31768 1865 31771 1917
rect 31713 1853 31725 1865
rect 31759 1853 31771 1865
rect 31713 1801 31716 1853
rect 31768 1801 31771 1853
rect 31713 1789 31725 1801
rect 31759 1789 31771 1801
rect 31713 1737 31716 1789
rect 31768 1737 31771 1789
rect 31713 1732 31771 1737
rect 31713 1725 31725 1732
rect 31759 1725 31771 1732
rect 31713 1673 31716 1725
rect 31768 1673 31771 1725
rect 31713 1661 31771 1673
rect 31713 1609 31716 1661
rect 31768 1609 31771 1661
rect 31713 1597 31771 1609
rect 31713 1545 31716 1597
rect 31768 1545 31771 1597
rect 31713 1533 31771 1545
rect 31713 1481 31716 1533
rect 31768 1481 31771 1533
rect 31713 1469 31771 1481
rect 31713 1417 31716 1469
rect 31768 1417 31771 1469
rect 31713 1410 31725 1417
rect 31759 1410 31771 1417
rect 31713 1405 31771 1410
rect 31713 1353 31716 1405
rect 31768 1353 31771 1405
rect 31713 1341 31725 1353
rect 31759 1341 31771 1353
rect 31713 1289 31716 1341
rect 31768 1289 31771 1341
rect 31713 1277 31725 1289
rect 31759 1277 31771 1289
rect 31713 1225 31716 1277
rect 31768 1225 31771 1277
rect 31713 1213 31725 1225
rect 31759 1213 31771 1225
rect 31713 1161 31716 1213
rect 31768 1161 31771 1213
rect 31713 1147 31771 1161
rect 31809 3133 31867 3147
rect 31809 3081 31812 3133
rect 31864 3081 31867 3133
rect 31809 3069 31821 3081
rect 31855 3069 31867 3081
rect 31809 3017 31812 3069
rect 31864 3017 31867 3069
rect 31809 3005 31821 3017
rect 31855 3005 31867 3017
rect 31809 2953 31812 3005
rect 31864 2953 31867 3005
rect 31809 2941 31821 2953
rect 31855 2941 31867 2953
rect 31809 2889 31812 2941
rect 31864 2889 31867 2941
rect 31809 2884 31867 2889
rect 31809 2877 31821 2884
rect 31855 2877 31867 2884
rect 31809 2825 31812 2877
rect 31864 2825 31867 2877
rect 31809 2813 31867 2825
rect 31809 2761 31812 2813
rect 31864 2761 31867 2813
rect 31809 2749 31867 2761
rect 31809 2697 31812 2749
rect 31864 2697 31867 2749
rect 31809 2685 31867 2697
rect 31809 2633 31812 2685
rect 31864 2633 31867 2685
rect 31809 2621 31867 2633
rect 31809 2569 31812 2621
rect 31864 2569 31867 2621
rect 31809 2562 31821 2569
rect 31855 2562 31867 2569
rect 31809 2557 31867 2562
rect 31809 2505 31812 2557
rect 31864 2505 31867 2557
rect 31809 2493 31821 2505
rect 31855 2493 31867 2505
rect 31809 2441 31812 2493
rect 31864 2441 31867 2493
rect 31809 2429 31821 2441
rect 31855 2429 31867 2441
rect 31809 2377 31812 2429
rect 31864 2377 31867 2429
rect 31809 2365 31821 2377
rect 31855 2365 31867 2377
rect 31809 2313 31812 2365
rect 31864 2313 31867 2365
rect 31809 2308 31867 2313
rect 31809 2301 31821 2308
rect 31855 2301 31867 2308
rect 31809 2249 31812 2301
rect 31864 2249 31867 2301
rect 31809 2237 31867 2249
rect 31809 2185 31812 2237
rect 31864 2185 31867 2237
rect 31809 2173 31867 2185
rect 31809 2121 31812 2173
rect 31864 2121 31867 2173
rect 31809 2109 31867 2121
rect 31809 2057 31812 2109
rect 31864 2057 31867 2109
rect 31809 2045 31867 2057
rect 31809 1993 31812 2045
rect 31864 1993 31867 2045
rect 31809 1986 31821 1993
rect 31855 1986 31867 1993
rect 31809 1981 31867 1986
rect 31809 1929 31812 1981
rect 31864 1929 31867 1981
rect 31809 1917 31821 1929
rect 31855 1917 31867 1929
rect 31809 1865 31812 1917
rect 31864 1865 31867 1917
rect 31809 1853 31821 1865
rect 31855 1853 31867 1865
rect 31809 1801 31812 1853
rect 31864 1801 31867 1853
rect 31809 1789 31821 1801
rect 31855 1789 31867 1801
rect 31809 1737 31812 1789
rect 31864 1737 31867 1789
rect 31809 1732 31867 1737
rect 31809 1725 31821 1732
rect 31855 1725 31867 1732
rect 31809 1673 31812 1725
rect 31864 1673 31867 1725
rect 31809 1661 31867 1673
rect 31809 1609 31812 1661
rect 31864 1609 31867 1661
rect 31809 1597 31867 1609
rect 31809 1545 31812 1597
rect 31864 1545 31867 1597
rect 31809 1533 31867 1545
rect 31809 1481 31812 1533
rect 31864 1481 31867 1533
rect 31809 1469 31867 1481
rect 31809 1417 31812 1469
rect 31864 1417 31867 1469
rect 31809 1410 31821 1417
rect 31855 1410 31867 1417
rect 31809 1405 31867 1410
rect 31809 1353 31812 1405
rect 31864 1353 31867 1405
rect 31809 1341 31821 1353
rect 31855 1341 31867 1353
rect 31809 1289 31812 1341
rect 31864 1289 31867 1341
rect 31809 1277 31821 1289
rect 31855 1277 31867 1289
rect 31809 1225 31812 1277
rect 31864 1225 31867 1277
rect 31809 1213 31821 1225
rect 31855 1213 31867 1225
rect 31809 1161 31812 1213
rect 31864 1161 31867 1213
rect 31809 1147 31867 1161
rect 31905 3133 31963 3147
rect 31905 3081 31908 3133
rect 31960 3081 31963 3133
rect 31905 3069 31917 3081
rect 31951 3069 31963 3081
rect 31905 3017 31908 3069
rect 31960 3017 31963 3069
rect 31905 3005 31917 3017
rect 31951 3005 31963 3017
rect 31905 2953 31908 3005
rect 31960 2953 31963 3005
rect 31905 2941 31917 2953
rect 31951 2941 31963 2953
rect 31905 2889 31908 2941
rect 31960 2889 31963 2941
rect 31905 2884 31963 2889
rect 31905 2877 31917 2884
rect 31951 2877 31963 2884
rect 31905 2825 31908 2877
rect 31960 2825 31963 2877
rect 31905 2813 31963 2825
rect 31905 2761 31908 2813
rect 31960 2761 31963 2813
rect 31905 2749 31963 2761
rect 31905 2697 31908 2749
rect 31960 2697 31963 2749
rect 31905 2685 31963 2697
rect 31905 2633 31908 2685
rect 31960 2633 31963 2685
rect 31905 2621 31963 2633
rect 31905 2569 31908 2621
rect 31960 2569 31963 2621
rect 31905 2562 31917 2569
rect 31951 2562 31963 2569
rect 31905 2557 31963 2562
rect 31905 2505 31908 2557
rect 31960 2505 31963 2557
rect 31905 2493 31917 2505
rect 31951 2493 31963 2505
rect 31905 2441 31908 2493
rect 31960 2441 31963 2493
rect 31905 2429 31917 2441
rect 31951 2429 31963 2441
rect 31905 2377 31908 2429
rect 31960 2377 31963 2429
rect 31905 2365 31917 2377
rect 31951 2365 31963 2377
rect 31905 2313 31908 2365
rect 31960 2313 31963 2365
rect 31905 2308 31963 2313
rect 31905 2301 31917 2308
rect 31951 2301 31963 2308
rect 31905 2249 31908 2301
rect 31960 2249 31963 2301
rect 31905 2237 31963 2249
rect 31905 2185 31908 2237
rect 31960 2185 31963 2237
rect 31905 2173 31963 2185
rect 31905 2121 31908 2173
rect 31960 2121 31963 2173
rect 31905 2109 31963 2121
rect 31905 2057 31908 2109
rect 31960 2057 31963 2109
rect 31905 2045 31963 2057
rect 31905 1993 31908 2045
rect 31960 1993 31963 2045
rect 31905 1986 31917 1993
rect 31951 1986 31963 1993
rect 31905 1981 31963 1986
rect 31905 1929 31908 1981
rect 31960 1929 31963 1981
rect 31905 1917 31917 1929
rect 31951 1917 31963 1929
rect 31905 1865 31908 1917
rect 31960 1865 31963 1917
rect 31905 1853 31917 1865
rect 31951 1853 31963 1865
rect 31905 1801 31908 1853
rect 31960 1801 31963 1853
rect 31905 1789 31917 1801
rect 31951 1789 31963 1801
rect 31905 1737 31908 1789
rect 31960 1737 31963 1789
rect 31905 1732 31963 1737
rect 31905 1725 31917 1732
rect 31951 1725 31963 1732
rect 31905 1673 31908 1725
rect 31960 1673 31963 1725
rect 31905 1661 31963 1673
rect 31905 1609 31908 1661
rect 31960 1609 31963 1661
rect 31905 1597 31963 1609
rect 31905 1545 31908 1597
rect 31960 1545 31963 1597
rect 31905 1533 31963 1545
rect 31905 1481 31908 1533
rect 31960 1481 31963 1533
rect 31905 1469 31963 1481
rect 31905 1417 31908 1469
rect 31960 1417 31963 1469
rect 31905 1410 31917 1417
rect 31951 1410 31963 1417
rect 31905 1405 31963 1410
rect 31905 1353 31908 1405
rect 31960 1353 31963 1405
rect 31905 1341 31917 1353
rect 31951 1341 31963 1353
rect 31905 1289 31908 1341
rect 31960 1289 31963 1341
rect 31905 1277 31917 1289
rect 31951 1277 31963 1289
rect 31905 1225 31908 1277
rect 31960 1225 31963 1277
rect 31905 1213 31917 1225
rect 31951 1213 31963 1225
rect 31905 1161 31908 1213
rect 31960 1161 31963 1213
rect 31905 1147 31963 1161
rect 32004 3133 32056 3147
rect 32004 3069 32013 3081
rect 32047 3069 32056 3081
rect 32004 3005 32013 3017
rect 32047 3005 32056 3017
rect 32004 2941 32013 2953
rect 32047 2941 32056 2953
rect 32004 2884 32056 2889
rect 32004 2877 32013 2884
rect 32047 2877 32056 2884
rect 32004 2813 32056 2825
rect 32004 2749 32056 2761
rect 32004 2685 32056 2697
rect 32004 2621 32056 2633
rect 32004 2562 32013 2569
rect 32047 2562 32056 2569
rect 32004 2557 32056 2562
rect 32004 2493 32013 2505
rect 32047 2493 32056 2505
rect 32004 2429 32013 2441
rect 32047 2429 32056 2441
rect 32004 2365 32013 2377
rect 32047 2365 32056 2377
rect 32004 2308 32056 2313
rect 32004 2301 32013 2308
rect 32047 2301 32056 2308
rect 32004 2237 32056 2249
rect 32004 2173 32056 2185
rect 32004 2109 32056 2121
rect 32004 2045 32056 2057
rect 32004 1986 32013 1993
rect 32047 1986 32056 1993
rect 32004 1981 32056 1986
rect 32004 1917 32013 1929
rect 32047 1917 32056 1929
rect 32004 1853 32013 1865
rect 32047 1853 32056 1865
rect 32004 1789 32013 1801
rect 32047 1789 32056 1801
rect 32004 1732 32056 1737
rect 32004 1725 32013 1732
rect 32047 1725 32056 1732
rect 32004 1661 32056 1673
rect 32004 1597 32056 1609
rect 32004 1533 32056 1545
rect 32004 1469 32056 1481
rect 32004 1410 32013 1417
rect 32047 1410 32056 1417
rect 32004 1405 32056 1410
rect 32004 1341 32013 1353
rect 32047 1341 32056 1353
rect 32004 1277 32013 1289
rect 32047 1277 32056 1289
rect 32004 1213 32013 1225
rect 32047 1213 32056 1225
rect 32004 1147 32056 1161
rect 32097 3133 32155 3147
rect 32097 3081 32100 3133
rect 32152 3081 32155 3133
rect 32097 3069 32109 3081
rect 32143 3069 32155 3081
rect 32097 3017 32100 3069
rect 32152 3017 32155 3069
rect 32097 3005 32109 3017
rect 32143 3005 32155 3017
rect 32097 2953 32100 3005
rect 32152 2953 32155 3005
rect 32097 2941 32109 2953
rect 32143 2941 32155 2953
rect 32097 2889 32100 2941
rect 32152 2889 32155 2941
rect 32097 2884 32155 2889
rect 32097 2877 32109 2884
rect 32143 2877 32155 2884
rect 32097 2825 32100 2877
rect 32152 2825 32155 2877
rect 32097 2813 32155 2825
rect 32097 2761 32100 2813
rect 32152 2761 32155 2813
rect 32097 2749 32155 2761
rect 32097 2697 32100 2749
rect 32152 2697 32155 2749
rect 32097 2685 32155 2697
rect 32097 2633 32100 2685
rect 32152 2633 32155 2685
rect 32097 2621 32155 2633
rect 32097 2569 32100 2621
rect 32152 2569 32155 2621
rect 32097 2562 32109 2569
rect 32143 2562 32155 2569
rect 32097 2557 32155 2562
rect 32097 2505 32100 2557
rect 32152 2505 32155 2557
rect 32097 2493 32109 2505
rect 32143 2493 32155 2505
rect 32097 2441 32100 2493
rect 32152 2441 32155 2493
rect 32097 2429 32109 2441
rect 32143 2429 32155 2441
rect 32097 2377 32100 2429
rect 32152 2377 32155 2429
rect 32097 2365 32109 2377
rect 32143 2365 32155 2377
rect 32097 2313 32100 2365
rect 32152 2313 32155 2365
rect 32097 2308 32155 2313
rect 32097 2301 32109 2308
rect 32143 2301 32155 2308
rect 32097 2249 32100 2301
rect 32152 2249 32155 2301
rect 32097 2237 32155 2249
rect 32097 2185 32100 2237
rect 32152 2185 32155 2237
rect 32097 2173 32155 2185
rect 32097 2121 32100 2173
rect 32152 2121 32155 2173
rect 32097 2109 32155 2121
rect 32097 2057 32100 2109
rect 32152 2057 32155 2109
rect 32097 2045 32155 2057
rect 32097 1993 32100 2045
rect 32152 1993 32155 2045
rect 32097 1986 32109 1993
rect 32143 1986 32155 1993
rect 32097 1981 32155 1986
rect 32097 1929 32100 1981
rect 32152 1929 32155 1981
rect 32097 1917 32109 1929
rect 32143 1917 32155 1929
rect 32097 1865 32100 1917
rect 32152 1865 32155 1917
rect 32097 1853 32109 1865
rect 32143 1853 32155 1865
rect 32097 1801 32100 1853
rect 32152 1801 32155 1853
rect 32097 1789 32109 1801
rect 32143 1789 32155 1801
rect 32097 1737 32100 1789
rect 32152 1737 32155 1789
rect 32097 1732 32155 1737
rect 32097 1725 32109 1732
rect 32143 1725 32155 1732
rect 32097 1673 32100 1725
rect 32152 1673 32155 1725
rect 32097 1661 32155 1673
rect 32097 1609 32100 1661
rect 32152 1609 32155 1661
rect 32097 1597 32155 1609
rect 32097 1545 32100 1597
rect 32152 1545 32155 1597
rect 32097 1533 32155 1545
rect 32097 1481 32100 1533
rect 32152 1481 32155 1533
rect 32097 1469 32155 1481
rect 32097 1417 32100 1469
rect 32152 1417 32155 1469
rect 32097 1410 32109 1417
rect 32143 1410 32155 1417
rect 32097 1405 32155 1410
rect 32097 1353 32100 1405
rect 32152 1353 32155 1405
rect 32097 1341 32109 1353
rect 32143 1341 32155 1353
rect 32097 1289 32100 1341
rect 32152 1289 32155 1341
rect 32097 1277 32109 1289
rect 32143 1277 32155 1289
rect 32097 1225 32100 1277
rect 32152 1225 32155 1277
rect 32097 1213 32109 1225
rect 32143 1213 32155 1225
rect 32097 1161 32100 1213
rect 32152 1161 32155 1213
rect 32097 1147 32155 1161
rect 32193 3133 32251 3147
rect 32193 3081 32196 3133
rect 32248 3081 32251 3133
rect 32193 3069 32205 3081
rect 32239 3069 32251 3081
rect 32193 3017 32196 3069
rect 32248 3017 32251 3069
rect 32193 3005 32205 3017
rect 32239 3005 32251 3017
rect 32193 2953 32196 3005
rect 32248 2953 32251 3005
rect 32193 2941 32205 2953
rect 32239 2941 32251 2953
rect 32193 2889 32196 2941
rect 32248 2889 32251 2941
rect 32193 2884 32251 2889
rect 32193 2877 32205 2884
rect 32239 2877 32251 2884
rect 32193 2825 32196 2877
rect 32248 2825 32251 2877
rect 32193 2813 32251 2825
rect 32193 2761 32196 2813
rect 32248 2761 32251 2813
rect 32193 2749 32251 2761
rect 32193 2697 32196 2749
rect 32248 2697 32251 2749
rect 32193 2685 32251 2697
rect 32193 2633 32196 2685
rect 32248 2633 32251 2685
rect 32193 2621 32251 2633
rect 32193 2569 32196 2621
rect 32248 2569 32251 2621
rect 32193 2562 32205 2569
rect 32239 2562 32251 2569
rect 32193 2557 32251 2562
rect 32193 2505 32196 2557
rect 32248 2505 32251 2557
rect 32193 2493 32205 2505
rect 32239 2493 32251 2505
rect 32193 2441 32196 2493
rect 32248 2441 32251 2493
rect 32193 2429 32205 2441
rect 32239 2429 32251 2441
rect 32193 2377 32196 2429
rect 32248 2377 32251 2429
rect 32193 2365 32205 2377
rect 32239 2365 32251 2377
rect 32193 2313 32196 2365
rect 32248 2313 32251 2365
rect 32193 2308 32251 2313
rect 32193 2301 32205 2308
rect 32239 2301 32251 2308
rect 32193 2249 32196 2301
rect 32248 2249 32251 2301
rect 32193 2237 32251 2249
rect 32193 2185 32196 2237
rect 32248 2185 32251 2237
rect 32193 2173 32251 2185
rect 32193 2121 32196 2173
rect 32248 2121 32251 2173
rect 32193 2109 32251 2121
rect 32193 2057 32196 2109
rect 32248 2057 32251 2109
rect 32193 2045 32251 2057
rect 32193 1993 32196 2045
rect 32248 1993 32251 2045
rect 32193 1986 32205 1993
rect 32239 1986 32251 1993
rect 32193 1981 32251 1986
rect 32193 1929 32196 1981
rect 32248 1929 32251 1981
rect 32193 1917 32205 1929
rect 32239 1917 32251 1929
rect 32193 1865 32196 1917
rect 32248 1865 32251 1917
rect 32193 1853 32205 1865
rect 32239 1853 32251 1865
rect 32193 1801 32196 1853
rect 32248 1801 32251 1853
rect 32193 1789 32205 1801
rect 32239 1789 32251 1801
rect 32193 1737 32196 1789
rect 32248 1737 32251 1789
rect 32193 1732 32251 1737
rect 32193 1725 32205 1732
rect 32239 1725 32251 1732
rect 32193 1673 32196 1725
rect 32248 1673 32251 1725
rect 32193 1661 32251 1673
rect 32193 1609 32196 1661
rect 32248 1609 32251 1661
rect 32193 1597 32251 1609
rect 32193 1545 32196 1597
rect 32248 1545 32251 1597
rect 32193 1533 32251 1545
rect 32193 1481 32196 1533
rect 32248 1481 32251 1533
rect 32193 1469 32251 1481
rect 32193 1417 32196 1469
rect 32248 1417 32251 1469
rect 32193 1410 32205 1417
rect 32239 1410 32251 1417
rect 32193 1405 32251 1410
rect 32193 1353 32196 1405
rect 32248 1353 32251 1405
rect 32193 1341 32205 1353
rect 32239 1341 32251 1353
rect 32193 1289 32196 1341
rect 32248 1289 32251 1341
rect 32193 1277 32205 1289
rect 32239 1277 32251 1289
rect 32193 1225 32196 1277
rect 32248 1225 32251 1277
rect 32193 1213 32205 1225
rect 32239 1213 32251 1225
rect 32193 1161 32196 1213
rect 32248 1161 32251 1213
rect 32193 1147 32251 1161
rect 32289 3133 32347 3147
rect 32289 3081 32292 3133
rect 32344 3081 32347 3133
rect 32289 3069 32301 3081
rect 32335 3069 32347 3081
rect 32289 3017 32292 3069
rect 32344 3017 32347 3069
rect 32289 3005 32301 3017
rect 32335 3005 32347 3017
rect 32289 2953 32292 3005
rect 32344 2953 32347 3005
rect 32289 2941 32301 2953
rect 32335 2941 32347 2953
rect 32289 2889 32292 2941
rect 32344 2889 32347 2941
rect 32289 2884 32347 2889
rect 32289 2877 32301 2884
rect 32335 2877 32347 2884
rect 32289 2825 32292 2877
rect 32344 2825 32347 2877
rect 32289 2813 32347 2825
rect 32289 2761 32292 2813
rect 32344 2761 32347 2813
rect 32289 2749 32347 2761
rect 32289 2697 32292 2749
rect 32344 2697 32347 2749
rect 32289 2685 32347 2697
rect 32289 2633 32292 2685
rect 32344 2633 32347 2685
rect 32289 2621 32347 2633
rect 32289 2569 32292 2621
rect 32344 2569 32347 2621
rect 32289 2562 32301 2569
rect 32335 2562 32347 2569
rect 32289 2557 32347 2562
rect 32289 2505 32292 2557
rect 32344 2505 32347 2557
rect 32289 2493 32301 2505
rect 32335 2493 32347 2505
rect 32289 2441 32292 2493
rect 32344 2441 32347 2493
rect 32289 2429 32301 2441
rect 32335 2429 32347 2441
rect 32289 2377 32292 2429
rect 32344 2377 32347 2429
rect 32289 2365 32301 2377
rect 32335 2365 32347 2377
rect 32289 2313 32292 2365
rect 32344 2313 32347 2365
rect 32289 2308 32347 2313
rect 32289 2301 32301 2308
rect 32335 2301 32347 2308
rect 32289 2249 32292 2301
rect 32344 2249 32347 2301
rect 32289 2237 32347 2249
rect 32289 2185 32292 2237
rect 32344 2185 32347 2237
rect 32289 2173 32347 2185
rect 32289 2121 32292 2173
rect 32344 2121 32347 2173
rect 32289 2109 32347 2121
rect 32289 2057 32292 2109
rect 32344 2057 32347 2109
rect 32289 2045 32347 2057
rect 32289 1993 32292 2045
rect 32344 1993 32347 2045
rect 32289 1986 32301 1993
rect 32335 1986 32347 1993
rect 32289 1981 32347 1986
rect 32289 1929 32292 1981
rect 32344 1929 32347 1981
rect 32289 1917 32301 1929
rect 32335 1917 32347 1929
rect 32289 1865 32292 1917
rect 32344 1865 32347 1917
rect 32289 1853 32301 1865
rect 32335 1853 32347 1865
rect 32289 1801 32292 1853
rect 32344 1801 32347 1853
rect 32289 1789 32301 1801
rect 32335 1789 32347 1801
rect 32289 1737 32292 1789
rect 32344 1737 32347 1789
rect 32289 1732 32347 1737
rect 32289 1725 32301 1732
rect 32335 1725 32347 1732
rect 32289 1673 32292 1725
rect 32344 1673 32347 1725
rect 32289 1661 32347 1673
rect 32289 1609 32292 1661
rect 32344 1609 32347 1661
rect 32289 1597 32347 1609
rect 32289 1545 32292 1597
rect 32344 1545 32347 1597
rect 32289 1533 32347 1545
rect 32289 1481 32292 1533
rect 32344 1481 32347 1533
rect 32289 1469 32347 1481
rect 32289 1417 32292 1469
rect 32344 1417 32347 1469
rect 32289 1410 32301 1417
rect 32335 1410 32347 1417
rect 32289 1405 32347 1410
rect 32289 1353 32292 1405
rect 32344 1353 32347 1405
rect 32289 1341 32301 1353
rect 32335 1341 32347 1353
rect 32289 1289 32292 1341
rect 32344 1289 32347 1341
rect 32289 1277 32301 1289
rect 32335 1277 32347 1289
rect 32289 1225 32292 1277
rect 32344 1225 32347 1277
rect 32289 1213 32301 1225
rect 32335 1213 32347 1225
rect 32289 1161 32292 1213
rect 32344 1161 32347 1213
rect 32289 1147 32347 1161
rect 32388 3133 32440 3147
rect 32388 3069 32397 3081
rect 32431 3069 32440 3081
rect 32388 3005 32397 3017
rect 32431 3005 32440 3017
rect 32388 2941 32397 2953
rect 32431 2941 32440 2953
rect 32388 2884 32440 2889
rect 32388 2877 32397 2884
rect 32431 2877 32440 2884
rect 32388 2813 32440 2825
rect 32388 2749 32440 2761
rect 32388 2685 32440 2697
rect 32388 2621 32440 2633
rect 32388 2562 32397 2569
rect 32431 2562 32440 2569
rect 32388 2557 32440 2562
rect 32388 2493 32397 2505
rect 32431 2493 32440 2505
rect 32388 2429 32397 2441
rect 32431 2429 32440 2441
rect 32388 2365 32397 2377
rect 32431 2365 32440 2377
rect 32388 2308 32440 2313
rect 32388 2301 32397 2308
rect 32431 2301 32440 2308
rect 32388 2237 32440 2249
rect 32388 2173 32440 2185
rect 32388 2109 32440 2121
rect 32388 2045 32440 2057
rect 32388 1986 32397 1993
rect 32431 1986 32440 1993
rect 32388 1981 32440 1986
rect 32388 1917 32397 1929
rect 32431 1917 32440 1929
rect 32388 1853 32397 1865
rect 32431 1853 32440 1865
rect 32388 1789 32397 1801
rect 32431 1789 32440 1801
rect 32388 1732 32440 1737
rect 32388 1725 32397 1732
rect 32431 1725 32440 1732
rect 32388 1661 32440 1673
rect 32388 1597 32440 1609
rect 32388 1533 32440 1545
rect 32388 1469 32440 1481
rect 32388 1410 32397 1417
rect 32431 1410 32440 1417
rect 32388 1405 32440 1410
rect 32388 1341 32397 1353
rect 32431 1341 32440 1353
rect 32388 1277 32397 1289
rect 32431 1277 32440 1289
rect 32388 1213 32397 1225
rect 32431 1213 32440 1225
rect 32388 1147 32440 1161
rect 32481 3133 32539 3147
rect 32481 3081 32484 3133
rect 32536 3081 32539 3133
rect 32481 3069 32493 3081
rect 32527 3069 32539 3081
rect 32481 3017 32484 3069
rect 32536 3017 32539 3069
rect 32481 3005 32493 3017
rect 32527 3005 32539 3017
rect 32481 2953 32484 3005
rect 32536 2953 32539 3005
rect 32481 2941 32493 2953
rect 32527 2941 32539 2953
rect 32481 2889 32484 2941
rect 32536 2889 32539 2941
rect 32481 2884 32539 2889
rect 32481 2877 32493 2884
rect 32527 2877 32539 2884
rect 32481 2825 32484 2877
rect 32536 2825 32539 2877
rect 32481 2813 32539 2825
rect 32481 2761 32484 2813
rect 32536 2761 32539 2813
rect 32481 2749 32539 2761
rect 32481 2697 32484 2749
rect 32536 2697 32539 2749
rect 32481 2685 32539 2697
rect 32481 2633 32484 2685
rect 32536 2633 32539 2685
rect 32481 2621 32539 2633
rect 32481 2569 32484 2621
rect 32536 2569 32539 2621
rect 32481 2562 32493 2569
rect 32527 2562 32539 2569
rect 32481 2557 32539 2562
rect 32481 2505 32484 2557
rect 32536 2505 32539 2557
rect 32481 2493 32493 2505
rect 32527 2493 32539 2505
rect 32481 2441 32484 2493
rect 32536 2441 32539 2493
rect 32481 2429 32493 2441
rect 32527 2429 32539 2441
rect 32481 2377 32484 2429
rect 32536 2377 32539 2429
rect 32481 2365 32493 2377
rect 32527 2365 32539 2377
rect 32481 2313 32484 2365
rect 32536 2313 32539 2365
rect 32481 2308 32539 2313
rect 32481 2301 32493 2308
rect 32527 2301 32539 2308
rect 32481 2249 32484 2301
rect 32536 2249 32539 2301
rect 32481 2237 32539 2249
rect 32481 2185 32484 2237
rect 32536 2185 32539 2237
rect 32481 2173 32539 2185
rect 32481 2121 32484 2173
rect 32536 2121 32539 2173
rect 32481 2109 32539 2121
rect 32481 2057 32484 2109
rect 32536 2057 32539 2109
rect 32481 2045 32539 2057
rect 32481 1993 32484 2045
rect 32536 1993 32539 2045
rect 32481 1986 32493 1993
rect 32527 1986 32539 1993
rect 32481 1981 32539 1986
rect 32481 1929 32484 1981
rect 32536 1929 32539 1981
rect 32481 1917 32493 1929
rect 32527 1917 32539 1929
rect 32481 1865 32484 1917
rect 32536 1865 32539 1917
rect 32481 1853 32493 1865
rect 32527 1853 32539 1865
rect 32481 1801 32484 1853
rect 32536 1801 32539 1853
rect 32481 1789 32493 1801
rect 32527 1789 32539 1801
rect 32481 1737 32484 1789
rect 32536 1737 32539 1789
rect 32481 1732 32539 1737
rect 32481 1725 32493 1732
rect 32527 1725 32539 1732
rect 32481 1673 32484 1725
rect 32536 1673 32539 1725
rect 32481 1661 32539 1673
rect 32481 1609 32484 1661
rect 32536 1609 32539 1661
rect 32481 1597 32539 1609
rect 32481 1545 32484 1597
rect 32536 1545 32539 1597
rect 32481 1533 32539 1545
rect 32481 1481 32484 1533
rect 32536 1481 32539 1533
rect 32481 1469 32539 1481
rect 32481 1417 32484 1469
rect 32536 1417 32539 1469
rect 32481 1410 32493 1417
rect 32527 1410 32539 1417
rect 32481 1405 32539 1410
rect 32481 1353 32484 1405
rect 32536 1353 32539 1405
rect 32481 1341 32493 1353
rect 32527 1341 32539 1353
rect 32481 1289 32484 1341
rect 32536 1289 32539 1341
rect 32481 1277 32493 1289
rect 32527 1277 32539 1289
rect 32481 1225 32484 1277
rect 32536 1225 32539 1277
rect 32481 1213 32493 1225
rect 32527 1213 32539 1225
rect 32481 1161 32484 1213
rect 32536 1161 32539 1213
rect 32481 1147 32539 1161
rect 32577 3133 32635 3147
rect 32577 3081 32580 3133
rect 32632 3081 32635 3133
rect 32577 3069 32589 3081
rect 32623 3069 32635 3081
rect 32577 3017 32580 3069
rect 32632 3017 32635 3069
rect 32577 3005 32589 3017
rect 32623 3005 32635 3017
rect 32577 2953 32580 3005
rect 32632 2953 32635 3005
rect 32577 2941 32589 2953
rect 32623 2941 32635 2953
rect 32577 2889 32580 2941
rect 32632 2889 32635 2941
rect 32577 2884 32635 2889
rect 32577 2877 32589 2884
rect 32623 2877 32635 2884
rect 32577 2825 32580 2877
rect 32632 2825 32635 2877
rect 32577 2813 32635 2825
rect 32577 2761 32580 2813
rect 32632 2761 32635 2813
rect 32577 2749 32635 2761
rect 32577 2697 32580 2749
rect 32632 2697 32635 2749
rect 32577 2685 32635 2697
rect 32577 2633 32580 2685
rect 32632 2633 32635 2685
rect 32577 2621 32635 2633
rect 32577 2569 32580 2621
rect 32632 2569 32635 2621
rect 32577 2562 32589 2569
rect 32623 2562 32635 2569
rect 32577 2557 32635 2562
rect 32577 2505 32580 2557
rect 32632 2505 32635 2557
rect 32577 2493 32589 2505
rect 32623 2493 32635 2505
rect 32577 2441 32580 2493
rect 32632 2441 32635 2493
rect 32577 2429 32589 2441
rect 32623 2429 32635 2441
rect 32577 2377 32580 2429
rect 32632 2377 32635 2429
rect 32577 2365 32589 2377
rect 32623 2365 32635 2377
rect 32577 2313 32580 2365
rect 32632 2313 32635 2365
rect 32577 2308 32635 2313
rect 32577 2301 32589 2308
rect 32623 2301 32635 2308
rect 32577 2249 32580 2301
rect 32632 2249 32635 2301
rect 32577 2237 32635 2249
rect 32577 2185 32580 2237
rect 32632 2185 32635 2237
rect 32577 2173 32635 2185
rect 32577 2121 32580 2173
rect 32632 2121 32635 2173
rect 32577 2109 32635 2121
rect 32577 2057 32580 2109
rect 32632 2057 32635 2109
rect 32577 2045 32635 2057
rect 32577 1993 32580 2045
rect 32632 1993 32635 2045
rect 32577 1986 32589 1993
rect 32623 1986 32635 1993
rect 32577 1981 32635 1986
rect 32577 1929 32580 1981
rect 32632 1929 32635 1981
rect 32577 1917 32589 1929
rect 32623 1917 32635 1929
rect 32577 1865 32580 1917
rect 32632 1865 32635 1917
rect 32577 1853 32589 1865
rect 32623 1853 32635 1865
rect 32577 1801 32580 1853
rect 32632 1801 32635 1853
rect 32577 1789 32589 1801
rect 32623 1789 32635 1801
rect 32577 1737 32580 1789
rect 32632 1737 32635 1789
rect 32577 1732 32635 1737
rect 32577 1725 32589 1732
rect 32623 1725 32635 1732
rect 32577 1673 32580 1725
rect 32632 1673 32635 1725
rect 32577 1661 32635 1673
rect 32577 1609 32580 1661
rect 32632 1609 32635 1661
rect 32577 1597 32635 1609
rect 32577 1545 32580 1597
rect 32632 1545 32635 1597
rect 32577 1533 32635 1545
rect 32577 1481 32580 1533
rect 32632 1481 32635 1533
rect 32577 1469 32635 1481
rect 32577 1417 32580 1469
rect 32632 1417 32635 1469
rect 32577 1410 32589 1417
rect 32623 1410 32635 1417
rect 32577 1405 32635 1410
rect 32577 1353 32580 1405
rect 32632 1353 32635 1405
rect 32577 1341 32589 1353
rect 32623 1341 32635 1353
rect 32577 1289 32580 1341
rect 32632 1289 32635 1341
rect 32577 1277 32589 1289
rect 32623 1277 32635 1289
rect 32577 1225 32580 1277
rect 32632 1225 32635 1277
rect 32577 1213 32589 1225
rect 32623 1213 32635 1225
rect 32577 1161 32580 1213
rect 32632 1161 32635 1213
rect 32577 1147 32635 1161
rect 32673 3133 32731 3147
rect 32673 3081 32676 3133
rect 32728 3081 32731 3133
rect 32673 3069 32685 3081
rect 32719 3069 32731 3081
rect 32673 3017 32676 3069
rect 32728 3017 32731 3069
rect 32673 3005 32685 3017
rect 32719 3005 32731 3017
rect 32673 2953 32676 3005
rect 32728 2953 32731 3005
rect 32673 2941 32685 2953
rect 32719 2941 32731 2953
rect 32673 2889 32676 2941
rect 32728 2889 32731 2941
rect 32673 2884 32731 2889
rect 32673 2877 32685 2884
rect 32719 2877 32731 2884
rect 32673 2825 32676 2877
rect 32728 2825 32731 2877
rect 32673 2813 32731 2825
rect 32673 2761 32676 2813
rect 32728 2761 32731 2813
rect 32673 2749 32731 2761
rect 32673 2697 32676 2749
rect 32728 2697 32731 2749
rect 32673 2685 32731 2697
rect 32673 2633 32676 2685
rect 32728 2633 32731 2685
rect 32673 2621 32731 2633
rect 32673 2569 32676 2621
rect 32728 2569 32731 2621
rect 32673 2562 32685 2569
rect 32719 2562 32731 2569
rect 32673 2557 32731 2562
rect 32673 2505 32676 2557
rect 32728 2505 32731 2557
rect 32673 2493 32685 2505
rect 32719 2493 32731 2505
rect 32673 2441 32676 2493
rect 32728 2441 32731 2493
rect 32673 2429 32685 2441
rect 32719 2429 32731 2441
rect 32673 2377 32676 2429
rect 32728 2377 32731 2429
rect 32673 2365 32685 2377
rect 32719 2365 32731 2377
rect 32673 2313 32676 2365
rect 32728 2313 32731 2365
rect 32673 2308 32731 2313
rect 32673 2301 32685 2308
rect 32719 2301 32731 2308
rect 32673 2249 32676 2301
rect 32728 2249 32731 2301
rect 32673 2237 32731 2249
rect 32673 2185 32676 2237
rect 32728 2185 32731 2237
rect 32673 2173 32731 2185
rect 32673 2121 32676 2173
rect 32728 2121 32731 2173
rect 32673 2109 32731 2121
rect 32673 2057 32676 2109
rect 32728 2057 32731 2109
rect 32673 2045 32731 2057
rect 32673 1993 32676 2045
rect 32728 1993 32731 2045
rect 32673 1986 32685 1993
rect 32719 1986 32731 1993
rect 32673 1981 32731 1986
rect 32673 1929 32676 1981
rect 32728 1929 32731 1981
rect 32673 1917 32685 1929
rect 32719 1917 32731 1929
rect 32673 1865 32676 1917
rect 32728 1865 32731 1917
rect 32673 1853 32685 1865
rect 32719 1853 32731 1865
rect 32673 1801 32676 1853
rect 32728 1801 32731 1853
rect 32673 1789 32685 1801
rect 32719 1789 32731 1801
rect 32673 1737 32676 1789
rect 32728 1737 32731 1789
rect 32673 1732 32731 1737
rect 32673 1725 32685 1732
rect 32719 1725 32731 1732
rect 32673 1673 32676 1725
rect 32728 1673 32731 1725
rect 32673 1661 32731 1673
rect 32673 1609 32676 1661
rect 32728 1609 32731 1661
rect 32673 1597 32731 1609
rect 32673 1545 32676 1597
rect 32728 1545 32731 1597
rect 32673 1533 32731 1545
rect 32673 1481 32676 1533
rect 32728 1481 32731 1533
rect 32673 1469 32731 1481
rect 32673 1417 32676 1469
rect 32728 1417 32731 1469
rect 32673 1410 32685 1417
rect 32719 1410 32731 1417
rect 32673 1405 32731 1410
rect 32673 1353 32676 1405
rect 32728 1353 32731 1405
rect 32673 1341 32685 1353
rect 32719 1341 32731 1353
rect 32673 1289 32676 1341
rect 32728 1289 32731 1341
rect 32673 1277 32685 1289
rect 32719 1277 32731 1289
rect 32673 1225 32676 1277
rect 32728 1225 32731 1277
rect 32673 1213 32685 1225
rect 32719 1213 32731 1225
rect 32673 1161 32676 1213
rect 32728 1161 32731 1213
rect 32673 1147 32731 1161
rect 32772 3133 32824 3147
rect 32772 3069 32781 3081
rect 32815 3069 32824 3081
rect 32772 3005 32781 3017
rect 32815 3005 32824 3017
rect 32772 2941 32781 2953
rect 32815 2941 32824 2953
rect 32772 2884 32824 2889
rect 32772 2877 32781 2884
rect 32815 2877 32824 2884
rect 32772 2813 32824 2825
rect 32772 2749 32824 2761
rect 32772 2685 32824 2697
rect 32772 2621 32824 2633
rect 32772 2562 32781 2569
rect 32815 2562 32824 2569
rect 32772 2557 32824 2562
rect 32772 2493 32781 2505
rect 32815 2493 32824 2505
rect 32772 2429 32781 2441
rect 32815 2429 32824 2441
rect 32772 2365 32781 2377
rect 32815 2365 32824 2377
rect 32772 2308 32824 2313
rect 32772 2301 32781 2308
rect 32815 2301 32824 2308
rect 32772 2237 32824 2249
rect 32772 2173 32824 2185
rect 32772 2109 32824 2121
rect 32772 2045 32824 2057
rect 32772 1986 32781 1993
rect 32815 1986 32824 1993
rect 32772 1981 32824 1986
rect 32772 1917 32781 1929
rect 32815 1917 32824 1929
rect 32772 1853 32781 1865
rect 32815 1853 32824 1865
rect 32772 1789 32781 1801
rect 32815 1789 32824 1801
rect 32772 1732 32824 1737
rect 32772 1725 32781 1732
rect 32815 1725 32824 1732
rect 32772 1661 32824 1673
rect 32772 1597 32824 1609
rect 32772 1533 32824 1545
rect 32772 1469 32824 1481
rect 32772 1410 32781 1417
rect 32815 1410 32824 1417
rect 32772 1405 32824 1410
rect 32772 1341 32781 1353
rect 32815 1341 32824 1353
rect 32772 1277 32781 1289
rect 32815 1277 32824 1289
rect 32772 1213 32781 1225
rect 32815 1213 32824 1225
rect 32772 1147 32824 1161
rect 32865 3133 32923 3147
rect 32865 3081 32868 3133
rect 32920 3081 32923 3133
rect 32865 3069 32877 3081
rect 32911 3069 32923 3081
rect 32865 3017 32868 3069
rect 32920 3017 32923 3069
rect 32865 3005 32877 3017
rect 32911 3005 32923 3017
rect 32865 2953 32868 3005
rect 32920 2953 32923 3005
rect 32865 2941 32877 2953
rect 32911 2941 32923 2953
rect 32865 2889 32868 2941
rect 32920 2889 32923 2941
rect 32865 2884 32923 2889
rect 32865 2877 32877 2884
rect 32911 2877 32923 2884
rect 32865 2825 32868 2877
rect 32920 2825 32923 2877
rect 32865 2813 32923 2825
rect 32865 2761 32868 2813
rect 32920 2761 32923 2813
rect 32865 2749 32923 2761
rect 32865 2697 32868 2749
rect 32920 2697 32923 2749
rect 32865 2685 32923 2697
rect 32865 2633 32868 2685
rect 32920 2633 32923 2685
rect 32865 2621 32923 2633
rect 32865 2569 32868 2621
rect 32920 2569 32923 2621
rect 32865 2562 32877 2569
rect 32911 2562 32923 2569
rect 32865 2557 32923 2562
rect 32865 2505 32868 2557
rect 32920 2505 32923 2557
rect 32865 2493 32877 2505
rect 32911 2493 32923 2505
rect 32865 2441 32868 2493
rect 32920 2441 32923 2493
rect 32865 2429 32877 2441
rect 32911 2429 32923 2441
rect 32865 2377 32868 2429
rect 32920 2377 32923 2429
rect 32865 2365 32877 2377
rect 32911 2365 32923 2377
rect 32865 2313 32868 2365
rect 32920 2313 32923 2365
rect 32865 2308 32923 2313
rect 32865 2301 32877 2308
rect 32911 2301 32923 2308
rect 32865 2249 32868 2301
rect 32920 2249 32923 2301
rect 32865 2237 32923 2249
rect 32865 2185 32868 2237
rect 32920 2185 32923 2237
rect 32865 2173 32923 2185
rect 32865 2121 32868 2173
rect 32920 2121 32923 2173
rect 32865 2109 32923 2121
rect 32865 2057 32868 2109
rect 32920 2057 32923 2109
rect 32865 2045 32923 2057
rect 32865 1993 32868 2045
rect 32920 1993 32923 2045
rect 32865 1986 32877 1993
rect 32911 1986 32923 1993
rect 32865 1981 32923 1986
rect 32865 1929 32868 1981
rect 32920 1929 32923 1981
rect 32865 1917 32877 1929
rect 32911 1917 32923 1929
rect 32865 1865 32868 1917
rect 32920 1865 32923 1917
rect 32865 1853 32877 1865
rect 32911 1853 32923 1865
rect 32865 1801 32868 1853
rect 32920 1801 32923 1853
rect 32865 1789 32877 1801
rect 32911 1789 32923 1801
rect 32865 1737 32868 1789
rect 32920 1737 32923 1789
rect 32865 1732 32923 1737
rect 32865 1725 32877 1732
rect 32911 1725 32923 1732
rect 32865 1673 32868 1725
rect 32920 1673 32923 1725
rect 32865 1661 32923 1673
rect 32865 1609 32868 1661
rect 32920 1609 32923 1661
rect 32865 1597 32923 1609
rect 32865 1545 32868 1597
rect 32920 1545 32923 1597
rect 32865 1533 32923 1545
rect 32865 1481 32868 1533
rect 32920 1481 32923 1533
rect 32865 1469 32923 1481
rect 32865 1417 32868 1469
rect 32920 1417 32923 1469
rect 32865 1410 32877 1417
rect 32911 1410 32923 1417
rect 32865 1405 32923 1410
rect 32865 1353 32868 1405
rect 32920 1353 32923 1405
rect 32865 1341 32877 1353
rect 32911 1341 32923 1353
rect 32865 1289 32868 1341
rect 32920 1289 32923 1341
rect 32865 1277 32877 1289
rect 32911 1277 32923 1289
rect 32865 1225 32868 1277
rect 32920 1225 32923 1277
rect 32865 1213 32877 1225
rect 32911 1213 32923 1225
rect 32865 1161 32868 1213
rect 32920 1161 32923 1213
rect 32865 1147 32923 1161
rect 32961 3133 33019 3147
rect 32961 3081 32964 3133
rect 33016 3081 33019 3133
rect 32961 3069 32973 3081
rect 33007 3069 33019 3081
rect 32961 3017 32964 3069
rect 33016 3017 33019 3069
rect 32961 3005 32973 3017
rect 33007 3005 33019 3017
rect 32961 2953 32964 3005
rect 33016 2953 33019 3005
rect 32961 2941 32973 2953
rect 33007 2941 33019 2953
rect 32961 2889 32964 2941
rect 33016 2889 33019 2941
rect 32961 2884 33019 2889
rect 32961 2877 32973 2884
rect 33007 2877 33019 2884
rect 32961 2825 32964 2877
rect 33016 2825 33019 2877
rect 32961 2813 33019 2825
rect 32961 2761 32964 2813
rect 33016 2761 33019 2813
rect 32961 2749 33019 2761
rect 32961 2697 32964 2749
rect 33016 2697 33019 2749
rect 32961 2685 33019 2697
rect 32961 2633 32964 2685
rect 33016 2633 33019 2685
rect 32961 2621 33019 2633
rect 32961 2569 32964 2621
rect 33016 2569 33019 2621
rect 32961 2562 32973 2569
rect 33007 2562 33019 2569
rect 32961 2557 33019 2562
rect 32961 2505 32964 2557
rect 33016 2505 33019 2557
rect 32961 2493 32973 2505
rect 33007 2493 33019 2505
rect 32961 2441 32964 2493
rect 33016 2441 33019 2493
rect 32961 2429 32973 2441
rect 33007 2429 33019 2441
rect 32961 2377 32964 2429
rect 33016 2377 33019 2429
rect 32961 2365 32973 2377
rect 33007 2365 33019 2377
rect 32961 2313 32964 2365
rect 33016 2313 33019 2365
rect 32961 2308 33019 2313
rect 32961 2301 32973 2308
rect 33007 2301 33019 2308
rect 32961 2249 32964 2301
rect 33016 2249 33019 2301
rect 32961 2237 33019 2249
rect 32961 2185 32964 2237
rect 33016 2185 33019 2237
rect 32961 2173 33019 2185
rect 32961 2121 32964 2173
rect 33016 2121 33019 2173
rect 32961 2109 33019 2121
rect 32961 2057 32964 2109
rect 33016 2057 33019 2109
rect 32961 2045 33019 2057
rect 32961 1993 32964 2045
rect 33016 1993 33019 2045
rect 32961 1986 32973 1993
rect 33007 1986 33019 1993
rect 32961 1981 33019 1986
rect 32961 1929 32964 1981
rect 33016 1929 33019 1981
rect 32961 1917 32973 1929
rect 33007 1917 33019 1929
rect 32961 1865 32964 1917
rect 33016 1865 33019 1917
rect 32961 1853 32973 1865
rect 33007 1853 33019 1865
rect 32961 1801 32964 1853
rect 33016 1801 33019 1853
rect 32961 1789 32973 1801
rect 33007 1789 33019 1801
rect 32961 1737 32964 1789
rect 33016 1737 33019 1789
rect 32961 1732 33019 1737
rect 32961 1725 32973 1732
rect 33007 1725 33019 1732
rect 32961 1673 32964 1725
rect 33016 1673 33019 1725
rect 32961 1661 33019 1673
rect 32961 1609 32964 1661
rect 33016 1609 33019 1661
rect 32961 1597 33019 1609
rect 32961 1545 32964 1597
rect 33016 1545 33019 1597
rect 32961 1533 33019 1545
rect 32961 1481 32964 1533
rect 33016 1481 33019 1533
rect 32961 1469 33019 1481
rect 32961 1417 32964 1469
rect 33016 1417 33019 1469
rect 32961 1410 32973 1417
rect 33007 1410 33019 1417
rect 32961 1405 33019 1410
rect 32961 1353 32964 1405
rect 33016 1353 33019 1405
rect 32961 1341 32973 1353
rect 33007 1341 33019 1353
rect 32961 1289 32964 1341
rect 33016 1289 33019 1341
rect 32961 1277 32973 1289
rect 33007 1277 33019 1289
rect 32961 1225 32964 1277
rect 33016 1225 33019 1277
rect 32961 1213 32973 1225
rect 33007 1213 33019 1225
rect 32961 1161 32964 1213
rect 33016 1161 33019 1213
rect 32961 1147 33019 1161
rect 33057 3133 33115 3147
rect 33057 3081 33060 3133
rect 33112 3081 33115 3133
rect 33057 3069 33069 3081
rect 33103 3069 33115 3081
rect 33057 3017 33060 3069
rect 33112 3017 33115 3069
rect 33057 3005 33069 3017
rect 33103 3005 33115 3017
rect 33057 2953 33060 3005
rect 33112 2953 33115 3005
rect 33057 2941 33069 2953
rect 33103 2941 33115 2953
rect 33057 2889 33060 2941
rect 33112 2889 33115 2941
rect 33057 2884 33115 2889
rect 33057 2877 33069 2884
rect 33103 2877 33115 2884
rect 33057 2825 33060 2877
rect 33112 2825 33115 2877
rect 33057 2813 33115 2825
rect 33057 2761 33060 2813
rect 33112 2761 33115 2813
rect 33057 2749 33115 2761
rect 33057 2697 33060 2749
rect 33112 2697 33115 2749
rect 33057 2685 33115 2697
rect 33057 2633 33060 2685
rect 33112 2633 33115 2685
rect 33057 2621 33115 2633
rect 33057 2569 33060 2621
rect 33112 2569 33115 2621
rect 33057 2562 33069 2569
rect 33103 2562 33115 2569
rect 33057 2557 33115 2562
rect 33057 2505 33060 2557
rect 33112 2505 33115 2557
rect 33057 2493 33069 2505
rect 33103 2493 33115 2505
rect 33057 2441 33060 2493
rect 33112 2441 33115 2493
rect 33057 2429 33069 2441
rect 33103 2429 33115 2441
rect 33057 2377 33060 2429
rect 33112 2377 33115 2429
rect 33057 2365 33069 2377
rect 33103 2365 33115 2377
rect 33057 2313 33060 2365
rect 33112 2313 33115 2365
rect 33057 2308 33115 2313
rect 33057 2301 33069 2308
rect 33103 2301 33115 2308
rect 33057 2249 33060 2301
rect 33112 2249 33115 2301
rect 33057 2237 33115 2249
rect 33057 2185 33060 2237
rect 33112 2185 33115 2237
rect 33057 2173 33115 2185
rect 33057 2121 33060 2173
rect 33112 2121 33115 2173
rect 33057 2109 33115 2121
rect 33057 2057 33060 2109
rect 33112 2057 33115 2109
rect 33057 2045 33115 2057
rect 33057 1993 33060 2045
rect 33112 1993 33115 2045
rect 33057 1986 33069 1993
rect 33103 1986 33115 1993
rect 33057 1981 33115 1986
rect 33057 1929 33060 1981
rect 33112 1929 33115 1981
rect 33057 1917 33069 1929
rect 33103 1917 33115 1929
rect 33057 1865 33060 1917
rect 33112 1865 33115 1917
rect 33057 1853 33069 1865
rect 33103 1853 33115 1865
rect 33057 1801 33060 1853
rect 33112 1801 33115 1853
rect 33057 1789 33069 1801
rect 33103 1789 33115 1801
rect 33057 1737 33060 1789
rect 33112 1737 33115 1789
rect 33057 1732 33115 1737
rect 33057 1725 33069 1732
rect 33103 1725 33115 1732
rect 33057 1673 33060 1725
rect 33112 1673 33115 1725
rect 33057 1661 33115 1673
rect 33057 1609 33060 1661
rect 33112 1609 33115 1661
rect 33057 1597 33115 1609
rect 33057 1545 33060 1597
rect 33112 1545 33115 1597
rect 33057 1533 33115 1545
rect 33057 1481 33060 1533
rect 33112 1481 33115 1533
rect 33057 1469 33115 1481
rect 33057 1417 33060 1469
rect 33112 1417 33115 1469
rect 33057 1410 33069 1417
rect 33103 1410 33115 1417
rect 33057 1405 33115 1410
rect 33057 1353 33060 1405
rect 33112 1353 33115 1405
rect 33057 1341 33069 1353
rect 33103 1341 33115 1353
rect 33057 1289 33060 1341
rect 33112 1289 33115 1341
rect 33057 1277 33069 1289
rect 33103 1277 33115 1289
rect 33057 1225 33060 1277
rect 33112 1225 33115 1277
rect 33057 1213 33069 1225
rect 33103 1213 33115 1225
rect 33057 1161 33060 1213
rect 33112 1161 33115 1213
rect 33057 1147 33115 1161
rect 33156 3133 33208 3147
rect 33156 3069 33165 3081
rect 33199 3069 33208 3081
rect 33156 3005 33165 3017
rect 33199 3005 33208 3017
rect 33156 2941 33165 2953
rect 33199 2941 33208 2953
rect 33156 2884 33208 2889
rect 33156 2877 33165 2884
rect 33199 2877 33208 2884
rect 33156 2813 33208 2825
rect 33156 2749 33208 2761
rect 33156 2685 33208 2697
rect 33156 2621 33208 2633
rect 33156 2562 33165 2569
rect 33199 2562 33208 2569
rect 33156 2557 33208 2562
rect 33156 2493 33165 2505
rect 33199 2493 33208 2505
rect 33156 2429 33165 2441
rect 33199 2429 33208 2441
rect 33156 2365 33165 2377
rect 33199 2365 33208 2377
rect 33156 2308 33208 2313
rect 33156 2301 33165 2308
rect 33199 2301 33208 2308
rect 33156 2237 33208 2249
rect 33156 2173 33208 2185
rect 33156 2109 33208 2121
rect 33156 2045 33208 2057
rect 33156 1986 33165 1993
rect 33199 1986 33208 1993
rect 33156 1981 33208 1986
rect 33156 1917 33165 1929
rect 33199 1917 33208 1929
rect 33156 1853 33165 1865
rect 33199 1853 33208 1865
rect 33156 1789 33165 1801
rect 33199 1789 33208 1801
rect 33156 1732 33208 1737
rect 33156 1725 33165 1732
rect 33199 1725 33208 1732
rect 33156 1661 33208 1673
rect 33156 1597 33208 1609
rect 33156 1533 33208 1545
rect 33156 1469 33208 1481
rect 33156 1410 33165 1417
rect 33199 1410 33208 1417
rect 33156 1405 33208 1410
rect 33156 1341 33165 1353
rect 33199 1341 33208 1353
rect 33156 1277 33165 1289
rect 33199 1277 33208 1289
rect 33156 1213 33165 1225
rect 33199 1213 33208 1225
rect 33156 1147 33208 1161
rect 33249 3133 33307 3147
rect 33249 3081 33252 3133
rect 33304 3081 33307 3133
rect 33249 3069 33261 3081
rect 33295 3069 33307 3081
rect 33249 3017 33252 3069
rect 33304 3017 33307 3069
rect 33249 3005 33261 3017
rect 33295 3005 33307 3017
rect 33249 2953 33252 3005
rect 33304 2953 33307 3005
rect 33249 2941 33261 2953
rect 33295 2941 33307 2953
rect 33249 2889 33252 2941
rect 33304 2889 33307 2941
rect 33249 2884 33307 2889
rect 33249 2877 33261 2884
rect 33295 2877 33307 2884
rect 33249 2825 33252 2877
rect 33304 2825 33307 2877
rect 33249 2813 33307 2825
rect 33249 2761 33252 2813
rect 33304 2761 33307 2813
rect 33249 2749 33307 2761
rect 33249 2697 33252 2749
rect 33304 2697 33307 2749
rect 33249 2685 33307 2697
rect 33249 2633 33252 2685
rect 33304 2633 33307 2685
rect 33249 2621 33307 2633
rect 33249 2569 33252 2621
rect 33304 2569 33307 2621
rect 33249 2562 33261 2569
rect 33295 2562 33307 2569
rect 33249 2557 33307 2562
rect 33249 2505 33252 2557
rect 33304 2505 33307 2557
rect 33249 2493 33261 2505
rect 33295 2493 33307 2505
rect 33249 2441 33252 2493
rect 33304 2441 33307 2493
rect 33249 2429 33261 2441
rect 33295 2429 33307 2441
rect 33249 2377 33252 2429
rect 33304 2377 33307 2429
rect 33249 2365 33261 2377
rect 33295 2365 33307 2377
rect 33249 2313 33252 2365
rect 33304 2313 33307 2365
rect 33249 2308 33307 2313
rect 33249 2301 33261 2308
rect 33295 2301 33307 2308
rect 33249 2249 33252 2301
rect 33304 2249 33307 2301
rect 33249 2237 33307 2249
rect 33249 2185 33252 2237
rect 33304 2185 33307 2237
rect 33249 2173 33307 2185
rect 33249 2121 33252 2173
rect 33304 2121 33307 2173
rect 33249 2109 33307 2121
rect 33249 2057 33252 2109
rect 33304 2057 33307 2109
rect 33249 2045 33307 2057
rect 33249 1993 33252 2045
rect 33304 1993 33307 2045
rect 33249 1986 33261 1993
rect 33295 1986 33307 1993
rect 33249 1981 33307 1986
rect 33249 1929 33252 1981
rect 33304 1929 33307 1981
rect 33249 1917 33261 1929
rect 33295 1917 33307 1929
rect 33249 1865 33252 1917
rect 33304 1865 33307 1917
rect 33249 1853 33261 1865
rect 33295 1853 33307 1865
rect 33249 1801 33252 1853
rect 33304 1801 33307 1853
rect 33249 1789 33261 1801
rect 33295 1789 33307 1801
rect 33249 1737 33252 1789
rect 33304 1737 33307 1789
rect 33249 1732 33307 1737
rect 33249 1725 33261 1732
rect 33295 1725 33307 1732
rect 33249 1673 33252 1725
rect 33304 1673 33307 1725
rect 33249 1661 33307 1673
rect 33249 1609 33252 1661
rect 33304 1609 33307 1661
rect 33249 1597 33307 1609
rect 33249 1545 33252 1597
rect 33304 1545 33307 1597
rect 33249 1533 33307 1545
rect 33249 1481 33252 1533
rect 33304 1481 33307 1533
rect 33249 1469 33307 1481
rect 33249 1417 33252 1469
rect 33304 1417 33307 1469
rect 33249 1410 33261 1417
rect 33295 1410 33307 1417
rect 33249 1405 33307 1410
rect 33249 1353 33252 1405
rect 33304 1353 33307 1405
rect 33249 1341 33261 1353
rect 33295 1341 33307 1353
rect 33249 1289 33252 1341
rect 33304 1289 33307 1341
rect 33249 1277 33261 1289
rect 33295 1277 33307 1289
rect 33249 1225 33252 1277
rect 33304 1225 33307 1277
rect 33249 1213 33261 1225
rect 33295 1213 33307 1225
rect 33249 1161 33252 1213
rect 33304 1161 33307 1213
rect 33249 1147 33307 1161
rect 33345 3133 33403 3147
rect 33345 3081 33348 3133
rect 33400 3081 33403 3133
rect 33345 3069 33357 3081
rect 33391 3069 33403 3081
rect 33345 3017 33348 3069
rect 33400 3017 33403 3069
rect 33345 3005 33357 3017
rect 33391 3005 33403 3017
rect 33345 2953 33348 3005
rect 33400 2953 33403 3005
rect 33345 2941 33357 2953
rect 33391 2941 33403 2953
rect 33345 2889 33348 2941
rect 33400 2889 33403 2941
rect 33345 2884 33403 2889
rect 33345 2877 33357 2884
rect 33391 2877 33403 2884
rect 33345 2825 33348 2877
rect 33400 2825 33403 2877
rect 33345 2813 33403 2825
rect 33345 2761 33348 2813
rect 33400 2761 33403 2813
rect 33345 2749 33403 2761
rect 33345 2697 33348 2749
rect 33400 2697 33403 2749
rect 33345 2685 33403 2697
rect 33345 2633 33348 2685
rect 33400 2633 33403 2685
rect 33345 2621 33403 2633
rect 33345 2569 33348 2621
rect 33400 2569 33403 2621
rect 33345 2562 33357 2569
rect 33391 2562 33403 2569
rect 33345 2557 33403 2562
rect 33345 2505 33348 2557
rect 33400 2505 33403 2557
rect 33345 2493 33357 2505
rect 33391 2493 33403 2505
rect 33345 2441 33348 2493
rect 33400 2441 33403 2493
rect 33345 2429 33357 2441
rect 33391 2429 33403 2441
rect 33345 2377 33348 2429
rect 33400 2377 33403 2429
rect 33345 2365 33357 2377
rect 33391 2365 33403 2377
rect 33345 2313 33348 2365
rect 33400 2313 33403 2365
rect 33345 2308 33403 2313
rect 33345 2301 33357 2308
rect 33391 2301 33403 2308
rect 33345 2249 33348 2301
rect 33400 2249 33403 2301
rect 33345 2237 33403 2249
rect 33345 2185 33348 2237
rect 33400 2185 33403 2237
rect 33345 2173 33403 2185
rect 33345 2121 33348 2173
rect 33400 2121 33403 2173
rect 33345 2109 33403 2121
rect 33345 2057 33348 2109
rect 33400 2057 33403 2109
rect 33345 2045 33403 2057
rect 33345 1993 33348 2045
rect 33400 1993 33403 2045
rect 33345 1986 33357 1993
rect 33391 1986 33403 1993
rect 33345 1981 33403 1986
rect 33345 1929 33348 1981
rect 33400 1929 33403 1981
rect 33345 1917 33357 1929
rect 33391 1917 33403 1929
rect 33345 1865 33348 1917
rect 33400 1865 33403 1917
rect 33345 1853 33357 1865
rect 33391 1853 33403 1865
rect 33345 1801 33348 1853
rect 33400 1801 33403 1853
rect 33345 1789 33357 1801
rect 33391 1789 33403 1801
rect 33345 1737 33348 1789
rect 33400 1737 33403 1789
rect 33345 1732 33403 1737
rect 33345 1725 33357 1732
rect 33391 1725 33403 1732
rect 33345 1673 33348 1725
rect 33400 1673 33403 1725
rect 33345 1661 33403 1673
rect 33345 1609 33348 1661
rect 33400 1609 33403 1661
rect 33345 1597 33403 1609
rect 33345 1545 33348 1597
rect 33400 1545 33403 1597
rect 33345 1533 33403 1545
rect 33345 1481 33348 1533
rect 33400 1481 33403 1533
rect 33345 1469 33403 1481
rect 33345 1417 33348 1469
rect 33400 1417 33403 1469
rect 33345 1410 33357 1417
rect 33391 1410 33403 1417
rect 33345 1405 33403 1410
rect 33345 1353 33348 1405
rect 33400 1353 33403 1405
rect 33345 1341 33357 1353
rect 33391 1341 33403 1353
rect 33345 1289 33348 1341
rect 33400 1289 33403 1341
rect 33345 1277 33357 1289
rect 33391 1277 33403 1289
rect 33345 1225 33348 1277
rect 33400 1225 33403 1277
rect 33345 1213 33357 1225
rect 33391 1213 33403 1225
rect 33345 1161 33348 1213
rect 33400 1161 33403 1213
rect 33345 1147 33403 1161
rect 33441 3133 33499 3147
rect 33441 3081 33444 3133
rect 33496 3081 33499 3133
rect 33441 3069 33453 3081
rect 33487 3069 33499 3081
rect 33441 3017 33444 3069
rect 33496 3017 33499 3069
rect 33441 3005 33453 3017
rect 33487 3005 33499 3017
rect 33441 2953 33444 3005
rect 33496 2953 33499 3005
rect 33441 2941 33453 2953
rect 33487 2941 33499 2953
rect 33441 2889 33444 2941
rect 33496 2889 33499 2941
rect 33441 2884 33499 2889
rect 33441 2877 33453 2884
rect 33487 2877 33499 2884
rect 33441 2825 33444 2877
rect 33496 2825 33499 2877
rect 33441 2813 33499 2825
rect 33441 2761 33444 2813
rect 33496 2761 33499 2813
rect 33441 2749 33499 2761
rect 33441 2697 33444 2749
rect 33496 2697 33499 2749
rect 33441 2685 33499 2697
rect 33441 2633 33444 2685
rect 33496 2633 33499 2685
rect 33441 2621 33499 2633
rect 33441 2569 33444 2621
rect 33496 2569 33499 2621
rect 33441 2562 33453 2569
rect 33487 2562 33499 2569
rect 33441 2557 33499 2562
rect 33441 2505 33444 2557
rect 33496 2505 33499 2557
rect 33441 2493 33453 2505
rect 33487 2493 33499 2505
rect 33441 2441 33444 2493
rect 33496 2441 33499 2493
rect 33441 2429 33453 2441
rect 33487 2429 33499 2441
rect 33441 2377 33444 2429
rect 33496 2377 33499 2429
rect 33441 2365 33453 2377
rect 33487 2365 33499 2377
rect 33441 2313 33444 2365
rect 33496 2313 33499 2365
rect 33441 2308 33499 2313
rect 33441 2301 33453 2308
rect 33487 2301 33499 2308
rect 33441 2249 33444 2301
rect 33496 2249 33499 2301
rect 33441 2237 33499 2249
rect 33441 2185 33444 2237
rect 33496 2185 33499 2237
rect 33441 2173 33499 2185
rect 33441 2121 33444 2173
rect 33496 2121 33499 2173
rect 33441 2109 33499 2121
rect 33441 2057 33444 2109
rect 33496 2057 33499 2109
rect 33441 2045 33499 2057
rect 33441 1993 33444 2045
rect 33496 1993 33499 2045
rect 33441 1986 33453 1993
rect 33487 1986 33499 1993
rect 33441 1981 33499 1986
rect 33441 1929 33444 1981
rect 33496 1929 33499 1981
rect 33441 1917 33453 1929
rect 33487 1917 33499 1929
rect 33441 1865 33444 1917
rect 33496 1865 33499 1917
rect 33441 1853 33453 1865
rect 33487 1853 33499 1865
rect 33441 1801 33444 1853
rect 33496 1801 33499 1853
rect 33441 1789 33453 1801
rect 33487 1789 33499 1801
rect 33441 1737 33444 1789
rect 33496 1737 33499 1789
rect 33441 1732 33499 1737
rect 33441 1725 33453 1732
rect 33487 1725 33499 1732
rect 33441 1673 33444 1725
rect 33496 1673 33499 1725
rect 33441 1661 33499 1673
rect 33441 1609 33444 1661
rect 33496 1609 33499 1661
rect 33441 1597 33499 1609
rect 33441 1545 33444 1597
rect 33496 1545 33499 1597
rect 33441 1533 33499 1545
rect 33441 1481 33444 1533
rect 33496 1481 33499 1533
rect 33441 1469 33499 1481
rect 33441 1417 33444 1469
rect 33496 1417 33499 1469
rect 33441 1410 33453 1417
rect 33487 1410 33499 1417
rect 33441 1405 33499 1410
rect 33441 1353 33444 1405
rect 33496 1353 33499 1405
rect 33441 1341 33453 1353
rect 33487 1341 33499 1353
rect 33441 1289 33444 1341
rect 33496 1289 33499 1341
rect 33441 1277 33453 1289
rect 33487 1277 33499 1289
rect 33441 1225 33444 1277
rect 33496 1225 33499 1277
rect 33441 1213 33453 1225
rect 33487 1213 33499 1225
rect 33441 1161 33444 1213
rect 33496 1161 33499 1213
rect 33441 1147 33499 1161
rect 33540 3133 33592 3147
rect 33540 3069 33549 3081
rect 33583 3069 33592 3081
rect 33540 3005 33549 3017
rect 33583 3005 33592 3017
rect 33540 2941 33549 2953
rect 33583 2941 33592 2953
rect 33540 2884 33592 2889
rect 33540 2877 33549 2884
rect 33583 2877 33592 2884
rect 33540 2813 33592 2825
rect 33540 2749 33592 2761
rect 33540 2685 33592 2697
rect 33540 2621 33592 2633
rect 33540 2562 33549 2569
rect 33583 2562 33592 2569
rect 33540 2557 33592 2562
rect 33540 2493 33549 2505
rect 33583 2493 33592 2505
rect 33540 2429 33549 2441
rect 33583 2429 33592 2441
rect 33540 2365 33549 2377
rect 33583 2365 33592 2377
rect 33540 2308 33592 2313
rect 33540 2301 33549 2308
rect 33583 2301 33592 2308
rect 33540 2237 33592 2249
rect 33540 2173 33592 2185
rect 33540 2109 33592 2121
rect 33540 2045 33592 2057
rect 33540 1986 33549 1993
rect 33583 1986 33592 1993
rect 33540 1981 33592 1986
rect 33540 1917 33549 1929
rect 33583 1917 33592 1929
rect 33540 1853 33549 1865
rect 33583 1853 33592 1865
rect 33540 1789 33549 1801
rect 33583 1789 33592 1801
rect 33540 1732 33592 1737
rect 33540 1725 33549 1732
rect 33583 1725 33592 1732
rect 33540 1661 33592 1673
rect 33540 1597 33592 1609
rect 33540 1533 33592 1545
rect 33540 1469 33592 1481
rect 33540 1410 33549 1417
rect 33583 1410 33592 1417
rect 33540 1405 33592 1410
rect 33540 1341 33549 1353
rect 33583 1341 33592 1353
rect 33540 1277 33549 1289
rect 33583 1277 33592 1289
rect 33540 1213 33549 1225
rect 33583 1213 33592 1225
rect 33540 1147 33592 1161
rect 33633 3133 33691 3147
rect 33633 3081 33636 3133
rect 33688 3081 33691 3133
rect 33633 3069 33645 3081
rect 33679 3069 33691 3081
rect 33633 3017 33636 3069
rect 33688 3017 33691 3069
rect 33633 3005 33645 3017
rect 33679 3005 33691 3017
rect 33633 2953 33636 3005
rect 33688 2953 33691 3005
rect 33633 2941 33645 2953
rect 33679 2941 33691 2953
rect 33633 2889 33636 2941
rect 33688 2889 33691 2941
rect 33633 2884 33691 2889
rect 33633 2877 33645 2884
rect 33679 2877 33691 2884
rect 33633 2825 33636 2877
rect 33688 2825 33691 2877
rect 33633 2813 33691 2825
rect 33633 2761 33636 2813
rect 33688 2761 33691 2813
rect 33633 2749 33691 2761
rect 33633 2697 33636 2749
rect 33688 2697 33691 2749
rect 33633 2685 33691 2697
rect 33633 2633 33636 2685
rect 33688 2633 33691 2685
rect 33633 2621 33691 2633
rect 33633 2569 33636 2621
rect 33688 2569 33691 2621
rect 33633 2562 33645 2569
rect 33679 2562 33691 2569
rect 33633 2557 33691 2562
rect 33633 2505 33636 2557
rect 33688 2505 33691 2557
rect 33633 2493 33645 2505
rect 33679 2493 33691 2505
rect 33633 2441 33636 2493
rect 33688 2441 33691 2493
rect 33633 2429 33645 2441
rect 33679 2429 33691 2441
rect 33633 2377 33636 2429
rect 33688 2377 33691 2429
rect 33633 2365 33645 2377
rect 33679 2365 33691 2377
rect 33633 2313 33636 2365
rect 33688 2313 33691 2365
rect 33633 2308 33691 2313
rect 33633 2301 33645 2308
rect 33679 2301 33691 2308
rect 33633 2249 33636 2301
rect 33688 2249 33691 2301
rect 33633 2237 33691 2249
rect 33633 2185 33636 2237
rect 33688 2185 33691 2237
rect 33633 2173 33691 2185
rect 33633 2121 33636 2173
rect 33688 2121 33691 2173
rect 33633 2109 33691 2121
rect 33633 2057 33636 2109
rect 33688 2057 33691 2109
rect 33633 2045 33691 2057
rect 33633 1993 33636 2045
rect 33688 1993 33691 2045
rect 33633 1986 33645 1993
rect 33679 1986 33691 1993
rect 33633 1981 33691 1986
rect 33633 1929 33636 1981
rect 33688 1929 33691 1981
rect 33633 1917 33645 1929
rect 33679 1917 33691 1929
rect 33633 1865 33636 1917
rect 33688 1865 33691 1917
rect 33633 1853 33645 1865
rect 33679 1853 33691 1865
rect 33633 1801 33636 1853
rect 33688 1801 33691 1853
rect 33633 1789 33645 1801
rect 33679 1789 33691 1801
rect 33633 1737 33636 1789
rect 33688 1737 33691 1789
rect 33633 1732 33691 1737
rect 33633 1725 33645 1732
rect 33679 1725 33691 1732
rect 33633 1673 33636 1725
rect 33688 1673 33691 1725
rect 33633 1661 33691 1673
rect 33633 1609 33636 1661
rect 33688 1609 33691 1661
rect 33633 1597 33691 1609
rect 33633 1545 33636 1597
rect 33688 1545 33691 1597
rect 33633 1533 33691 1545
rect 33633 1481 33636 1533
rect 33688 1481 33691 1533
rect 33633 1469 33691 1481
rect 33633 1417 33636 1469
rect 33688 1417 33691 1469
rect 33633 1410 33645 1417
rect 33679 1410 33691 1417
rect 33633 1405 33691 1410
rect 33633 1353 33636 1405
rect 33688 1353 33691 1405
rect 33633 1341 33645 1353
rect 33679 1341 33691 1353
rect 33633 1289 33636 1341
rect 33688 1289 33691 1341
rect 33633 1277 33645 1289
rect 33679 1277 33691 1289
rect 33633 1225 33636 1277
rect 33688 1225 33691 1277
rect 33633 1213 33645 1225
rect 33679 1213 33691 1225
rect 33633 1161 33636 1213
rect 33688 1161 33691 1213
rect 33633 1147 33691 1161
rect 33729 3133 33787 3147
rect 33729 3081 33732 3133
rect 33784 3081 33787 3133
rect 33729 3069 33741 3081
rect 33775 3069 33787 3081
rect 33729 3017 33732 3069
rect 33784 3017 33787 3069
rect 33729 3005 33741 3017
rect 33775 3005 33787 3017
rect 33729 2953 33732 3005
rect 33784 2953 33787 3005
rect 33729 2941 33741 2953
rect 33775 2941 33787 2953
rect 33729 2889 33732 2941
rect 33784 2889 33787 2941
rect 33729 2884 33787 2889
rect 33729 2877 33741 2884
rect 33775 2877 33787 2884
rect 33729 2825 33732 2877
rect 33784 2825 33787 2877
rect 33729 2813 33787 2825
rect 33729 2761 33732 2813
rect 33784 2761 33787 2813
rect 33729 2749 33787 2761
rect 33729 2697 33732 2749
rect 33784 2697 33787 2749
rect 33729 2685 33787 2697
rect 33729 2633 33732 2685
rect 33784 2633 33787 2685
rect 33729 2621 33787 2633
rect 33729 2569 33732 2621
rect 33784 2569 33787 2621
rect 33729 2562 33741 2569
rect 33775 2562 33787 2569
rect 33729 2557 33787 2562
rect 33729 2505 33732 2557
rect 33784 2505 33787 2557
rect 33729 2493 33741 2505
rect 33775 2493 33787 2505
rect 33729 2441 33732 2493
rect 33784 2441 33787 2493
rect 33729 2429 33741 2441
rect 33775 2429 33787 2441
rect 33729 2377 33732 2429
rect 33784 2377 33787 2429
rect 33729 2365 33741 2377
rect 33775 2365 33787 2377
rect 33729 2313 33732 2365
rect 33784 2313 33787 2365
rect 33729 2308 33787 2313
rect 33729 2301 33741 2308
rect 33775 2301 33787 2308
rect 33729 2249 33732 2301
rect 33784 2249 33787 2301
rect 33729 2237 33787 2249
rect 33729 2185 33732 2237
rect 33784 2185 33787 2237
rect 33729 2173 33787 2185
rect 33729 2121 33732 2173
rect 33784 2121 33787 2173
rect 33729 2109 33787 2121
rect 33729 2057 33732 2109
rect 33784 2057 33787 2109
rect 33729 2045 33787 2057
rect 33729 1993 33732 2045
rect 33784 1993 33787 2045
rect 33729 1986 33741 1993
rect 33775 1986 33787 1993
rect 33729 1981 33787 1986
rect 33729 1929 33732 1981
rect 33784 1929 33787 1981
rect 33729 1917 33741 1929
rect 33775 1917 33787 1929
rect 33729 1865 33732 1917
rect 33784 1865 33787 1917
rect 33729 1853 33741 1865
rect 33775 1853 33787 1865
rect 33729 1801 33732 1853
rect 33784 1801 33787 1853
rect 33729 1789 33741 1801
rect 33775 1789 33787 1801
rect 33729 1737 33732 1789
rect 33784 1737 33787 1789
rect 33729 1732 33787 1737
rect 33729 1725 33741 1732
rect 33775 1725 33787 1732
rect 33729 1673 33732 1725
rect 33784 1673 33787 1725
rect 33729 1661 33787 1673
rect 33729 1609 33732 1661
rect 33784 1609 33787 1661
rect 33729 1597 33787 1609
rect 33729 1545 33732 1597
rect 33784 1545 33787 1597
rect 33729 1533 33787 1545
rect 33729 1481 33732 1533
rect 33784 1481 33787 1533
rect 33729 1469 33787 1481
rect 33729 1417 33732 1469
rect 33784 1417 33787 1469
rect 33729 1410 33741 1417
rect 33775 1410 33787 1417
rect 33729 1405 33787 1410
rect 33729 1353 33732 1405
rect 33784 1353 33787 1405
rect 33729 1341 33741 1353
rect 33775 1341 33787 1353
rect 33729 1289 33732 1341
rect 33784 1289 33787 1341
rect 33729 1277 33741 1289
rect 33775 1277 33787 1289
rect 33729 1225 33732 1277
rect 33784 1225 33787 1277
rect 33729 1213 33741 1225
rect 33775 1213 33787 1225
rect 33729 1161 33732 1213
rect 33784 1161 33787 1213
rect 33729 1147 33787 1161
rect 33825 3133 33883 3147
rect 33825 3081 33828 3133
rect 33880 3081 33883 3133
rect 33825 3069 33837 3081
rect 33871 3069 33883 3081
rect 33825 3017 33828 3069
rect 33880 3017 33883 3069
rect 33825 3005 33837 3017
rect 33871 3005 33883 3017
rect 33825 2953 33828 3005
rect 33880 2953 33883 3005
rect 33825 2941 33837 2953
rect 33871 2941 33883 2953
rect 33825 2889 33828 2941
rect 33880 2889 33883 2941
rect 33825 2884 33883 2889
rect 33825 2877 33837 2884
rect 33871 2877 33883 2884
rect 33825 2825 33828 2877
rect 33880 2825 33883 2877
rect 33825 2813 33883 2825
rect 33825 2761 33828 2813
rect 33880 2761 33883 2813
rect 33825 2749 33883 2761
rect 33825 2697 33828 2749
rect 33880 2697 33883 2749
rect 33825 2685 33883 2697
rect 33825 2633 33828 2685
rect 33880 2633 33883 2685
rect 33825 2621 33883 2633
rect 33825 2569 33828 2621
rect 33880 2569 33883 2621
rect 33825 2562 33837 2569
rect 33871 2562 33883 2569
rect 33825 2557 33883 2562
rect 33825 2505 33828 2557
rect 33880 2505 33883 2557
rect 33825 2493 33837 2505
rect 33871 2493 33883 2505
rect 33825 2441 33828 2493
rect 33880 2441 33883 2493
rect 33825 2429 33837 2441
rect 33871 2429 33883 2441
rect 33825 2377 33828 2429
rect 33880 2377 33883 2429
rect 33825 2365 33837 2377
rect 33871 2365 33883 2377
rect 33825 2313 33828 2365
rect 33880 2313 33883 2365
rect 33825 2308 33883 2313
rect 33825 2301 33837 2308
rect 33871 2301 33883 2308
rect 33825 2249 33828 2301
rect 33880 2249 33883 2301
rect 33825 2237 33883 2249
rect 33825 2185 33828 2237
rect 33880 2185 33883 2237
rect 33825 2173 33883 2185
rect 33825 2121 33828 2173
rect 33880 2121 33883 2173
rect 33825 2109 33883 2121
rect 33825 2057 33828 2109
rect 33880 2057 33883 2109
rect 33825 2045 33883 2057
rect 33825 1993 33828 2045
rect 33880 1993 33883 2045
rect 33825 1986 33837 1993
rect 33871 1986 33883 1993
rect 33825 1981 33883 1986
rect 33825 1929 33828 1981
rect 33880 1929 33883 1981
rect 33825 1917 33837 1929
rect 33871 1917 33883 1929
rect 33825 1865 33828 1917
rect 33880 1865 33883 1917
rect 33825 1853 33837 1865
rect 33871 1853 33883 1865
rect 33825 1801 33828 1853
rect 33880 1801 33883 1853
rect 33825 1789 33837 1801
rect 33871 1789 33883 1801
rect 33825 1737 33828 1789
rect 33880 1737 33883 1789
rect 33825 1732 33883 1737
rect 33825 1725 33837 1732
rect 33871 1725 33883 1732
rect 33825 1673 33828 1725
rect 33880 1673 33883 1725
rect 33825 1661 33883 1673
rect 33825 1609 33828 1661
rect 33880 1609 33883 1661
rect 33825 1597 33883 1609
rect 33825 1545 33828 1597
rect 33880 1545 33883 1597
rect 33825 1533 33883 1545
rect 33825 1481 33828 1533
rect 33880 1481 33883 1533
rect 33825 1469 33883 1481
rect 33825 1417 33828 1469
rect 33880 1417 33883 1469
rect 33825 1410 33837 1417
rect 33871 1410 33883 1417
rect 33825 1405 33883 1410
rect 33825 1353 33828 1405
rect 33880 1353 33883 1405
rect 33825 1341 33837 1353
rect 33871 1341 33883 1353
rect 33825 1289 33828 1341
rect 33880 1289 33883 1341
rect 33825 1277 33837 1289
rect 33871 1277 33883 1289
rect 33825 1225 33828 1277
rect 33880 1225 33883 1277
rect 33825 1213 33837 1225
rect 33871 1213 33883 1225
rect 33825 1161 33828 1213
rect 33880 1161 33883 1213
rect 33825 1147 33883 1161
rect 33924 3133 33976 3147
rect 33924 3069 33933 3081
rect 33967 3069 33976 3081
rect 33924 3005 33933 3017
rect 33967 3005 33976 3017
rect 33924 2941 33933 2953
rect 33967 2941 33976 2953
rect 33924 2884 33976 2889
rect 33924 2877 33933 2884
rect 33967 2877 33976 2884
rect 33924 2813 33976 2825
rect 33924 2749 33976 2761
rect 33924 2685 33976 2697
rect 33924 2621 33976 2633
rect 33924 2562 33933 2569
rect 33967 2562 33976 2569
rect 33924 2557 33976 2562
rect 33924 2493 33933 2505
rect 33967 2493 33976 2505
rect 33924 2429 33933 2441
rect 33967 2429 33976 2441
rect 33924 2365 33933 2377
rect 33967 2365 33976 2377
rect 33924 2308 33976 2313
rect 33924 2301 33933 2308
rect 33967 2301 33976 2308
rect 33924 2237 33976 2249
rect 33924 2173 33976 2185
rect 33924 2109 33976 2121
rect 33924 2045 33976 2057
rect 33924 1986 33933 1993
rect 33967 1986 33976 1993
rect 33924 1981 33976 1986
rect 33924 1917 33933 1929
rect 33967 1917 33976 1929
rect 33924 1853 33933 1865
rect 33967 1853 33976 1865
rect 33924 1789 33933 1801
rect 33967 1789 33976 1801
rect 33924 1732 33976 1737
rect 33924 1725 33933 1732
rect 33967 1725 33976 1732
rect 33924 1661 33976 1673
rect 33924 1597 33976 1609
rect 33924 1533 33976 1545
rect 33924 1469 33976 1481
rect 33924 1410 33933 1417
rect 33967 1410 33976 1417
rect 33924 1405 33976 1410
rect 33924 1341 33933 1353
rect 33967 1341 33976 1353
rect 33924 1277 33933 1289
rect 33967 1277 33976 1289
rect 33924 1213 33933 1225
rect 33967 1213 33976 1225
rect 33924 1147 33976 1161
rect 34017 3133 34075 3147
rect 34017 3081 34020 3133
rect 34072 3081 34075 3133
rect 34017 3069 34029 3081
rect 34063 3069 34075 3081
rect 34017 3017 34020 3069
rect 34072 3017 34075 3069
rect 34017 3005 34029 3017
rect 34063 3005 34075 3017
rect 34017 2953 34020 3005
rect 34072 2953 34075 3005
rect 34017 2941 34029 2953
rect 34063 2941 34075 2953
rect 34017 2889 34020 2941
rect 34072 2889 34075 2941
rect 34017 2884 34075 2889
rect 34017 2877 34029 2884
rect 34063 2877 34075 2884
rect 34017 2825 34020 2877
rect 34072 2825 34075 2877
rect 34017 2813 34075 2825
rect 34017 2761 34020 2813
rect 34072 2761 34075 2813
rect 34017 2749 34075 2761
rect 34017 2697 34020 2749
rect 34072 2697 34075 2749
rect 34017 2685 34075 2697
rect 34017 2633 34020 2685
rect 34072 2633 34075 2685
rect 34017 2621 34075 2633
rect 34017 2569 34020 2621
rect 34072 2569 34075 2621
rect 34017 2562 34029 2569
rect 34063 2562 34075 2569
rect 34017 2557 34075 2562
rect 34017 2505 34020 2557
rect 34072 2505 34075 2557
rect 34017 2493 34029 2505
rect 34063 2493 34075 2505
rect 34017 2441 34020 2493
rect 34072 2441 34075 2493
rect 34017 2429 34029 2441
rect 34063 2429 34075 2441
rect 34017 2377 34020 2429
rect 34072 2377 34075 2429
rect 34017 2365 34029 2377
rect 34063 2365 34075 2377
rect 34017 2313 34020 2365
rect 34072 2313 34075 2365
rect 34017 2308 34075 2313
rect 34017 2301 34029 2308
rect 34063 2301 34075 2308
rect 34017 2249 34020 2301
rect 34072 2249 34075 2301
rect 34017 2237 34075 2249
rect 34017 2185 34020 2237
rect 34072 2185 34075 2237
rect 34017 2173 34075 2185
rect 34017 2121 34020 2173
rect 34072 2121 34075 2173
rect 34017 2109 34075 2121
rect 34017 2057 34020 2109
rect 34072 2057 34075 2109
rect 34017 2045 34075 2057
rect 34017 1993 34020 2045
rect 34072 1993 34075 2045
rect 34017 1986 34029 1993
rect 34063 1986 34075 1993
rect 34017 1981 34075 1986
rect 34017 1929 34020 1981
rect 34072 1929 34075 1981
rect 34017 1917 34029 1929
rect 34063 1917 34075 1929
rect 34017 1865 34020 1917
rect 34072 1865 34075 1917
rect 34017 1853 34029 1865
rect 34063 1853 34075 1865
rect 34017 1801 34020 1853
rect 34072 1801 34075 1853
rect 34017 1789 34029 1801
rect 34063 1789 34075 1801
rect 34017 1737 34020 1789
rect 34072 1737 34075 1789
rect 34017 1732 34075 1737
rect 34017 1725 34029 1732
rect 34063 1725 34075 1732
rect 34017 1673 34020 1725
rect 34072 1673 34075 1725
rect 34017 1661 34075 1673
rect 34017 1609 34020 1661
rect 34072 1609 34075 1661
rect 34017 1597 34075 1609
rect 34017 1545 34020 1597
rect 34072 1545 34075 1597
rect 34017 1533 34075 1545
rect 34017 1481 34020 1533
rect 34072 1481 34075 1533
rect 34017 1469 34075 1481
rect 34017 1417 34020 1469
rect 34072 1417 34075 1469
rect 34017 1410 34029 1417
rect 34063 1410 34075 1417
rect 34017 1405 34075 1410
rect 34017 1353 34020 1405
rect 34072 1353 34075 1405
rect 34017 1341 34029 1353
rect 34063 1341 34075 1353
rect 34017 1289 34020 1341
rect 34072 1289 34075 1341
rect 34017 1277 34029 1289
rect 34063 1277 34075 1289
rect 34017 1225 34020 1277
rect 34072 1225 34075 1277
rect 34017 1213 34029 1225
rect 34063 1213 34075 1225
rect 34017 1161 34020 1213
rect 34072 1161 34075 1213
rect 34017 1147 34075 1161
rect 34113 3133 34171 3147
rect 34113 3081 34116 3133
rect 34168 3081 34171 3133
rect 34113 3069 34125 3081
rect 34159 3069 34171 3081
rect 34113 3017 34116 3069
rect 34168 3017 34171 3069
rect 34113 3005 34125 3017
rect 34159 3005 34171 3017
rect 34113 2953 34116 3005
rect 34168 2953 34171 3005
rect 34113 2941 34125 2953
rect 34159 2941 34171 2953
rect 34113 2889 34116 2941
rect 34168 2889 34171 2941
rect 34113 2884 34171 2889
rect 34113 2877 34125 2884
rect 34159 2877 34171 2884
rect 34113 2825 34116 2877
rect 34168 2825 34171 2877
rect 34113 2813 34171 2825
rect 34113 2761 34116 2813
rect 34168 2761 34171 2813
rect 34113 2749 34171 2761
rect 34113 2697 34116 2749
rect 34168 2697 34171 2749
rect 34113 2685 34171 2697
rect 34113 2633 34116 2685
rect 34168 2633 34171 2685
rect 34113 2621 34171 2633
rect 34113 2569 34116 2621
rect 34168 2569 34171 2621
rect 34113 2562 34125 2569
rect 34159 2562 34171 2569
rect 34113 2557 34171 2562
rect 34113 2505 34116 2557
rect 34168 2505 34171 2557
rect 34113 2493 34125 2505
rect 34159 2493 34171 2505
rect 34113 2441 34116 2493
rect 34168 2441 34171 2493
rect 34113 2429 34125 2441
rect 34159 2429 34171 2441
rect 34113 2377 34116 2429
rect 34168 2377 34171 2429
rect 34113 2365 34125 2377
rect 34159 2365 34171 2377
rect 34113 2313 34116 2365
rect 34168 2313 34171 2365
rect 34113 2308 34171 2313
rect 34113 2301 34125 2308
rect 34159 2301 34171 2308
rect 34113 2249 34116 2301
rect 34168 2249 34171 2301
rect 34113 2237 34171 2249
rect 34113 2185 34116 2237
rect 34168 2185 34171 2237
rect 34113 2173 34171 2185
rect 34113 2121 34116 2173
rect 34168 2121 34171 2173
rect 34113 2109 34171 2121
rect 34113 2057 34116 2109
rect 34168 2057 34171 2109
rect 34113 2045 34171 2057
rect 34113 1993 34116 2045
rect 34168 1993 34171 2045
rect 34113 1986 34125 1993
rect 34159 1986 34171 1993
rect 34113 1981 34171 1986
rect 34113 1929 34116 1981
rect 34168 1929 34171 1981
rect 34113 1917 34125 1929
rect 34159 1917 34171 1929
rect 34113 1865 34116 1917
rect 34168 1865 34171 1917
rect 34113 1853 34125 1865
rect 34159 1853 34171 1865
rect 34113 1801 34116 1853
rect 34168 1801 34171 1853
rect 34113 1789 34125 1801
rect 34159 1789 34171 1801
rect 34113 1737 34116 1789
rect 34168 1737 34171 1789
rect 34113 1732 34171 1737
rect 34113 1725 34125 1732
rect 34159 1725 34171 1732
rect 34113 1673 34116 1725
rect 34168 1673 34171 1725
rect 34113 1661 34171 1673
rect 34113 1609 34116 1661
rect 34168 1609 34171 1661
rect 34113 1597 34171 1609
rect 34113 1545 34116 1597
rect 34168 1545 34171 1597
rect 34113 1533 34171 1545
rect 34113 1481 34116 1533
rect 34168 1481 34171 1533
rect 34113 1469 34171 1481
rect 34113 1417 34116 1469
rect 34168 1417 34171 1469
rect 34113 1410 34125 1417
rect 34159 1410 34171 1417
rect 34113 1405 34171 1410
rect 34113 1353 34116 1405
rect 34168 1353 34171 1405
rect 34113 1341 34125 1353
rect 34159 1341 34171 1353
rect 34113 1289 34116 1341
rect 34168 1289 34171 1341
rect 34113 1277 34125 1289
rect 34159 1277 34171 1289
rect 34113 1225 34116 1277
rect 34168 1225 34171 1277
rect 34113 1213 34125 1225
rect 34159 1213 34171 1225
rect 34113 1161 34116 1213
rect 34168 1161 34171 1213
rect 34113 1147 34171 1161
rect 34209 3133 34267 3147
rect 34209 3081 34212 3133
rect 34264 3081 34267 3133
rect 34209 3069 34221 3081
rect 34255 3069 34267 3081
rect 34209 3017 34212 3069
rect 34264 3017 34267 3069
rect 34209 3005 34221 3017
rect 34255 3005 34267 3017
rect 34209 2953 34212 3005
rect 34264 2953 34267 3005
rect 34209 2941 34221 2953
rect 34255 2941 34267 2953
rect 34209 2889 34212 2941
rect 34264 2889 34267 2941
rect 34209 2884 34267 2889
rect 34209 2877 34221 2884
rect 34255 2877 34267 2884
rect 34209 2825 34212 2877
rect 34264 2825 34267 2877
rect 34209 2813 34267 2825
rect 34209 2761 34212 2813
rect 34264 2761 34267 2813
rect 34209 2749 34267 2761
rect 34209 2697 34212 2749
rect 34264 2697 34267 2749
rect 34209 2685 34267 2697
rect 34209 2633 34212 2685
rect 34264 2633 34267 2685
rect 34209 2621 34267 2633
rect 34209 2569 34212 2621
rect 34264 2569 34267 2621
rect 34209 2562 34221 2569
rect 34255 2562 34267 2569
rect 34209 2557 34267 2562
rect 34209 2505 34212 2557
rect 34264 2505 34267 2557
rect 34209 2493 34221 2505
rect 34255 2493 34267 2505
rect 34209 2441 34212 2493
rect 34264 2441 34267 2493
rect 34209 2429 34221 2441
rect 34255 2429 34267 2441
rect 34209 2377 34212 2429
rect 34264 2377 34267 2429
rect 34209 2365 34221 2377
rect 34255 2365 34267 2377
rect 34209 2313 34212 2365
rect 34264 2313 34267 2365
rect 34209 2308 34267 2313
rect 34209 2301 34221 2308
rect 34255 2301 34267 2308
rect 34209 2249 34212 2301
rect 34264 2249 34267 2301
rect 34209 2237 34267 2249
rect 34209 2185 34212 2237
rect 34264 2185 34267 2237
rect 34209 2173 34267 2185
rect 34209 2121 34212 2173
rect 34264 2121 34267 2173
rect 34209 2109 34267 2121
rect 34209 2057 34212 2109
rect 34264 2057 34267 2109
rect 34209 2045 34267 2057
rect 34209 1993 34212 2045
rect 34264 1993 34267 2045
rect 34209 1986 34221 1993
rect 34255 1986 34267 1993
rect 34209 1981 34267 1986
rect 34209 1929 34212 1981
rect 34264 1929 34267 1981
rect 34209 1917 34221 1929
rect 34255 1917 34267 1929
rect 34209 1865 34212 1917
rect 34264 1865 34267 1917
rect 34209 1853 34221 1865
rect 34255 1853 34267 1865
rect 34209 1801 34212 1853
rect 34264 1801 34267 1853
rect 34209 1789 34221 1801
rect 34255 1789 34267 1801
rect 34209 1737 34212 1789
rect 34264 1737 34267 1789
rect 34209 1732 34267 1737
rect 34209 1725 34221 1732
rect 34255 1725 34267 1732
rect 34209 1673 34212 1725
rect 34264 1673 34267 1725
rect 34209 1661 34267 1673
rect 34209 1609 34212 1661
rect 34264 1609 34267 1661
rect 34209 1597 34267 1609
rect 34209 1545 34212 1597
rect 34264 1545 34267 1597
rect 34209 1533 34267 1545
rect 34209 1481 34212 1533
rect 34264 1481 34267 1533
rect 34209 1469 34267 1481
rect 34209 1417 34212 1469
rect 34264 1417 34267 1469
rect 34209 1410 34221 1417
rect 34255 1410 34267 1417
rect 34209 1405 34267 1410
rect 34209 1353 34212 1405
rect 34264 1353 34267 1405
rect 34209 1341 34221 1353
rect 34255 1341 34267 1353
rect 34209 1289 34212 1341
rect 34264 1289 34267 1341
rect 34209 1277 34221 1289
rect 34255 1277 34267 1289
rect 34209 1225 34212 1277
rect 34264 1225 34267 1277
rect 34209 1213 34221 1225
rect 34255 1213 34267 1225
rect 34209 1161 34212 1213
rect 34264 1161 34267 1213
rect 34209 1147 34267 1161
rect 34308 3133 34360 3147
rect 34308 3069 34317 3081
rect 34351 3069 34360 3081
rect 34308 3005 34317 3017
rect 34351 3005 34360 3017
rect 34308 2941 34317 2953
rect 34351 2941 34360 2953
rect 34308 2884 34360 2889
rect 34308 2877 34317 2884
rect 34351 2877 34360 2884
rect 34308 2813 34360 2825
rect 34308 2749 34360 2761
rect 34308 2685 34360 2697
rect 34308 2621 34360 2633
rect 34308 2562 34317 2569
rect 34351 2562 34360 2569
rect 34308 2557 34360 2562
rect 34308 2493 34317 2505
rect 34351 2493 34360 2505
rect 34308 2429 34317 2441
rect 34351 2429 34360 2441
rect 34308 2365 34317 2377
rect 34351 2365 34360 2377
rect 34308 2308 34360 2313
rect 34308 2301 34317 2308
rect 34351 2301 34360 2308
rect 34308 2237 34360 2249
rect 34308 2173 34360 2185
rect 34308 2109 34360 2121
rect 34308 2045 34360 2057
rect 34308 1986 34317 1993
rect 34351 1986 34360 1993
rect 34308 1981 34360 1986
rect 34308 1917 34317 1929
rect 34351 1917 34360 1929
rect 34308 1853 34317 1865
rect 34351 1853 34360 1865
rect 34308 1789 34317 1801
rect 34351 1789 34360 1801
rect 34308 1732 34360 1737
rect 34308 1725 34317 1732
rect 34351 1725 34360 1732
rect 34308 1661 34360 1673
rect 34308 1597 34360 1609
rect 34308 1533 34360 1545
rect 34308 1469 34360 1481
rect 34308 1410 34317 1417
rect 34351 1410 34360 1417
rect 34308 1405 34360 1410
rect 34308 1341 34317 1353
rect 34351 1341 34360 1353
rect 34308 1277 34317 1289
rect 34351 1277 34360 1289
rect 34308 1213 34317 1225
rect 34351 1213 34360 1225
rect 34308 1147 34360 1161
rect 34401 3133 34459 3147
rect 34401 3081 34404 3133
rect 34456 3081 34459 3133
rect 34401 3069 34413 3081
rect 34447 3069 34459 3081
rect 34401 3017 34404 3069
rect 34456 3017 34459 3069
rect 34401 3005 34413 3017
rect 34447 3005 34459 3017
rect 34401 2953 34404 3005
rect 34456 2953 34459 3005
rect 34401 2941 34413 2953
rect 34447 2941 34459 2953
rect 34401 2889 34404 2941
rect 34456 2889 34459 2941
rect 34401 2884 34459 2889
rect 34401 2877 34413 2884
rect 34447 2877 34459 2884
rect 34401 2825 34404 2877
rect 34456 2825 34459 2877
rect 34401 2813 34459 2825
rect 34401 2761 34404 2813
rect 34456 2761 34459 2813
rect 34401 2749 34459 2761
rect 34401 2697 34404 2749
rect 34456 2697 34459 2749
rect 34401 2685 34459 2697
rect 34401 2633 34404 2685
rect 34456 2633 34459 2685
rect 34401 2621 34459 2633
rect 34401 2569 34404 2621
rect 34456 2569 34459 2621
rect 34401 2562 34413 2569
rect 34447 2562 34459 2569
rect 34401 2557 34459 2562
rect 34401 2505 34404 2557
rect 34456 2505 34459 2557
rect 34401 2493 34413 2505
rect 34447 2493 34459 2505
rect 34401 2441 34404 2493
rect 34456 2441 34459 2493
rect 34401 2429 34413 2441
rect 34447 2429 34459 2441
rect 34401 2377 34404 2429
rect 34456 2377 34459 2429
rect 34401 2365 34413 2377
rect 34447 2365 34459 2377
rect 34401 2313 34404 2365
rect 34456 2313 34459 2365
rect 34401 2308 34459 2313
rect 34401 2301 34413 2308
rect 34447 2301 34459 2308
rect 34401 2249 34404 2301
rect 34456 2249 34459 2301
rect 34401 2237 34459 2249
rect 34401 2185 34404 2237
rect 34456 2185 34459 2237
rect 34401 2173 34459 2185
rect 34401 2121 34404 2173
rect 34456 2121 34459 2173
rect 34401 2109 34459 2121
rect 34401 2057 34404 2109
rect 34456 2057 34459 2109
rect 34401 2045 34459 2057
rect 34401 1993 34404 2045
rect 34456 1993 34459 2045
rect 34401 1986 34413 1993
rect 34447 1986 34459 1993
rect 34401 1981 34459 1986
rect 34401 1929 34404 1981
rect 34456 1929 34459 1981
rect 34401 1917 34413 1929
rect 34447 1917 34459 1929
rect 34401 1865 34404 1917
rect 34456 1865 34459 1917
rect 34401 1853 34413 1865
rect 34447 1853 34459 1865
rect 34401 1801 34404 1853
rect 34456 1801 34459 1853
rect 34401 1789 34413 1801
rect 34447 1789 34459 1801
rect 34401 1737 34404 1789
rect 34456 1737 34459 1789
rect 34401 1732 34459 1737
rect 34401 1725 34413 1732
rect 34447 1725 34459 1732
rect 34401 1673 34404 1725
rect 34456 1673 34459 1725
rect 34401 1661 34459 1673
rect 34401 1609 34404 1661
rect 34456 1609 34459 1661
rect 34401 1597 34459 1609
rect 34401 1545 34404 1597
rect 34456 1545 34459 1597
rect 34401 1533 34459 1545
rect 34401 1481 34404 1533
rect 34456 1481 34459 1533
rect 34401 1469 34459 1481
rect 34401 1417 34404 1469
rect 34456 1417 34459 1469
rect 34401 1410 34413 1417
rect 34447 1410 34459 1417
rect 34401 1405 34459 1410
rect 34401 1353 34404 1405
rect 34456 1353 34459 1405
rect 34401 1341 34413 1353
rect 34447 1341 34459 1353
rect 34401 1289 34404 1341
rect 34456 1289 34459 1341
rect 34401 1277 34413 1289
rect 34447 1277 34459 1289
rect 34401 1225 34404 1277
rect 34456 1225 34459 1277
rect 34401 1213 34413 1225
rect 34447 1213 34459 1225
rect 34401 1161 34404 1213
rect 34456 1161 34459 1213
rect 34401 1147 34459 1161
rect 34497 3133 34555 3147
rect 34497 3081 34500 3133
rect 34552 3081 34555 3133
rect 34497 3069 34509 3081
rect 34543 3069 34555 3081
rect 34497 3017 34500 3069
rect 34552 3017 34555 3069
rect 34497 3005 34509 3017
rect 34543 3005 34555 3017
rect 34497 2953 34500 3005
rect 34552 2953 34555 3005
rect 34497 2941 34509 2953
rect 34543 2941 34555 2953
rect 34497 2889 34500 2941
rect 34552 2889 34555 2941
rect 34497 2884 34555 2889
rect 34497 2877 34509 2884
rect 34543 2877 34555 2884
rect 34497 2825 34500 2877
rect 34552 2825 34555 2877
rect 34497 2813 34555 2825
rect 34497 2761 34500 2813
rect 34552 2761 34555 2813
rect 34497 2749 34555 2761
rect 34497 2697 34500 2749
rect 34552 2697 34555 2749
rect 34497 2685 34555 2697
rect 34497 2633 34500 2685
rect 34552 2633 34555 2685
rect 34497 2621 34555 2633
rect 34497 2569 34500 2621
rect 34552 2569 34555 2621
rect 34497 2562 34509 2569
rect 34543 2562 34555 2569
rect 34497 2557 34555 2562
rect 34497 2505 34500 2557
rect 34552 2505 34555 2557
rect 34497 2493 34509 2505
rect 34543 2493 34555 2505
rect 34497 2441 34500 2493
rect 34552 2441 34555 2493
rect 34497 2429 34509 2441
rect 34543 2429 34555 2441
rect 34497 2377 34500 2429
rect 34552 2377 34555 2429
rect 34497 2365 34509 2377
rect 34543 2365 34555 2377
rect 34497 2313 34500 2365
rect 34552 2313 34555 2365
rect 34497 2308 34555 2313
rect 34497 2301 34509 2308
rect 34543 2301 34555 2308
rect 34497 2249 34500 2301
rect 34552 2249 34555 2301
rect 34497 2237 34555 2249
rect 34497 2185 34500 2237
rect 34552 2185 34555 2237
rect 34497 2173 34555 2185
rect 34497 2121 34500 2173
rect 34552 2121 34555 2173
rect 34497 2109 34555 2121
rect 34497 2057 34500 2109
rect 34552 2057 34555 2109
rect 34497 2045 34555 2057
rect 34497 1993 34500 2045
rect 34552 1993 34555 2045
rect 34497 1986 34509 1993
rect 34543 1986 34555 1993
rect 34497 1981 34555 1986
rect 34497 1929 34500 1981
rect 34552 1929 34555 1981
rect 34497 1917 34509 1929
rect 34543 1917 34555 1929
rect 34497 1865 34500 1917
rect 34552 1865 34555 1917
rect 34497 1853 34509 1865
rect 34543 1853 34555 1865
rect 34497 1801 34500 1853
rect 34552 1801 34555 1853
rect 34497 1789 34509 1801
rect 34543 1789 34555 1801
rect 34497 1737 34500 1789
rect 34552 1737 34555 1789
rect 34497 1732 34555 1737
rect 34497 1725 34509 1732
rect 34543 1725 34555 1732
rect 34497 1673 34500 1725
rect 34552 1673 34555 1725
rect 34497 1661 34555 1673
rect 34497 1609 34500 1661
rect 34552 1609 34555 1661
rect 34497 1597 34555 1609
rect 34497 1545 34500 1597
rect 34552 1545 34555 1597
rect 34497 1533 34555 1545
rect 34497 1481 34500 1533
rect 34552 1481 34555 1533
rect 34497 1469 34555 1481
rect 34497 1417 34500 1469
rect 34552 1417 34555 1469
rect 34497 1410 34509 1417
rect 34543 1410 34555 1417
rect 34497 1405 34555 1410
rect 34497 1353 34500 1405
rect 34552 1353 34555 1405
rect 34497 1341 34509 1353
rect 34543 1341 34555 1353
rect 34497 1289 34500 1341
rect 34552 1289 34555 1341
rect 34497 1277 34509 1289
rect 34543 1277 34555 1289
rect 34497 1225 34500 1277
rect 34552 1225 34555 1277
rect 34497 1213 34509 1225
rect 34543 1213 34555 1225
rect 34497 1161 34500 1213
rect 34552 1161 34555 1213
rect 34497 1147 34555 1161
rect 34593 3133 34651 3147
rect 34593 3081 34596 3133
rect 34648 3081 34651 3133
rect 34593 3069 34605 3081
rect 34639 3069 34651 3081
rect 34593 3017 34596 3069
rect 34648 3017 34651 3069
rect 34593 3005 34605 3017
rect 34639 3005 34651 3017
rect 34593 2953 34596 3005
rect 34648 2953 34651 3005
rect 34593 2941 34605 2953
rect 34639 2941 34651 2953
rect 34593 2889 34596 2941
rect 34648 2889 34651 2941
rect 34593 2884 34651 2889
rect 34593 2877 34605 2884
rect 34639 2877 34651 2884
rect 34593 2825 34596 2877
rect 34648 2825 34651 2877
rect 34593 2813 34651 2825
rect 34593 2761 34596 2813
rect 34648 2761 34651 2813
rect 34593 2749 34651 2761
rect 34593 2697 34596 2749
rect 34648 2697 34651 2749
rect 34593 2685 34651 2697
rect 34593 2633 34596 2685
rect 34648 2633 34651 2685
rect 34593 2621 34651 2633
rect 34593 2569 34596 2621
rect 34648 2569 34651 2621
rect 34593 2562 34605 2569
rect 34639 2562 34651 2569
rect 34593 2557 34651 2562
rect 34593 2505 34596 2557
rect 34648 2505 34651 2557
rect 34593 2493 34605 2505
rect 34639 2493 34651 2505
rect 34593 2441 34596 2493
rect 34648 2441 34651 2493
rect 34593 2429 34605 2441
rect 34639 2429 34651 2441
rect 34593 2377 34596 2429
rect 34648 2377 34651 2429
rect 34593 2365 34605 2377
rect 34639 2365 34651 2377
rect 34593 2313 34596 2365
rect 34648 2313 34651 2365
rect 34593 2308 34651 2313
rect 34593 2301 34605 2308
rect 34639 2301 34651 2308
rect 34593 2249 34596 2301
rect 34648 2249 34651 2301
rect 34593 2237 34651 2249
rect 34593 2185 34596 2237
rect 34648 2185 34651 2237
rect 34593 2173 34651 2185
rect 34593 2121 34596 2173
rect 34648 2121 34651 2173
rect 34593 2109 34651 2121
rect 34593 2057 34596 2109
rect 34648 2057 34651 2109
rect 34593 2045 34651 2057
rect 34593 1993 34596 2045
rect 34648 1993 34651 2045
rect 34593 1986 34605 1993
rect 34639 1986 34651 1993
rect 34593 1981 34651 1986
rect 34593 1929 34596 1981
rect 34648 1929 34651 1981
rect 34593 1917 34605 1929
rect 34639 1917 34651 1929
rect 34593 1865 34596 1917
rect 34648 1865 34651 1917
rect 34593 1853 34605 1865
rect 34639 1853 34651 1865
rect 34593 1801 34596 1853
rect 34648 1801 34651 1853
rect 34593 1789 34605 1801
rect 34639 1789 34651 1801
rect 34593 1737 34596 1789
rect 34648 1737 34651 1789
rect 34593 1732 34651 1737
rect 34593 1725 34605 1732
rect 34639 1725 34651 1732
rect 34593 1673 34596 1725
rect 34648 1673 34651 1725
rect 34593 1661 34651 1673
rect 34593 1609 34596 1661
rect 34648 1609 34651 1661
rect 34593 1597 34651 1609
rect 34593 1545 34596 1597
rect 34648 1545 34651 1597
rect 34593 1533 34651 1545
rect 34593 1481 34596 1533
rect 34648 1481 34651 1533
rect 34593 1469 34651 1481
rect 34593 1417 34596 1469
rect 34648 1417 34651 1469
rect 34593 1410 34605 1417
rect 34639 1410 34651 1417
rect 34593 1405 34651 1410
rect 34593 1353 34596 1405
rect 34648 1353 34651 1405
rect 34593 1341 34605 1353
rect 34639 1341 34651 1353
rect 34593 1289 34596 1341
rect 34648 1289 34651 1341
rect 34593 1277 34605 1289
rect 34639 1277 34651 1289
rect 34593 1225 34596 1277
rect 34648 1225 34651 1277
rect 34593 1213 34605 1225
rect 34639 1213 34651 1225
rect 34593 1161 34596 1213
rect 34648 1161 34651 1213
rect 34593 1147 34651 1161
rect 34692 3133 34744 3147
rect 34692 3069 34701 3081
rect 34735 3069 34744 3081
rect 34692 3005 34701 3017
rect 34735 3005 34744 3017
rect 34692 2941 34701 2953
rect 34735 2941 34744 2953
rect 34692 2884 34744 2889
rect 34692 2877 34701 2884
rect 34735 2877 34744 2884
rect 34692 2813 34744 2825
rect 34692 2749 34744 2761
rect 34692 2685 34744 2697
rect 34692 2621 34744 2633
rect 34692 2562 34701 2569
rect 34735 2562 34744 2569
rect 34692 2557 34744 2562
rect 34692 2493 34701 2505
rect 34735 2493 34744 2505
rect 34692 2429 34701 2441
rect 34735 2429 34744 2441
rect 34692 2365 34701 2377
rect 34735 2365 34744 2377
rect 34692 2308 34744 2313
rect 34692 2301 34701 2308
rect 34735 2301 34744 2308
rect 34692 2237 34744 2249
rect 34692 2173 34744 2185
rect 34692 2109 34744 2121
rect 34692 2045 34744 2057
rect 34692 1986 34701 1993
rect 34735 1986 34744 1993
rect 34692 1981 34744 1986
rect 34692 1917 34701 1929
rect 34735 1917 34744 1929
rect 34692 1853 34701 1865
rect 34735 1853 34744 1865
rect 34692 1789 34701 1801
rect 34735 1789 34744 1801
rect 34692 1732 34744 1737
rect 34692 1725 34701 1732
rect 34735 1725 34744 1732
rect 34692 1661 34744 1673
rect 34692 1597 34744 1609
rect 34692 1533 34744 1545
rect 34692 1469 34744 1481
rect 34692 1410 34701 1417
rect 34735 1410 34744 1417
rect 34692 1405 34744 1410
rect 34692 1341 34701 1353
rect 34735 1341 34744 1353
rect 34692 1277 34701 1289
rect 34735 1277 34744 1289
rect 34692 1213 34701 1225
rect 34735 1213 34744 1225
rect 34692 1147 34744 1161
rect 34785 3133 34843 3147
rect 34785 3081 34788 3133
rect 34840 3081 34843 3133
rect 34785 3069 34797 3081
rect 34831 3069 34843 3081
rect 34785 3017 34788 3069
rect 34840 3017 34843 3069
rect 34785 3005 34797 3017
rect 34831 3005 34843 3017
rect 34785 2953 34788 3005
rect 34840 2953 34843 3005
rect 34785 2941 34797 2953
rect 34831 2941 34843 2953
rect 34785 2889 34788 2941
rect 34840 2889 34843 2941
rect 34785 2884 34843 2889
rect 34785 2877 34797 2884
rect 34831 2877 34843 2884
rect 34785 2825 34788 2877
rect 34840 2825 34843 2877
rect 34785 2813 34843 2825
rect 34785 2761 34788 2813
rect 34840 2761 34843 2813
rect 34785 2749 34843 2761
rect 34785 2697 34788 2749
rect 34840 2697 34843 2749
rect 34785 2685 34843 2697
rect 34785 2633 34788 2685
rect 34840 2633 34843 2685
rect 34785 2621 34843 2633
rect 34785 2569 34788 2621
rect 34840 2569 34843 2621
rect 34785 2562 34797 2569
rect 34831 2562 34843 2569
rect 34785 2557 34843 2562
rect 34785 2505 34788 2557
rect 34840 2505 34843 2557
rect 34785 2493 34797 2505
rect 34831 2493 34843 2505
rect 34785 2441 34788 2493
rect 34840 2441 34843 2493
rect 34785 2429 34797 2441
rect 34831 2429 34843 2441
rect 34785 2377 34788 2429
rect 34840 2377 34843 2429
rect 34785 2365 34797 2377
rect 34831 2365 34843 2377
rect 34785 2313 34788 2365
rect 34840 2313 34843 2365
rect 34785 2308 34843 2313
rect 34785 2301 34797 2308
rect 34831 2301 34843 2308
rect 34785 2249 34788 2301
rect 34840 2249 34843 2301
rect 34785 2237 34843 2249
rect 34785 2185 34788 2237
rect 34840 2185 34843 2237
rect 34785 2173 34843 2185
rect 34785 2121 34788 2173
rect 34840 2121 34843 2173
rect 34785 2109 34843 2121
rect 34785 2057 34788 2109
rect 34840 2057 34843 2109
rect 34785 2045 34843 2057
rect 34785 1993 34788 2045
rect 34840 1993 34843 2045
rect 34785 1986 34797 1993
rect 34831 1986 34843 1993
rect 34785 1981 34843 1986
rect 34785 1929 34788 1981
rect 34840 1929 34843 1981
rect 34785 1917 34797 1929
rect 34831 1917 34843 1929
rect 34785 1865 34788 1917
rect 34840 1865 34843 1917
rect 34785 1853 34797 1865
rect 34831 1853 34843 1865
rect 34785 1801 34788 1853
rect 34840 1801 34843 1853
rect 34785 1789 34797 1801
rect 34831 1789 34843 1801
rect 34785 1737 34788 1789
rect 34840 1737 34843 1789
rect 34785 1732 34843 1737
rect 34785 1725 34797 1732
rect 34831 1725 34843 1732
rect 34785 1673 34788 1725
rect 34840 1673 34843 1725
rect 34785 1661 34843 1673
rect 34785 1609 34788 1661
rect 34840 1609 34843 1661
rect 34785 1597 34843 1609
rect 34785 1545 34788 1597
rect 34840 1545 34843 1597
rect 34785 1533 34843 1545
rect 34785 1481 34788 1533
rect 34840 1481 34843 1533
rect 34785 1469 34843 1481
rect 34785 1417 34788 1469
rect 34840 1417 34843 1469
rect 34785 1410 34797 1417
rect 34831 1410 34843 1417
rect 34785 1405 34843 1410
rect 34785 1353 34788 1405
rect 34840 1353 34843 1405
rect 34785 1341 34797 1353
rect 34831 1341 34843 1353
rect 34785 1289 34788 1341
rect 34840 1289 34843 1341
rect 34785 1277 34797 1289
rect 34831 1277 34843 1289
rect 34785 1225 34788 1277
rect 34840 1225 34843 1277
rect 34785 1213 34797 1225
rect 34831 1213 34843 1225
rect 34785 1161 34788 1213
rect 34840 1161 34843 1213
rect 34785 1147 34843 1161
rect 34881 3133 34939 3147
rect 34881 3081 34884 3133
rect 34936 3081 34939 3133
rect 34881 3069 34893 3081
rect 34927 3069 34939 3081
rect 34881 3017 34884 3069
rect 34936 3017 34939 3069
rect 34881 3005 34893 3017
rect 34927 3005 34939 3017
rect 34881 2953 34884 3005
rect 34936 2953 34939 3005
rect 34881 2941 34893 2953
rect 34927 2941 34939 2953
rect 34881 2889 34884 2941
rect 34936 2889 34939 2941
rect 34881 2884 34939 2889
rect 34881 2877 34893 2884
rect 34927 2877 34939 2884
rect 34881 2825 34884 2877
rect 34936 2825 34939 2877
rect 34881 2813 34939 2825
rect 34881 2761 34884 2813
rect 34936 2761 34939 2813
rect 34881 2749 34939 2761
rect 34881 2697 34884 2749
rect 34936 2697 34939 2749
rect 34881 2685 34939 2697
rect 34881 2633 34884 2685
rect 34936 2633 34939 2685
rect 34881 2621 34939 2633
rect 34881 2569 34884 2621
rect 34936 2569 34939 2621
rect 34881 2562 34893 2569
rect 34927 2562 34939 2569
rect 34881 2557 34939 2562
rect 34881 2505 34884 2557
rect 34936 2505 34939 2557
rect 34881 2493 34893 2505
rect 34927 2493 34939 2505
rect 34881 2441 34884 2493
rect 34936 2441 34939 2493
rect 34881 2429 34893 2441
rect 34927 2429 34939 2441
rect 34881 2377 34884 2429
rect 34936 2377 34939 2429
rect 34881 2365 34893 2377
rect 34927 2365 34939 2377
rect 34881 2313 34884 2365
rect 34936 2313 34939 2365
rect 34881 2308 34939 2313
rect 34881 2301 34893 2308
rect 34927 2301 34939 2308
rect 34881 2249 34884 2301
rect 34936 2249 34939 2301
rect 34881 2237 34939 2249
rect 34881 2185 34884 2237
rect 34936 2185 34939 2237
rect 34881 2173 34939 2185
rect 34881 2121 34884 2173
rect 34936 2121 34939 2173
rect 34881 2109 34939 2121
rect 34881 2057 34884 2109
rect 34936 2057 34939 2109
rect 34881 2045 34939 2057
rect 34881 1993 34884 2045
rect 34936 1993 34939 2045
rect 34881 1986 34893 1993
rect 34927 1986 34939 1993
rect 34881 1981 34939 1986
rect 34881 1929 34884 1981
rect 34936 1929 34939 1981
rect 34881 1917 34893 1929
rect 34927 1917 34939 1929
rect 34881 1865 34884 1917
rect 34936 1865 34939 1917
rect 34881 1853 34893 1865
rect 34927 1853 34939 1865
rect 34881 1801 34884 1853
rect 34936 1801 34939 1853
rect 34881 1789 34893 1801
rect 34927 1789 34939 1801
rect 34881 1737 34884 1789
rect 34936 1737 34939 1789
rect 34881 1732 34939 1737
rect 34881 1725 34893 1732
rect 34927 1725 34939 1732
rect 34881 1673 34884 1725
rect 34936 1673 34939 1725
rect 34881 1661 34939 1673
rect 34881 1609 34884 1661
rect 34936 1609 34939 1661
rect 34881 1597 34939 1609
rect 34881 1545 34884 1597
rect 34936 1545 34939 1597
rect 34881 1533 34939 1545
rect 34881 1481 34884 1533
rect 34936 1481 34939 1533
rect 34881 1469 34939 1481
rect 34881 1417 34884 1469
rect 34936 1417 34939 1469
rect 34881 1410 34893 1417
rect 34927 1410 34939 1417
rect 34881 1405 34939 1410
rect 34881 1353 34884 1405
rect 34936 1353 34939 1405
rect 34881 1341 34893 1353
rect 34927 1341 34939 1353
rect 34881 1289 34884 1341
rect 34936 1289 34939 1341
rect 34881 1277 34893 1289
rect 34927 1277 34939 1289
rect 34881 1225 34884 1277
rect 34936 1225 34939 1277
rect 34881 1213 34893 1225
rect 34927 1213 34939 1225
rect 34881 1161 34884 1213
rect 34936 1161 34939 1213
rect 34881 1147 34939 1161
rect 34977 3133 35035 3147
rect 34977 3081 34980 3133
rect 35032 3081 35035 3133
rect 34977 3069 34989 3081
rect 35023 3069 35035 3081
rect 34977 3017 34980 3069
rect 35032 3017 35035 3069
rect 34977 3005 34989 3017
rect 35023 3005 35035 3017
rect 34977 2953 34980 3005
rect 35032 2953 35035 3005
rect 34977 2941 34989 2953
rect 35023 2941 35035 2953
rect 34977 2889 34980 2941
rect 35032 2889 35035 2941
rect 34977 2884 35035 2889
rect 34977 2877 34989 2884
rect 35023 2877 35035 2884
rect 34977 2825 34980 2877
rect 35032 2825 35035 2877
rect 34977 2813 35035 2825
rect 34977 2761 34980 2813
rect 35032 2761 35035 2813
rect 34977 2749 35035 2761
rect 34977 2697 34980 2749
rect 35032 2697 35035 2749
rect 34977 2685 35035 2697
rect 34977 2633 34980 2685
rect 35032 2633 35035 2685
rect 34977 2621 35035 2633
rect 34977 2569 34980 2621
rect 35032 2569 35035 2621
rect 34977 2562 34989 2569
rect 35023 2562 35035 2569
rect 34977 2557 35035 2562
rect 34977 2505 34980 2557
rect 35032 2505 35035 2557
rect 34977 2493 34989 2505
rect 35023 2493 35035 2505
rect 34977 2441 34980 2493
rect 35032 2441 35035 2493
rect 34977 2429 34989 2441
rect 35023 2429 35035 2441
rect 34977 2377 34980 2429
rect 35032 2377 35035 2429
rect 34977 2365 34989 2377
rect 35023 2365 35035 2377
rect 34977 2313 34980 2365
rect 35032 2313 35035 2365
rect 34977 2308 35035 2313
rect 34977 2301 34989 2308
rect 35023 2301 35035 2308
rect 34977 2249 34980 2301
rect 35032 2249 35035 2301
rect 34977 2237 35035 2249
rect 34977 2185 34980 2237
rect 35032 2185 35035 2237
rect 34977 2173 35035 2185
rect 34977 2121 34980 2173
rect 35032 2121 35035 2173
rect 34977 2109 35035 2121
rect 34977 2057 34980 2109
rect 35032 2057 35035 2109
rect 34977 2045 35035 2057
rect 34977 1993 34980 2045
rect 35032 1993 35035 2045
rect 34977 1986 34989 1993
rect 35023 1986 35035 1993
rect 34977 1981 35035 1986
rect 34977 1929 34980 1981
rect 35032 1929 35035 1981
rect 34977 1917 34989 1929
rect 35023 1917 35035 1929
rect 34977 1865 34980 1917
rect 35032 1865 35035 1917
rect 34977 1853 34989 1865
rect 35023 1853 35035 1865
rect 34977 1801 34980 1853
rect 35032 1801 35035 1853
rect 34977 1789 34989 1801
rect 35023 1789 35035 1801
rect 34977 1737 34980 1789
rect 35032 1737 35035 1789
rect 34977 1732 35035 1737
rect 34977 1725 34989 1732
rect 35023 1725 35035 1732
rect 34977 1673 34980 1725
rect 35032 1673 35035 1725
rect 34977 1661 35035 1673
rect 34977 1609 34980 1661
rect 35032 1609 35035 1661
rect 34977 1597 35035 1609
rect 34977 1545 34980 1597
rect 35032 1545 35035 1597
rect 34977 1533 35035 1545
rect 34977 1481 34980 1533
rect 35032 1481 35035 1533
rect 34977 1469 35035 1481
rect 34977 1417 34980 1469
rect 35032 1417 35035 1469
rect 34977 1410 34989 1417
rect 35023 1410 35035 1417
rect 34977 1405 35035 1410
rect 34977 1353 34980 1405
rect 35032 1353 35035 1405
rect 34977 1341 34989 1353
rect 35023 1341 35035 1353
rect 34977 1289 34980 1341
rect 35032 1289 35035 1341
rect 34977 1277 34989 1289
rect 35023 1277 35035 1289
rect 34977 1225 34980 1277
rect 35032 1225 35035 1277
rect 34977 1213 34989 1225
rect 35023 1213 35035 1225
rect 34977 1161 34980 1213
rect 35032 1161 35035 1213
rect 34977 1147 35035 1161
rect 35076 3133 35128 3147
rect 35076 3069 35085 3081
rect 35119 3069 35128 3081
rect 35076 3005 35085 3017
rect 35119 3005 35128 3017
rect 35076 2941 35085 2953
rect 35119 2941 35128 2953
rect 35076 2884 35128 2889
rect 35076 2877 35085 2884
rect 35119 2877 35128 2884
rect 35076 2813 35128 2825
rect 35076 2749 35128 2761
rect 35076 2685 35128 2697
rect 35076 2621 35128 2633
rect 35076 2562 35085 2569
rect 35119 2562 35128 2569
rect 35076 2557 35128 2562
rect 35076 2493 35085 2505
rect 35119 2493 35128 2505
rect 35076 2429 35085 2441
rect 35119 2429 35128 2441
rect 35076 2365 35085 2377
rect 35119 2365 35128 2377
rect 35076 2308 35128 2313
rect 35076 2301 35085 2308
rect 35119 2301 35128 2308
rect 35076 2237 35128 2249
rect 35076 2173 35128 2185
rect 35076 2109 35128 2121
rect 35076 2045 35128 2057
rect 35076 1986 35085 1993
rect 35119 1986 35128 1993
rect 35076 1981 35128 1986
rect 35076 1917 35085 1929
rect 35119 1917 35128 1929
rect 35076 1853 35085 1865
rect 35119 1853 35128 1865
rect 35076 1789 35085 1801
rect 35119 1789 35128 1801
rect 35076 1732 35128 1737
rect 35076 1725 35085 1732
rect 35119 1725 35128 1732
rect 35076 1661 35128 1673
rect 35076 1597 35128 1609
rect 35076 1533 35128 1545
rect 35076 1469 35128 1481
rect 35076 1410 35085 1417
rect 35119 1410 35128 1417
rect 35076 1405 35128 1410
rect 35076 1341 35085 1353
rect 35119 1341 35128 1353
rect 35076 1277 35085 1289
rect 35119 1277 35128 1289
rect 35076 1213 35085 1225
rect 35119 1213 35128 1225
rect 35076 1147 35128 1161
rect 35169 3133 35227 3147
rect 35169 3081 35172 3133
rect 35224 3081 35227 3133
rect 35169 3069 35181 3081
rect 35215 3069 35227 3081
rect 35169 3017 35172 3069
rect 35224 3017 35227 3069
rect 35169 3005 35181 3017
rect 35215 3005 35227 3017
rect 35169 2953 35172 3005
rect 35224 2953 35227 3005
rect 35169 2941 35181 2953
rect 35215 2941 35227 2953
rect 35169 2889 35172 2941
rect 35224 2889 35227 2941
rect 35169 2884 35227 2889
rect 35169 2877 35181 2884
rect 35215 2877 35227 2884
rect 35169 2825 35172 2877
rect 35224 2825 35227 2877
rect 35169 2813 35227 2825
rect 35169 2761 35172 2813
rect 35224 2761 35227 2813
rect 35169 2749 35227 2761
rect 35169 2697 35172 2749
rect 35224 2697 35227 2749
rect 35169 2685 35227 2697
rect 35169 2633 35172 2685
rect 35224 2633 35227 2685
rect 35169 2621 35227 2633
rect 35169 2569 35172 2621
rect 35224 2569 35227 2621
rect 35169 2562 35181 2569
rect 35215 2562 35227 2569
rect 35169 2557 35227 2562
rect 35169 2505 35172 2557
rect 35224 2505 35227 2557
rect 35169 2493 35181 2505
rect 35215 2493 35227 2505
rect 35169 2441 35172 2493
rect 35224 2441 35227 2493
rect 35169 2429 35181 2441
rect 35215 2429 35227 2441
rect 35169 2377 35172 2429
rect 35224 2377 35227 2429
rect 35169 2365 35181 2377
rect 35215 2365 35227 2377
rect 35169 2313 35172 2365
rect 35224 2313 35227 2365
rect 35169 2308 35227 2313
rect 35169 2301 35181 2308
rect 35215 2301 35227 2308
rect 35169 2249 35172 2301
rect 35224 2249 35227 2301
rect 35169 2237 35227 2249
rect 35169 2185 35172 2237
rect 35224 2185 35227 2237
rect 35169 2173 35227 2185
rect 35169 2121 35172 2173
rect 35224 2121 35227 2173
rect 35169 2109 35227 2121
rect 35169 2057 35172 2109
rect 35224 2057 35227 2109
rect 35169 2045 35227 2057
rect 35169 1993 35172 2045
rect 35224 1993 35227 2045
rect 35169 1986 35181 1993
rect 35215 1986 35227 1993
rect 35169 1981 35227 1986
rect 35169 1929 35172 1981
rect 35224 1929 35227 1981
rect 35169 1917 35181 1929
rect 35215 1917 35227 1929
rect 35169 1865 35172 1917
rect 35224 1865 35227 1917
rect 35169 1853 35181 1865
rect 35215 1853 35227 1865
rect 35169 1801 35172 1853
rect 35224 1801 35227 1853
rect 35169 1789 35181 1801
rect 35215 1789 35227 1801
rect 35169 1737 35172 1789
rect 35224 1737 35227 1789
rect 35169 1732 35227 1737
rect 35169 1725 35181 1732
rect 35215 1725 35227 1732
rect 35169 1673 35172 1725
rect 35224 1673 35227 1725
rect 35169 1661 35227 1673
rect 35169 1609 35172 1661
rect 35224 1609 35227 1661
rect 35169 1597 35227 1609
rect 35169 1545 35172 1597
rect 35224 1545 35227 1597
rect 35169 1533 35227 1545
rect 35169 1481 35172 1533
rect 35224 1481 35227 1533
rect 35169 1469 35227 1481
rect 35169 1417 35172 1469
rect 35224 1417 35227 1469
rect 35169 1410 35181 1417
rect 35215 1410 35227 1417
rect 35169 1405 35227 1410
rect 35169 1353 35172 1405
rect 35224 1353 35227 1405
rect 35169 1341 35181 1353
rect 35215 1341 35227 1353
rect 35169 1289 35172 1341
rect 35224 1289 35227 1341
rect 35169 1277 35181 1289
rect 35215 1277 35227 1289
rect 35169 1225 35172 1277
rect 35224 1225 35227 1277
rect 35169 1213 35181 1225
rect 35215 1213 35227 1225
rect 35169 1161 35172 1213
rect 35224 1161 35227 1213
rect 35169 1147 35227 1161
rect 35265 3133 35323 3147
rect 35265 3081 35268 3133
rect 35320 3081 35323 3133
rect 35265 3069 35277 3081
rect 35311 3069 35323 3081
rect 35265 3017 35268 3069
rect 35320 3017 35323 3069
rect 35265 3005 35277 3017
rect 35311 3005 35323 3017
rect 35265 2953 35268 3005
rect 35320 2953 35323 3005
rect 35265 2941 35277 2953
rect 35311 2941 35323 2953
rect 35265 2889 35268 2941
rect 35320 2889 35323 2941
rect 35265 2884 35323 2889
rect 35265 2877 35277 2884
rect 35311 2877 35323 2884
rect 35265 2825 35268 2877
rect 35320 2825 35323 2877
rect 35265 2813 35323 2825
rect 35265 2761 35268 2813
rect 35320 2761 35323 2813
rect 35265 2749 35323 2761
rect 35265 2697 35268 2749
rect 35320 2697 35323 2749
rect 35265 2685 35323 2697
rect 35265 2633 35268 2685
rect 35320 2633 35323 2685
rect 35265 2621 35323 2633
rect 35265 2569 35268 2621
rect 35320 2569 35323 2621
rect 35265 2562 35277 2569
rect 35311 2562 35323 2569
rect 35265 2557 35323 2562
rect 35265 2505 35268 2557
rect 35320 2505 35323 2557
rect 35265 2493 35277 2505
rect 35311 2493 35323 2505
rect 35265 2441 35268 2493
rect 35320 2441 35323 2493
rect 35265 2429 35277 2441
rect 35311 2429 35323 2441
rect 35265 2377 35268 2429
rect 35320 2377 35323 2429
rect 35265 2365 35277 2377
rect 35311 2365 35323 2377
rect 35265 2313 35268 2365
rect 35320 2313 35323 2365
rect 35265 2308 35323 2313
rect 35265 2301 35277 2308
rect 35311 2301 35323 2308
rect 35265 2249 35268 2301
rect 35320 2249 35323 2301
rect 35265 2237 35323 2249
rect 35265 2185 35268 2237
rect 35320 2185 35323 2237
rect 35265 2173 35323 2185
rect 35265 2121 35268 2173
rect 35320 2121 35323 2173
rect 35265 2109 35323 2121
rect 35265 2057 35268 2109
rect 35320 2057 35323 2109
rect 35265 2045 35323 2057
rect 35265 1993 35268 2045
rect 35320 1993 35323 2045
rect 35265 1986 35277 1993
rect 35311 1986 35323 1993
rect 35265 1981 35323 1986
rect 35265 1929 35268 1981
rect 35320 1929 35323 1981
rect 35265 1917 35277 1929
rect 35311 1917 35323 1929
rect 35265 1865 35268 1917
rect 35320 1865 35323 1917
rect 35265 1853 35277 1865
rect 35311 1853 35323 1865
rect 35265 1801 35268 1853
rect 35320 1801 35323 1853
rect 35265 1789 35277 1801
rect 35311 1789 35323 1801
rect 35265 1737 35268 1789
rect 35320 1737 35323 1789
rect 35265 1732 35323 1737
rect 35265 1725 35277 1732
rect 35311 1725 35323 1732
rect 35265 1673 35268 1725
rect 35320 1673 35323 1725
rect 35265 1661 35323 1673
rect 35265 1609 35268 1661
rect 35320 1609 35323 1661
rect 35265 1597 35323 1609
rect 35265 1545 35268 1597
rect 35320 1545 35323 1597
rect 35265 1533 35323 1545
rect 35265 1481 35268 1533
rect 35320 1481 35323 1533
rect 35265 1469 35323 1481
rect 35265 1417 35268 1469
rect 35320 1417 35323 1469
rect 35265 1410 35277 1417
rect 35311 1410 35323 1417
rect 35265 1405 35323 1410
rect 35265 1353 35268 1405
rect 35320 1353 35323 1405
rect 35265 1341 35277 1353
rect 35311 1341 35323 1353
rect 35265 1289 35268 1341
rect 35320 1289 35323 1341
rect 35265 1277 35277 1289
rect 35311 1277 35323 1289
rect 35265 1225 35268 1277
rect 35320 1225 35323 1277
rect 35265 1213 35277 1225
rect 35311 1213 35323 1225
rect 35265 1161 35268 1213
rect 35320 1161 35323 1213
rect 35265 1147 35323 1161
rect 35361 3133 35419 3147
rect 35361 3081 35364 3133
rect 35416 3081 35419 3133
rect 35361 3069 35373 3081
rect 35407 3069 35419 3081
rect 35361 3017 35364 3069
rect 35416 3017 35419 3069
rect 35361 3005 35373 3017
rect 35407 3005 35419 3017
rect 35361 2953 35364 3005
rect 35416 2953 35419 3005
rect 35361 2941 35373 2953
rect 35407 2941 35419 2953
rect 35361 2889 35364 2941
rect 35416 2889 35419 2941
rect 35361 2884 35419 2889
rect 35361 2877 35373 2884
rect 35407 2877 35419 2884
rect 35361 2825 35364 2877
rect 35416 2825 35419 2877
rect 35361 2813 35419 2825
rect 35361 2761 35364 2813
rect 35416 2761 35419 2813
rect 35361 2749 35419 2761
rect 35361 2697 35364 2749
rect 35416 2697 35419 2749
rect 35361 2685 35419 2697
rect 35361 2633 35364 2685
rect 35416 2633 35419 2685
rect 35361 2621 35419 2633
rect 35361 2569 35364 2621
rect 35416 2569 35419 2621
rect 35361 2562 35373 2569
rect 35407 2562 35419 2569
rect 35361 2557 35419 2562
rect 35361 2505 35364 2557
rect 35416 2505 35419 2557
rect 35361 2493 35373 2505
rect 35407 2493 35419 2505
rect 35361 2441 35364 2493
rect 35416 2441 35419 2493
rect 35361 2429 35373 2441
rect 35407 2429 35419 2441
rect 35361 2377 35364 2429
rect 35416 2377 35419 2429
rect 35361 2365 35373 2377
rect 35407 2365 35419 2377
rect 35361 2313 35364 2365
rect 35416 2313 35419 2365
rect 35361 2308 35419 2313
rect 35361 2301 35373 2308
rect 35407 2301 35419 2308
rect 35361 2249 35364 2301
rect 35416 2249 35419 2301
rect 35361 2237 35419 2249
rect 35361 2185 35364 2237
rect 35416 2185 35419 2237
rect 35361 2173 35419 2185
rect 35361 2121 35364 2173
rect 35416 2121 35419 2173
rect 35361 2109 35419 2121
rect 35361 2057 35364 2109
rect 35416 2057 35419 2109
rect 35361 2045 35419 2057
rect 35361 1993 35364 2045
rect 35416 1993 35419 2045
rect 35361 1986 35373 1993
rect 35407 1986 35419 1993
rect 35361 1981 35419 1986
rect 35361 1929 35364 1981
rect 35416 1929 35419 1981
rect 35361 1917 35373 1929
rect 35407 1917 35419 1929
rect 35361 1865 35364 1917
rect 35416 1865 35419 1917
rect 35361 1853 35373 1865
rect 35407 1853 35419 1865
rect 35361 1801 35364 1853
rect 35416 1801 35419 1853
rect 35361 1789 35373 1801
rect 35407 1789 35419 1801
rect 35361 1737 35364 1789
rect 35416 1737 35419 1789
rect 35361 1732 35419 1737
rect 35361 1725 35373 1732
rect 35407 1725 35419 1732
rect 35361 1673 35364 1725
rect 35416 1673 35419 1725
rect 35361 1661 35419 1673
rect 35361 1609 35364 1661
rect 35416 1609 35419 1661
rect 35361 1597 35419 1609
rect 35361 1545 35364 1597
rect 35416 1545 35419 1597
rect 35361 1533 35419 1545
rect 35361 1481 35364 1533
rect 35416 1481 35419 1533
rect 35361 1469 35419 1481
rect 35361 1417 35364 1469
rect 35416 1417 35419 1469
rect 35361 1410 35373 1417
rect 35407 1410 35419 1417
rect 35361 1405 35419 1410
rect 35361 1353 35364 1405
rect 35416 1353 35419 1405
rect 35361 1341 35373 1353
rect 35407 1341 35419 1353
rect 35361 1289 35364 1341
rect 35416 1289 35419 1341
rect 35361 1277 35373 1289
rect 35407 1277 35419 1289
rect 35361 1225 35364 1277
rect 35416 1225 35419 1277
rect 35361 1213 35373 1225
rect 35407 1213 35419 1225
rect 35361 1161 35364 1213
rect 35416 1161 35419 1213
rect 35361 1147 35419 1161
rect 35460 3133 35512 3147
rect 35460 3069 35469 3081
rect 35503 3069 35512 3081
rect 35460 3005 35469 3017
rect 35503 3005 35512 3017
rect 35460 2941 35469 2953
rect 35503 2941 35512 2953
rect 35460 2884 35512 2889
rect 35460 2877 35469 2884
rect 35503 2877 35512 2884
rect 35460 2813 35512 2825
rect 35460 2749 35512 2761
rect 35460 2685 35512 2697
rect 35460 2621 35512 2633
rect 35460 2562 35469 2569
rect 35503 2562 35512 2569
rect 35460 2557 35512 2562
rect 35460 2493 35469 2505
rect 35503 2493 35512 2505
rect 35460 2429 35469 2441
rect 35503 2429 35512 2441
rect 35460 2365 35469 2377
rect 35503 2365 35512 2377
rect 35460 2308 35512 2313
rect 35460 2301 35469 2308
rect 35503 2301 35512 2308
rect 35460 2237 35512 2249
rect 35460 2173 35512 2185
rect 35460 2109 35512 2121
rect 35460 2045 35512 2057
rect 35460 1986 35469 1993
rect 35503 1986 35512 1993
rect 35460 1981 35512 1986
rect 35460 1917 35469 1929
rect 35503 1917 35512 1929
rect 35460 1853 35469 1865
rect 35503 1853 35512 1865
rect 35460 1789 35469 1801
rect 35503 1789 35512 1801
rect 35460 1732 35512 1737
rect 35460 1725 35469 1732
rect 35503 1725 35512 1732
rect 35460 1661 35512 1673
rect 35460 1597 35512 1609
rect 35460 1533 35512 1545
rect 35460 1469 35512 1481
rect 35460 1410 35469 1417
rect 35503 1410 35512 1417
rect 35460 1405 35512 1410
rect 35460 1341 35469 1353
rect 35503 1341 35512 1353
rect 35460 1277 35469 1289
rect 35503 1277 35512 1289
rect 35460 1213 35469 1225
rect 35503 1213 35512 1225
rect 35460 1147 35512 1161
rect 35553 3133 35611 3147
rect 35553 3081 35556 3133
rect 35608 3081 35611 3133
rect 35553 3069 35565 3081
rect 35599 3069 35611 3081
rect 35553 3017 35556 3069
rect 35608 3017 35611 3069
rect 35553 3005 35565 3017
rect 35599 3005 35611 3017
rect 35553 2953 35556 3005
rect 35608 2953 35611 3005
rect 35553 2941 35565 2953
rect 35599 2941 35611 2953
rect 35553 2889 35556 2941
rect 35608 2889 35611 2941
rect 35553 2884 35611 2889
rect 35553 2877 35565 2884
rect 35599 2877 35611 2884
rect 35553 2825 35556 2877
rect 35608 2825 35611 2877
rect 35553 2813 35611 2825
rect 35553 2761 35556 2813
rect 35608 2761 35611 2813
rect 35553 2749 35611 2761
rect 35553 2697 35556 2749
rect 35608 2697 35611 2749
rect 35553 2685 35611 2697
rect 35553 2633 35556 2685
rect 35608 2633 35611 2685
rect 35553 2621 35611 2633
rect 35553 2569 35556 2621
rect 35608 2569 35611 2621
rect 35553 2562 35565 2569
rect 35599 2562 35611 2569
rect 35553 2557 35611 2562
rect 35553 2505 35556 2557
rect 35608 2505 35611 2557
rect 35553 2493 35565 2505
rect 35599 2493 35611 2505
rect 35553 2441 35556 2493
rect 35608 2441 35611 2493
rect 35553 2429 35565 2441
rect 35599 2429 35611 2441
rect 35553 2377 35556 2429
rect 35608 2377 35611 2429
rect 35553 2365 35565 2377
rect 35599 2365 35611 2377
rect 35553 2313 35556 2365
rect 35608 2313 35611 2365
rect 35553 2308 35611 2313
rect 35553 2301 35565 2308
rect 35599 2301 35611 2308
rect 35553 2249 35556 2301
rect 35608 2249 35611 2301
rect 35553 2237 35611 2249
rect 35553 2185 35556 2237
rect 35608 2185 35611 2237
rect 35553 2173 35611 2185
rect 35553 2121 35556 2173
rect 35608 2121 35611 2173
rect 35553 2109 35611 2121
rect 35553 2057 35556 2109
rect 35608 2057 35611 2109
rect 35553 2045 35611 2057
rect 35553 1993 35556 2045
rect 35608 1993 35611 2045
rect 35553 1986 35565 1993
rect 35599 1986 35611 1993
rect 35553 1981 35611 1986
rect 35553 1929 35556 1981
rect 35608 1929 35611 1981
rect 35553 1917 35565 1929
rect 35599 1917 35611 1929
rect 35553 1865 35556 1917
rect 35608 1865 35611 1917
rect 35553 1853 35565 1865
rect 35599 1853 35611 1865
rect 35553 1801 35556 1853
rect 35608 1801 35611 1853
rect 35553 1789 35565 1801
rect 35599 1789 35611 1801
rect 35553 1737 35556 1789
rect 35608 1737 35611 1789
rect 35553 1732 35611 1737
rect 35553 1725 35565 1732
rect 35599 1725 35611 1732
rect 35553 1673 35556 1725
rect 35608 1673 35611 1725
rect 35553 1661 35611 1673
rect 35553 1609 35556 1661
rect 35608 1609 35611 1661
rect 35553 1597 35611 1609
rect 35553 1545 35556 1597
rect 35608 1545 35611 1597
rect 35553 1533 35611 1545
rect 35553 1481 35556 1533
rect 35608 1481 35611 1533
rect 35553 1469 35611 1481
rect 35553 1417 35556 1469
rect 35608 1417 35611 1469
rect 35553 1410 35565 1417
rect 35599 1410 35611 1417
rect 35553 1405 35611 1410
rect 35553 1353 35556 1405
rect 35608 1353 35611 1405
rect 35553 1341 35565 1353
rect 35599 1341 35611 1353
rect 35553 1289 35556 1341
rect 35608 1289 35611 1341
rect 35553 1277 35565 1289
rect 35599 1277 35611 1289
rect 35553 1225 35556 1277
rect 35608 1225 35611 1277
rect 35553 1213 35565 1225
rect 35599 1213 35611 1225
rect 35553 1161 35556 1213
rect 35608 1161 35611 1213
rect 35553 1147 35611 1161
rect 35649 3133 35707 3147
rect 35649 3081 35652 3133
rect 35704 3081 35707 3133
rect 35649 3069 35661 3081
rect 35695 3069 35707 3081
rect 35649 3017 35652 3069
rect 35704 3017 35707 3069
rect 35649 3005 35661 3017
rect 35695 3005 35707 3017
rect 35649 2953 35652 3005
rect 35704 2953 35707 3005
rect 35649 2941 35661 2953
rect 35695 2941 35707 2953
rect 35649 2889 35652 2941
rect 35704 2889 35707 2941
rect 35649 2884 35707 2889
rect 35649 2877 35661 2884
rect 35695 2877 35707 2884
rect 35649 2825 35652 2877
rect 35704 2825 35707 2877
rect 35649 2813 35707 2825
rect 35649 2761 35652 2813
rect 35704 2761 35707 2813
rect 35649 2749 35707 2761
rect 35649 2697 35652 2749
rect 35704 2697 35707 2749
rect 35649 2685 35707 2697
rect 35649 2633 35652 2685
rect 35704 2633 35707 2685
rect 35649 2621 35707 2633
rect 35649 2569 35652 2621
rect 35704 2569 35707 2621
rect 35649 2562 35661 2569
rect 35695 2562 35707 2569
rect 35649 2557 35707 2562
rect 35649 2505 35652 2557
rect 35704 2505 35707 2557
rect 35649 2493 35661 2505
rect 35695 2493 35707 2505
rect 35649 2441 35652 2493
rect 35704 2441 35707 2493
rect 35649 2429 35661 2441
rect 35695 2429 35707 2441
rect 35649 2377 35652 2429
rect 35704 2377 35707 2429
rect 35649 2365 35661 2377
rect 35695 2365 35707 2377
rect 35649 2313 35652 2365
rect 35704 2313 35707 2365
rect 35649 2308 35707 2313
rect 35649 2301 35661 2308
rect 35695 2301 35707 2308
rect 35649 2249 35652 2301
rect 35704 2249 35707 2301
rect 35649 2237 35707 2249
rect 35649 2185 35652 2237
rect 35704 2185 35707 2237
rect 35649 2173 35707 2185
rect 35649 2121 35652 2173
rect 35704 2121 35707 2173
rect 35649 2109 35707 2121
rect 35649 2057 35652 2109
rect 35704 2057 35707 2109
rect 35649 2045 35707 2057
rect 35649 1993 35652 2045
rect 35704 1993 35707 2045
rect 35649 1986 35661 1993
rect 35695 1986 35707 1993
rect 35649 1981 35707 1986
rect 35649 1929 35652 1981
rect 35704 1929 35707 1981
rect 35649 1917 35661 1929
rect 35695 1917 35707 1929
rect 35649 1865 35652 1917
rect 35704 1865 35707 1917
rect 35649 1853 35661 1865
rect 35695 1853 35707 1865
rect 35649 1801 35652 1853
rect 35704 1801 35707 1853
rect 35649 1789 35661 1801
rect 35695 1789 35707 1801
rect 35649 1737 35652 1789
rect 35704 1737 35707 1789
rect 35649 1732 35707 1737
rect 35649 1725 35661 1732
rect 35695 1725 35707 1732
rect 35649 1673 35652 1725
rect 35704 1673 35707 1725
rect 35649 1661 35707 1673
rect 35649 1609 35652 1661
rect 35704 1609 35707 1661
rect 35649 1597 35707 1609
rect 35649 1545 35652 1597
rect 35704 1545 35707 1597
rect 35649 1533 35707 1545
rect 35649 1481 35652 1533
rect 35704 1481 35707 1533
rect 35649 1469 35707 1481
rect 35649 1417 35652 1469
rect 35704 1417 35707 1469
rect 35649 1410 35661 1417
rect 35695 1410 35707 1417
rect 35649 1405 35707 1410
rect 35649 1353 35652 1405
rect 35704 1353 35707 1405
rect 35649 1341 35661 1353
rect 35695 1341 35707 1353
rect 35649 1289 35652 1341
rect 35704 1289 35707 1341
rect 35649 1277 35661 1289
rect 35695 1277 35707 1289
rect 35649 1225 35652 1277
rect 35704 1225 35707 1277
rect 35649 1213 35661 1225
rect 35695 1213 35707 1225
rect 35649 1161 35652 1213
rect 35704 1161 35707 1213
rect 35649 1147 35707 1161
rect 35745 3133 35803 3147
rect 35745 3081 35748 3133
rect 35800 3081 35803 3133
rect 35745 3069 35757 3081
rect 35791 3069 35803 3081
rect 35745 3017 35748 3069
rect 35800 3017 35803 3069
rect 35745 3005 35757 3017
rect 35791 3005 35803 3017
rect 35745 2953 35748 3005
rect 35800 2953 35803 3005
rect 35745 2941 35757 2953
rect 35791 2941 35803 2953
rect 35745 2889 35748 2941
rect 35800 2889 35803 2941
rect 35745 2884 35803 2889
rect 35745 2877 35757 2884
rect 35791 2877 35803 2884
rect 35745 2825 35748 2877
rect 35800 2825 35803 2877
rect 35745 2813 35803 2825
rect 35745 2761 35748 2813
rect 35800 2761 35803 2813
rect 35745 2749 35803 2761
rect 35745 2697 35748 2749
rect 35800 2697 35803 2749
rect 35745 2685 35803 2697
rect 35745 2633 35748 2685
rect 35800 2633 35803 2685
rect 35745 2621 35803 2633
rect 35745 2569 35748 2621
rect 35800 2569 35803 2621
rect 35745 2562 35757 2569
rect 35791 2562 35803 2569
rect 35745 2557 35803 2562
rect 35745 2505 35748 2557
rect 35800 2505 35803 2557
rect 35745 2493 35757 2505
rect 35791 2493 35803 2505
rect 35745 2441 35748 2493
rect 35800 2441 35803 2493
rect 35745 2429 35757 2441
rect 35791 2429 35803 2441
rect 35745 2377 35748 2429
rect 35800 2377 35803 2429
rect 35745 2365 35757 2377
rect 35791 2365 35803 2377
rect 35745 2313 35748 2365
rect 35800 2313 35803 2365
rect 35745 2308 35803 2313
rect 35745 2301 35757 2308
rect 35791 2301 35803 2308
rect 35745 2249 35748 2301
rect 35800 2249 35803 2301
rect 35745 2237 35803 2249
rect 35745 2185 35748 2237
rect 35800 2185 35803 2237
rect 35745 2173 35803 2185
rect 35745 2121 35748 2173
rect 35800 2121 35803 2173
rect 35745 2109 35803 2121
rect 35745 2057 35748 2109
rect 35800 2057 35803 2109
rect 35745 2045 35803 2057
rect 35745 1993 35748 2045
rect 35800 1993 35803 2045
rect 35745 1986 35757 1993
rect 35791 1986 35803 1993
rect 35745 1981 35803 1986
rect 35745 1929 35748 1981
rect 35800 1929 35803 1981
rect 35745 1917 35757 1929
rect 35791 1917 35803 1929
rect 35745 1865 35748 1917
rect 35800 1865 35803 1917
rect 35745 1853 35757 1865
rect 35791 1853 35803 1865
rect 35745 1801 35748 1853
rect 35800 1801 35803 1853
rect 35745 1789 35757 1801
rect 35791 1789 35803 1801
rect 35745 1737 35748 1789
rect 35800 1737 35803 1789
rect 35745 1732 35803 1737
rect 35745 1725 35757 1732
rect 35791 1725 35803 1732
rect 35745 1673 35748 1725
rect 35800 1673 35803 1725
rect 35745 1661 35803 1673
rect 35745 1609 35748 1661
rect 35800 1609 35803 1661
rect 35745 1597 35803 1609
rect 35745 1545 35748 1597
rect 35800 1545 35803 1597
rect 35745 1533 35803 1545
rect 35745 1481 35748 1533
rect 35800 1481 35803 1533
rect 35745 1469 35803 1481
rect 35745 1417 35748 1469
rect 35800 1417 35803 1469
rect 35745 1410 35757 1417
rect 35791 1410 35803 1417
rect 35745 1405 35803 1410
rect 35745 1353 35748 1405
rect 35800 1353 35803 1405
rect 35745 1341 35757 1353
rect 35791 1341 35803 1353
rect 35745 1289 35748 1341
rect 35800 1289 35803 1341
rect 35745 1277 35757 1289
rect 35791 1277 35803 1289
rect 35745 1225 35748 1277
rect 35800 1225 35803 1277
rect 35745 1213 35757 1225
rect 35791 1213 35803 1225
rect 35745 1161 35748 1213
rect 35800 1161 35803 1213
rect 35745 1147 35803 1161
rect 35844 3133 35896 3147
rect 35844 3069 35853 3081
rect 35887 3069 35896 3081
rect 35844 3005 35853 3017
rect 35887 3005 35896 3017
rect 35844 2941 35853 2953
rect 35887 2941 35896 2953
rect 35844 2884 35896 2889
rect 35844 2877 35853 2884
rect 35887 2877 35896 2884
rect 35844 2813 35896 2825
rect 35844 2749 35896 2761
rect 35844 2685 35896 2697
rect 35844 2621 35896 2633
rect 35844 2562 35853 2569
rect 35887 2562 35896 2569
rect 35844 2557 35896 2562
rect 35844 2493 35853 2505
rect 35887 2493 35896 2505
rect 35844 2429 35853 2441
rect 35887 2429 35896 2441
rect 35844 2365 35853 2377
rect 35887 2365 35896 2377
rect 35844 2308 35896 2313
rect 35844 2301 35853 2308
rect 35887 2301 35896 2308
rect 35844 2237 35896 2249
rect 35844 2173 35896 2185
rect 35844 2109 35896 2121
rect 35844 2045 35896 2057
rect 35844 1986 35853 1993
rect 35887 1986 35896 1993
rect 35844 1981 35896 1986
rect 35844 1917 35853 1929
rect 35887 1917 35896 1929
rect 35844 1853 35853 1865
rect 35887 1853 35896 1865
rect 35844 1789 35853 1801
rect 35887 1789 35896 1801
rect 35844 1732 35896 1737
rect 35844 1725 35853 1732
rect 35887 1725 35896 1732
rect 35844 1661 35896 1673
rect 35844 1597 35896 1609
rect 35844 1533 35896 1545
rect 35844 1469 35896 1481
rect 35844 1410 35853 1417
rect 35887 1410 35896 1417
rect 35844 1405 35896 1410
rect 35844 1341 35853 1353
rect 35887 1341 35896 1353
rect 35844 1277 35853 1289
rect 35887 1277 35896 1289
rect 35844 1213 35853 1225
rect 35887 1213 35896 1225
rect 35844 1147 35896 1161
rect 35937 3133 35995 3147
rect 35937 3081 35940 3133
rect 35992 3081 35995 3133
rect 35937 3069 35949 3081
rect 35983 3069 35995 3081
rect 35937 3017 35940 3069
rect 35992 3017 35995 3069
rect 35937 3005 35949 3017
rect 35983 3005 35995 3017
rect 35937 2953 35940 3005
rect 35992 2953 35995 3005
rect 35937 2941 35949 2953
rect 35983 2941 35995 2953
rect 35937 2889 35940 2941
rect 35992 2889 35995 2941
rect 35937 2884 35995 2889
rect 35937 2877 35949 2884
rect 35983 2877 35995 2884
rect 35937 2825 35940 2877
rect 35992 2825 35995 2877
rect 35937 2813 35995 2825
rect 35937 2761 35940 2813
rect 35992 2761 35995 2813
rect 35937 2749 35995 2761
rect 35937 2697 35940 2749
rect 35992 2697 35995 2749
rect 35937 2685 35995 2697
rect 35937 2633 35940 2685
rect 35992 2633 35995 2685
rect 35937 2621 35995 2633
rect 35937 2569 35940 2621
rect 35992 2569 35995 2621
rect 35937 2562 35949 2569
rect 35983 2562 35995 2569
rect 35937 2557 35995 2562
rect 35937 2505 35940 2557
rect 35992 2505 35995 2557
rect 35937 2493 35949 2505
rect 35983 2493 35995 2505
rect 35937 2441 35940 2493
rect 35992 2441 35995 2493
rect 35937 2429 35949 2441
rect 35983 2429 35995 2441
rect 35937 2377 35940 2429
rect 35992 2377 35995 2429
rect 35937 2365 35949 2377
rect 35983 2365 35995 2377
rect 35937 2313 35940 2365
rect 35992 2313 35995 2365
rect 35937 2308 35995 2313
rect 35937 2301 35949 2308
rect 35983 2301 35995 2308
rect 35937 2249 35940 2301
rect 35992 2249 35995 2301
rect 35937 2237 35995 2249
rect 35937 2185 35940 2237
rect 35992 2185 35995 2237
rect 35937 2173 35995 2185
rect 35937 2121 35940 2173
rect 35992 2121 35995 2173
rect 35937 2109 35995 2121
rect 35937 2057 35940 2109
rect 35992 2057 35995 2109
rect 35937 2045 35995 2057
rect 35937 1993 35940 2045
rect 35992 1993 35995 2045
rect 35937 1986 35949 1993
rect 35983 1986 35995 1993
rect 35937 1981 35995 1986
rect 35937 1929 35940 1981
rect 35992 1929 35995 1981
rect 35937 1917 35949 1929
rect 35983 1917 35995 1929
rect 35937 1865 35940 1917
rect 35992 1865 35995 1917
rect 35937 1853 35949 1865
rect 35983 1853 35995 1865
rect 35937 1801 35940 1853
rect 35992 1801 35995 1853
rect 35937 1789 35949 1801
rect 35983 1789 35995 1801
rect 35937 1737 35940 1789
rect 35992 1737 35995 1789
rect 35937 1732 35995 1737
rect 35937 1725 35949 1732
rect 35983 1725 35995 1732
rect 35937 1673 35940 1725
rect 35992 1673 35995 1725
rect 35937 1661 35995 1673
rect 35937 1609 35940 1661
rect 35992 1609 35995 1661
rect 35937 1597 35995 1609
rect 35937 1545 35940 1597
rect 35992 1545 35995 1597
rect 35937 1533 35995 1545
rect 35937 1481 35940 1533
rect 35992 1481 35995 1533
rect 35937 1469 35995 1481
rect 35937 1417 35940 1469
rect 35992 1417 35995 1469
rect 35937 1410 35949 1417
rect 35983 1410 35995 1417
rect 35937 1405 35995 1410
rect 35937 1353 35940 1405
rect 35992 1353 35995 1405
rect 35937 1341 35949 1353
rect 35983 1341 35995 1353
rect 35937 1289 35940 1341
rect 35992 1289 35995 1341
rect 35937 1277 35949 1289
rect 35983 1277 35995 1289
rect 35937 1225 35940 1277
rect 35992 1225 35995 1277
rect 35937 1213 35949 1225
rect 35983 1213 35995 1225
rect 35937 1161 35940 1213
rect 35992 1161 35995 1213
rect 35937 1147 35995 1161
rect 36033 3133 36091 3147
rect 36033 3081 36036 3133
rect 36088 3081 36091 3133
rect 36033 3069 36045 3081
rect 36079 3069 36091 3081
rect 36033 3017 36036 3069
rect 36088 3017 36091 3069
rect 36033 3005 36045 3017
rect 36079 3005 36091 3017
rect 36033 2953 36036 3005
rect 36088 2953 36091 3005
rect 36033 2941 36045 2953
rect 36079 2941 36091 2953
rect 36033 2889 36036 2941
rect 36088 2889 36091 2941
rect 36033 2884 36091 2889
rect 36033 2877 36045 2884
rect 36079 2877 36091 2884
rect 36033 2825 36036 2877
rect 36088 2825 36091 2877
rect 36033 2813 36091 2825
rect 36033 2761 36036 2813
rect 36088 2761 36091 2813
rect 36033 2749 36091 2761
rect 36033 2697 36036 2749
rect 36088 2697 36091 2749
rect 36033 2685 36091 2697
rect 36033 2633 36036 2685
rect 36088 2633 36091 2685
rect 36033 2621 36091 2633
rect 36033 2569 36036 2621
rect 36088 2569 36091 2621
rect 36033 2562 36045 2569
rect 36079 2562 36091 2569
rect 36033 2557 36091 2562
rect 36033 2505 36036 2557
rect 36088 2505 36091 2557
rect 36033 2493 36045 2505
rect 36079 2493 36091 2505
rect 36033 2441 36036 2493
rect 36088 2441 36091 2493
rect 36033 2429 36045 2441
rect 36079 2429 36091 2441
rect 36033 2377 36036 2429
rect 36088 2377 36091 2429
rect 36033 2365 36045 2377
rect 36079 2365 36091 2377
rect 36033 2313 36036 2365
rect 36088 2313 36091 2365
rect 36033 2308 36091 2313
rect 36033 2301 36045 2308
rect 36079 2301 36091 2308
rect 36033 2249 36036 2301
rect 36088 2249 36091 2301
rect 36033 2237 36091 2249
rect 36033 2185 36036 2237
rect 36088 2185 36091 2237
rect 36033 2173 36091 2185
rect 36033 2121 36036 2173
rect 36088 2121 36091 2173
rect 36033 2109 36091 2121
rect 36033 2057 36036 2109
rect 36088 2057 36091 2109
rect 36033 2045 36091 2057
rect 36033 1993 36036 2045
rect 36088 1993 36091 2045
rect 36033 1986 36045 1993
rect 36079 1986 36091 1993
rect 36033 1981 36091 1986
rect 36033 1929 36036 1981
rect 36088 1929 36091 1981
rect 36033 1917 36045 1929
rect 36079 1917 36091 1929
rect 36033 1865 36036 1917
rect 36088 1865 36091 1917
rect 36033 1853 36045 1865
rect 36079 1853 36091 1865
rect 36033 1801 36036 1853
rect 36088 1801 36091 1853
rect 36033 1789 36045 1801
rect 36079 1789 36091 1801
rect 36033 1737 36036 1789
rect 36088 1737 36091 1789
rect 36033 1732 36091 1737
rect 36033 1725 36045 1732
rect 36079 1725 36091 1732
rect 36033 1673 36036 1725
rect 36088 1673 36091 1725
rect 36033 1661 36091 1673
rect 36033 1609 36036 1661
rect 36088 1609 36091 1661
rect 36033 1597 36091 1609
rect 36033 1545 36036 1597
rect 36088 1545 36091 1597
rect 36033 1533 36091 1545
rect 36033 1481 36036 1533
rect 36088 1481 36091 1533
rect 36033 1469 36091 1481
rect 36033 1417 36036 1469
rect 36088 1417 36091 1469
rect 36033 1410 36045 1417
rect 36079 1410 36091 1417
rect 36033 1405 36091 1410
rect 36033 1353 36036 1405
rect 36088 1353 36091 1405
rect 36033 1341 36045 1353
rect 36079 1341 36091 1353
rect 36033 1289 36036 1341
rect 36088 1289 36091 1341
rect 36033 1277 36045 1289
rect 36079 1277 36091 1289
rect 36033 1225 36036 1277
rect 36088 1225 36091 1277
rect 36033 1213 36045 1225
rect 36079 1213 36091 1225
rect 36033 1161 36036 1213
rect 36088 1161 36091 1213
rect 36033 1147 36091 1161
rect 36129 3133 36187 3147
rect 36129 3081 36132 3133
rect 36184 3081 36187 3133
rect 36129 3069 36141 3081
rect 36175 3069 36187 3081
rect 36129 3017 36132 3069
rect 36184 3017 36187 3069
rect 36129 3005 36141 3017
rect 36175 3005 36187 3017
rect 36129 2953 36132 3005
rect 36184 2953 36187 3005
rect 36129 2941 36141 2953
rect 36175 2941 36187 2953
rect 36129 2889 36132 2941
rect 36184 2889 36187 2941
rect 36129 2884 36187 2889
rect 36129 2877 36141 2884
rect 36175 2877 36187 2884
rect 36129 2825 36132 2877
rect 36184 2825 36187 2877
rect 36129 2813 36187 2825
rect 36129 2761 36132 2813
rect 36184 2761 36187 2813
rect 36129 2749 36187 2761
rect 36129 2697 36132 2749
rect 36184 2697 36187 2749
rect 36129 2685 36187 2697
rect 36129 2633 36132 2685
rect 36184 2633 36187 2685
rect 36129 2621 36187 2633
rect 36129 2569 36132 2621
rect 36184 2569 36187 2621
rect 36129 2562 36141 2569
rect 36175 2562 36187 2569
rect 36129 2557 36187 2562
rect 36129 2505 36132 2557
rect 36184 2505 36187 2557
rect 36129 2493 36141 2505
rect 36175 2493 36187 2505
rect 36129 2441 36132 2493
rect 36184 2441 36187 2493
rect 36129 2429 36141 2441
rect 36175 2429 36187 2441
rect 36129 2377 36132 2429
rect 36184 2377 36187 2429
rect 36129 2365 36141 2377
rect 36175 2365 36187 2377
rect 36129 2313 36132 2365
rect 36184 2313 36187 2365
rect 36129 2308 36187 2313
rect 36129 2301 36141 2308
rect 36175 2301 36187 2308
rect 36129 2249 36132 2301
rect 36184 2249 36187 2301
rect 36129 2237 36187 2249
rect 36129 2185 36132 2237
rect 36184 2185 36187 2237
rect 36129 2173 36187 2185
rect 36129 2121 36132 2173
rect 36184 2121 36187 2173
rect 36129 2109 36187 2121
rect 36129 2057 36132 2109
rect 36184 2057 36187 2109
rect 36129 2045 36187 2057
rect 36129 1993 36132 2045
rect 36184 1993 36187 2045
rect 36129 1986 36141 1993
rect 36175 1986 36187 1993
rect 36129 1981 36187 1986
rect 36129 1929 36132 1981
rect 36184 1929 36187 1981
rect 36129 1917 36141 1929
rect 36175 1917 36187 1929
rect 36129 1865 36132 1917
rect 36184 1865 36187 1917
rect 36129 1853 36141 1865
rect 36175 1853 36187 1865
rect 36129 1801 36132 1853
rect 36184 1801 36187 1853
rect 36129 1789 36141 1801
rect 36175 1789 36187 1801
rect 36129 1737 36132 1789
rect 36184 1737 36187 1789
rect 36129 1732 36187 1737
rect 36129 1725 36141 1732
rect 36175 1725 36187 1732
rect 36129 1673 36132 1725
rect 36184 1673 36187 1725
rect 36129 1661 36187 1673
rect 36129 1609 36132 1661
rect 36184 1609 36187 1661
rect 36129 1597 36187 1609
rect 36129 1545 36132 1597
rect 36184 1545 36187 1597
rect 36129 1533 36187 1545
rect 36129 1481 36132 1533
rect 36184 1481 36187 1533
rect 36129 1469 36187 1481
rect 36129 1417 36132 1469
rect 36184 1417 36187 1469
rect 36129 1410 36141 1417
rect 36175 1410 36187 1417
rect 36129 1405 36187 1410
rect 36129 1353 36132 1405
rect 36184 1353 36187 1405
rect 36129 1341 36141 1353
rect 36175 1341 36187 1353
rect 36129 1289 36132 1341
rect 36184 1289 36187 1341
rect 36129 1277 36141 1289
rect 36175 1277 36187 1289
rect 36129 1225 36132 1277
rect 36184 1225 36187 1277
rect 36129 1213 36141 1225
rect 36175 1213 36187 1225
rect 36129 1161 36132 1213
rect 36184 1161 36187 1213
rect 36129 1147 36187 1161
rect 36228 3133 36280 3147
rect 36228 3069 36237 3081
rect 36271 3069 36280 3081
rect 36228 3005 36237 3017
rect 36271 3005 36280 3017
rect 36228 2941 36237 2953
rect 36271 2941 36280 2953
rect 36228 2884 36280 2889
rect 36228 2877 36237 2884
rect 36271 2877 36280 2884
rect 36228 2813 36280 2825
rect 36228 2749 36280 2761
rect 36228 2685 36280 2697
rect 36228 2621 36280 2633
rect 36228 2562 36237 2569
rect 36271 2562 36280 2569
rect 36228 2557 36280 2562
rect 36228 2493 36237 2505
rect 36271 2493 36280 2505
rect 36228 2429 36237 2441
rect 36271 2429 36280 2441
rect 36228 2365 36237 2377
rect 36271 2365 36280 2377
rect 36228 2308 36280 2313
rect 36228 2301 36237 2308
rect 36271 2301 36280 2308
rect 36228 2237 36280 2249
rect 36228 2173 36280 2185
rect 36228 2109 36280 2121
rect 36228 2045 36280 2057
rect 36228 1986 36237 1993
rect 36271 1986 36280 1993
rect 36228 1981 36280 1986
rect 36228 1917 36237 1929
rect 36271 1917 36280 1929
rect 36228 1853 36237 1865
rect 36271 1853 36280 1865
rect 36228 1789 36237 1801
rect 36271 1789 36280 1801
rect 36228 1732 36280 1737
rect 36228 1725 36237 1732
rect 36271 1725 36280 1732
rect 36228 1661 36280 1673
rect 36228 1597 36280 1609
rect 36228 1533 36280 1545
rect 36228 1469 36280 1481
rect 36228 1410 36237 1417
rect 36271 1410 36280 1417
rect 36228 1405 36280 1410
rect 36228 1341 36237 1353
rect 36271 1341 36280 1353
rect 36228 1277 36237 1289
rect 36271 1277 36280 1289
rect 36228 1213 36237 1225
rect 36271 1213 36280 1225
rect 36228 1147 36280 1161
rect 36321 3133 36379 3147
rect 36321 3081 36324 3133
rect 36376 3081 36379 3133
rect 36321 3069 36333 3081
rect 36367 3069 36379 3081
rect 36321 3017 36324 3069
rect 36376 3017 36379 3069
rect 36321 3005 36333 3017
rect 36367 3005 36379 3017
rect 36321 2953 36324 3005
rect 36376 2953 36379 3005
rect 36321 2941 36333 2953
rect 36367 2941 36379 2953
rect 36321 2889 36324 2941
rect 36376 2889 36379 2941
rect 36321 2884 36379 2889
rect 36321 2877 36333 2884
rect 36367 2877 36379 2884
rect 36321 2825 36324 2877
rect 36376 2825 36379 2877
rect 36321 2813 36379 2825
rect 36321 2761 36324 2813
rect 36376 2761 36379 2813
rect 36321 2749 36379 2761
rect 36321 2697 36324 2749
rect 36376 2697 36379 2749
rect 36321 2685 36379 2697
rect 36321 2633 36324 2685
rect 36376 2633 36379 2685
rect 36321 2621 36379 2633
rect 36321 2569 36324 2621
rect 36376 2569 36379 2621
rect 36321 2562 36333 2569
rect 36367 2562 36379 2569
rect 36321 2557 36379 2562
rect 36321 2505 36324 2557
rect 36376 2505 36379 2557
rect 36321 2493 36333 2505
rect 36367 2493 36379 2505
rect 36321 2441 36324 2493
rect 36376 2441 36379 2493
rect 36321 2429 36333 2441
rect 36367 2429 36379 2441
rect 36321 2377 36324 2429
rect 36376 2377 36379 2429
rect 36321 2365 36333 2377
rect 36367 2365 36379 2377
rect 36321 2313 36324 2365
rect 36376 2313 36379 2365
rect 36321 2308 36379 2313
rect 36321 2301 36333 2308
rect 36367 2301 36379 2308
rect 36321 2249 36324 2301
rect 36376 2249 36379 2301
rect 36321 2237 36379 2249
rect 36321 2185 36324 2237
rect 36376 2185 36379 2237
rect 36321 2173 36379 2185
rect 36321 2121 36324 2173
rect 36376 2121 36379 2173
rect 36321 2109 36379 2121
rect 36321 2057 36324 2109
rect 36376 2057 36379 2109
rect 36321 2045 36379 2057
rect 36321 1993 36324 2045
rect 36376 1993 36379 2045
rect 36321 1986 36333 1993
rect 36367 1986 36379 1993
rect 36321 1981 36379 1986
rect 36321 1929 36324 1981
rect 36376 1929 36379 1981
rect 36321 1917 36333 1929
rect 36367 1917 36379 1929
rect 36321 1865 36324 1917
rect 36376 1865 36379 1917
rect 36321 1853 36333 1865
rect 36367 1853 36379 1865
rect 36321 1801 36324 1853
rect 36376 1801 36379 1853
rect 36321 1789 36333 1801
rect 36367 1789 36379 1801
rect 36321 1737 36324 1789
rect 36376 1737 36379 1789
rect 36321 1732 36379 1737
rect 36321 1725 36333 1732
rect 36367 1725 36379 1732
rect 36321 1673 36324 1725
rect 36376 1673 36379 1725
rect 36321 1661 36379 1673
rect 36321 1609 36324 1661
rect 36376 1609 36379 1661
rect 36321 1597 36379 1609
rect 36321 1545 36324 1597
rect 36376 1545 36379 1597
rect 36321 1533 36379 1545
rect 36321 1481 36324 1533
rect 36376 1481 36379 1533
rect 36321 1469 36379 1481
rect 36321 1417 36324 1469
rect 36376 1417 36379 1469
rect 36321 1410 36333 1417
rect 36367 1410 36379 1417
rect 36321 1405 36379 1410
rect 36321 1353 36324 1405
rect 36376 1353 36379 1405
rect 36321 1341 36333 1353
rect 36367 1341 36379 1353
rect 36321 1289 36324 1341
rect 36376 1289 36379 1341
rect 36321 1277 36333 1289
rect 36367 1277 36379 1289
rect 36321 1225 36324 1277
rect 36376 1225 36379 1277
rect 36321 1213 36333 1225
rect 36367 1213 36379 1225
rect 36321 1161 36324 1213
rect 36376 1161 36379 1213
rect 36321 1147 36379 1161
rect 36417 3133 36475 3147
rect 36417 3081 36420 3133
rect 36472 3081 36475 3133
rect 36417 3069 36429 3081
rect 36463 3069 36475 3081
rect 36417 3017 36420 3069
rect 36472 3017 36475 3069
rect 36417 3005 36429 3017
rect 36463 3005 36475 3017
rect 36417 2953 36420 3005
rect 36472 2953 36475 3005
rect 36417 2941 36429 2953
rect 36463 2941 36475 2953
rect 36417 2889 36420 2941
rect 36472 2889 36475 2941
rect 36417 2884 36475 2889
rect 36417 2877 36429 2884
rect 36463 2877 36475 2884
rect 36417 2825 36420 2877
rect 36472 2825 36475 2877
rect 36417 2813 36475 2825
rect 36417 2761 36420 2813
rect 36472 2761 36475 2813
rect 36417 2749 36475 2761
rect 36417 2697 36420 2749
rect 36472 2697 36475 2749
rect 36417 2685 36475 2697
rect 36417 2633 36420 2685
rect 36472 2633 36475 2685
rect 36417 2621 36475 2633
rect 36417 2569 36420 2621
rect 36472 2569 36475 2621
rect 36417 2562 36429 2569
rect 36463 2562 36475 2569
rect 36417 2557 36475 2562
rect 36417 2505 36420 2557
rect 36472 2505 36475 2557
rect 36417 2493 36429 2505
rect 36463 2493 36475 2505
rect 36417 2441 36420 2493
rect 36472 2441 36475 2493
rect 36417 2429 36429 2441
rect 36463 2429 36475 2441
rect 36417 2377 36420 2429
rect 36472 2377 36475 2429
rect 36417 2365 36429 2377
rect 36463 2365 36475 2377
rect 36417 2313 36420 2365
rect 36472 2313 36475 2365
rect 36417 2308 36475 2313
rect 36417 2301 36429 2308
rect 36463 2301 36475 2308
rect 36417 2249 36420 2301
rect 36472 2249 36475 2301
rect 36417 2237 36475 2249
rect 36417 2185 36420 2237
rect 36472 2185 36475 2237
rect 36417 2173 36475 2185
rect 36417 2121 36420 2173
rect 36472 2121 36475 2173
rect 36417 2109 36475 2121
rect 36417 2057 36420 2109
rect 36472 2057 36475 2109
rect 36417 2045 36475 2057
rect 36417 1993 36420 2045
rect 36472 1993 36475 2045
rect 36417 1986 36429 1993
rect 36463 1986 36475 1993
rect 36417 1981 36475 1986
rect 36417 1929 36420 1981
rect 36472 1929 36475 1981
rect 36417 1917 36429 1929
rect 36463 1917 36475 1929
rect 36417 1865 36420 1917
rect 36472 1865 36475 1917
rect 36417 1853 36429 1865
rect 36463 1853 36475 1865
rect 36417 1801 36420 1853
rect 36472 1801 36475 1853
rect 36417 1789 36429 1801
rect 36463 1789 36475 1801
rect 36417 1737 36420 1789
rect 36472 1737 36475 1789
rect 36417 1732 36475 1737
rect 36417 1725 36429 1732
rect 36463 1725 36475 1732
rect 36417 1673 36420 1725
rect 36472 1673 36475 1725
rect 36417 1661 36475 1673
rect 36417 1609 36420 1661
rect 36472 1609 36475 1661
rect 36417 1597 36475 1609
rect 36417 1545 36420 1597
rect 36472 1545 36475 1597
rect 36417 1533 36475 1545
rect 36417 1481 36420 1533
rect 36472 1481 36475 1533
rect 36417 1469 36475 1481
rect 36417 1417 36420 1469
rect 36472 1417 36475 1469
rect 36417 1410 36429 1417
rect 36463 1410 36475 1417
rect 36417 1405 36475 1410
rect 36417 1353 36420 1405
rect 36472 1353 36475 1405
rect 36417 1341 36429 1353
rect 36463 1341 36475 1353
rect 36417 1289 36420 1341
rect 36472 1289 36475 1341
rect 36417 1277 36429 1289
rect 36463 1277 36475 1289
rect 36417 1225 36420 1277
rect 36472 1225 36475 1277
rect 36417 1213 36429 1225
rect 36463 1213 36475 1225
rect 36417 1161 36420 1213
rect 36472 1161 36475 1213
rect 36417 1147 36475 1161
rect 36513 3133 36571 3147
rect 36513 3081 36516 3133
rect 36568 3081 36571 3133
rect 36513 3069 36525 3081
rect 36559 3069 36571 3081
rect 36513 3017 36516 3069
rect 36568 3017 36571 3069
rect 36513 3005 36525 3017
rect 36559 3005 36571 3017
rect 36513 2953 36516 3005
rect 36568 2953 36571 3005
rect 36513 2941 36525 2953
rect 36559 2941 36571 2953
rect 36513 2889 36516 2941
rect 36568 2889 36571 2941
rect 36513 2884 36571 2889
rect 36513 2877 36525 2884
rect 36559 2877 36571 2884
rect 36513 2825 36516 2877
rect 36568 2825 36571 2877
rect 36513 2813 36571 2825
rect 36513 2761 36516 2813
rect 36568 2761 36571 2813
rect 36513 2749 36571 2761
rect 36513 2697 36516 2749
rect 36568 2697 36571 2749
rect 36513 2685 36571 2697
rect 36513 2633 36516 2685
rect 36568 2633 36571 2685
rect 36513 2621 36571 2633
rect 36513 2569 36516 2621
rect 36568 2569 36571 2621
rect 36513 2562 36525 2569
rect 36559 2562 36571 2569
rect 36513 2557 36571 2562
rect 36513 2505 36516 2557
rect 36568 2505 36571 2557
rect 36513 2493 36525 2505
rect 36559 2493 36571 2505
rect 36513 2441 36516 2493
rect 36568 2441 36571 2493
rect 36513 2429 36525 2441
rect 36559 2429 36571 2441
rect 36513 2377 36516 2429
rect 36568 2377 36571 2429
rect 36513 2365 36525 2377
rect 36559 2365 36571 2377
rect 36513 2313 36516 2365
rect 36568 2313 36571 2365
rect 36513 2308 36571 2313
rect 36513 2301 36525 2308
rect 36559 2301 36571 2308
rect 36513 2249 36516 2301
rect 36568 2249 36571 2301
rect 36513 2237 36571 2249
rect 36513 2185 36516 2237
rect 36568 2185 36571 2237
rect 36513 2173 36571 2185
rect 36513 2121 36516 2173
rect 36568 2121 36571 2173
rect 36513 2109 36571 2121
rect 36513 2057 36516 2109
rect 36568 2057 36571 2109
rect 36513 2045 36571 2057
rect 36513 1993 36516 2045
rect 36568 1993 36571 2045
rect 36513 1986 36525 1993
rect 36559 1986 36571 1993
rect 36513 1981 36571 1986
rect 36513 1929 36516 1981
rect 36568 1929 36571 1981
rect 36513 1917 36525 1929
rect 36559 1917 36571 1929
rect 36513 1865 36516 1917
rect 36568 1865 36571 1917
rect 36513 1853 36525 1865
rect 36559 1853 36571 1865
rect 36513 1801 36516 1853
rect 36568 1801 36571 1853
rect 36513 1789 36525 1801
rect 36559 1789 36571 1801
rect 36513 1737 36516 1789
rect 36568 1737 36571 1789
rect 36513 1732 36571 1737
rect 36513 1725 36525 1732
rect 36559 1725 36571 1732
rect 36513 1673 36516 1725
rect 36568 1673 36571 1725
rect 36513 1661 36571 1673
rect 36513 1609 36516 1661
rect 36568 1609 36571 1661
rect 36513 1597 36571 1609
rect 36513 1545 36516 1597
rect 36568 1545 36571 1597
rect 36513 1533 36571 1545
rect 36513 1481 36516 1533
rect 36568 1481 36571 1533
rect 36513 1469 36571 1481
rect 36513 1417 36516 1469
rect 36568 1417 36571 1469
rect 36513 1410 36525 1417
rect 36559 1410 36571 1417
rect 36513 1405 36571 1410
rect 36513 1353 36516 1405
rect 36568 1353 36571 1405
rect 36513 1341 36525 1353
rect 36559 1341 36571 1353
rect 36513 1289 36516 1341
rect 36568 1289 36571 1341
rect 36513 1277 36525 1289
rect 36559 1277 36571 1289
rect 36513 1225 36516 1277
rect 36568 1225 36571 1277
rect 36513 1213 36525 1225
rect 36559 1213 36571 1225
rect 36513 1161 36516 1213
rect 36568 1161 36571 1213
rect 36513 1147 36571 1161
rect 36612 3133 36664 3147
rect 36612 3069 36621 3081
rect 36655 3069 36664 3081
rect 36612 3005 36621 3017
rect 36655 3005 36664 3017
rect 36612 2941 36621 2953
rect 36655 2941 36664 2953
rect 36612 2884 36664 2889
rect 36612 2877 36621 2884
rect 36655 2877 36664 2884
rect 36612 2813 36664 2825
rect 36612 2749 36664 2761
rect 36612 2685 36664 2697
rect 36612 2621 36664 2633
rect 36612 2562 36621 2569
rect 36655 2562 36664 2569
rect 36612 2557 36664 2562
rect 36612 2493 36621 2505
rect 36655 2493 36664 2505
rect 36612 2429 36621 2441
rect 36655 2429 36664 2441
rect 36612 2365 36621 2377
rect 36655 2365 36664 2377
rect 36612 2308 36664 2313
rect 36612 2301 36621 2308
rect 36655 2301 36664 2308
rect 36612 2237 36664 2249
rect 36612 2173 36664 2185
rect 36612 2109 36664 2121
rect 36612 2045 36664 2057
rect 36612 1986 36621 1993
rect 36655 1986 36664 1993
rect 36612 1981 36664 1986
rect 36612 1917 36621 1929
rect 36655 1917 36664 1929
rect 36612 1853 36621 1865
rect 36655 1853 36664 1865
rect 36612 1789 36621 1801
rect 36655 1789 36664 1801
rect 36612 1732 36664 1737
rect 36612 1725 36621 1732
rect 36655 1725 36664 1732
rect 36612 1661 36664 1673
rect 36612 1597 36664 1609
rect 36612 1533 36664 1545
rect 36612 1469 36664 1481
rect 36612 1410 36621 1417
rect 36655 1410 36664 1417
rect 36612 1405 36664 1410
rect 36612 1341 36621 1353
rect 36655 1341 36664 1353
rect 36612 1277 36621 1289
rect 36655 1277 36664 1289
rect 36612 1213 36621 1225
rect 36655 1213 36664 1225
rect 36612 1147 36664 1161
rect 36705 3133 36763 3147
rect 36705 3081 36708 3133
rect 36760 3081 36763 3133
rect 36705 3069 36717 3081
rect 36751 3069 36763 3081
rect 36705 3017 36708 3069
rect 36760 3017 36763 3069
rect 36705 3005 36717 3017
rect 36751 3005 36763 3017
rect 36705 2953 36708 3005
rect 36760 2953 36763 3005
rect 36705 2941 36717 2953
rect 36751 2941 36763 2953
rect 36705 2889 36708 2941
rect 36760 2889 36763 2941
rect 36705 2884 36763 2889
rect 36705 2877 36717 2884
rect 36751 2877 36763 2884
rect 36705 2825 36708 2877
rect 36760 2825 36763 2877
rect 36705 2813 36763 2825
rect 36705 2761 36708 2813
rect 36760 2761 36763 2813
rect 36705 2749 36763 2761
rect 36705 2697 36708 2749
rect 36760 2697 36763 2749
rect 36705 2685 36763 2697
rect 36705 2633 36708 2685
rect 36760 2633 36763 2685
rect 36705 2621 36763 2633
rect 36705 2569 36708 2621
rect 36760 2569 36763 2621
rect 36705 2562 36717 2569
rect 36751 2562 36763 2569
rect 36705 2557 36763 2562
rect 36705 2505 36708 2557
rect 36760 2505 36763 2557
rect 36705 2493 36717 2505
rect 36751 2493 36763 2505
rect 36705 2441 36708 2493
rect 36760 2441 36763 2493
rect 36705 2429 36717 2441
rect 36751 2429 36763 2441
rect 36705 2377 36708 2429
rect 36760 2377 36763 2429
rect 36705 2365 36717 2377
rect 36751 2365 36763 2377
rect 36705 2313 36708 2365
rect 36760 2313 36763 2365
rect 36705 2308 36763 2313
rect 36705 2301 36717 2308
rect 36751 2301 36763 2308
rect 36705 2249 36708 2301
rect 36760 2249 36763 2301
rect 36705 2237 36763 2249
rect 36705 2185 36708 2237
rect 36760 2185 36763 2237
rect 36705 2173 36763 2185
rect 36705 2121 36708 2173
rect 36760 2121 36763 2173
rect 36705 2109 36763 2121
rect 36705 2057 36708 2109
rect 36760 2057 36763 2109
rect 36705 2045 36763 2057
rect 36705 1993 36708 2045
rect 36760 1993 36763 2045
rect 36705 1986 36717 1993
rect 36751 1986 36763 1993
rect 36705 1981 36763 1986
rect 36705 1929 36708 1981
rect 36760 1929 36763 1981
rect 36705 1917 36717 1929
rect 36751 1917 36763 1929
rect 36705 1865 36708 1917
rect 36760 1865 36763 1917
rect 36705 1853 36717 1865
rect 36751 1853 36763 1865
rect 36705 1801 36708 1853
rect 36760 1801 36763 1853
rect 36705 1789 36717 1801
rect 36751 1789 36763 1801
rect 36705 1737 36708 1789
rect 36760 1737 36763 1789
rect 36705 1732 36763 1737
rect 36705 1725 36717 1732
rect 36751 1725 36763 1732
rect 36705 1673 36708 1725
rect 36760 1673 36763 1725
rect 36705 1661 36763 1673
rect 36705 1609 36708 1661
rect 36760 1609 36763 1661
rect 36705 1597 36763 1609
rect 36705 1545 36708 1597
rect 36760 1545 36763 1597
rect 36705 1533 36763 1545
rect 36705 1481 36708 1533
rect 36760 1481 36763 1533
rect 36705 1469 36763 1481
rect 36705 1417 36708 1469
rect 36760 1417 36763 1469
rect 36705 1410 36717 1417
rect 36751 1410 36763 1417
rect 36705 1405 36763 1410
rect 36705 1353 36708 1405
rect 36760 1353 36763 1405
rect 36705 1341 36717 1353
rect 36751 1341 36763 1353
rect 36705 1289 36708 1341
rect 36760 1289 36763 1341
rect 36705 1277 36717 1289
rect 36751 1277 36763 1289
rect 36705 1225 36708 1277
rect 36760 1225 36763 1277
rect 36705 1213 36717 1225
rect 36751 1213 36763 1225
rect 36705 1161 36708 1213
rect 36760 1161 36763 1213
rect 36705 1147 36763 1161
rect 36801 3133 36859 3147
rect 36801 3081 36804 3133
rect 36856 3081 36859 3133
rect 36801 3069 36813 3081
rect 36847 3069 36859 3081
rect 36801 3017 36804 3069
rect 36856 3017 36859 3069
rect 36801 3005 36813 3017
rect 36847 3005 36859 3017
rect 36801 2953 36804 3005
rect 36856 2953 36859 3005
rect 36801 2941 36813 2953
rect 36847 2941 36859 2953
rect 36801 2889 36804 2941
rect 36856 2889 36859 2941
rect 36801 2884 36859 2889
rect 36801 2877 36813 2884
rect 36847 2877 36859 2884
rect 36801 2825 36804 2877
rect 36856 2825 36859 2877
rect 36801 2813 36859 2825
rect 36801 2761 36804 2813
rect 36856 2761 36859 2813
rect 36801 2749 36859 2761
rect 36801 2697 36804 2749
rect 36856 2697 36859 2749
rect 36801 2685 36859 2697
rect 36801 2633 36804 2685
rect 36856 2633 36859 2685
rect 36801 2621 36859 2633
rect 36801 2569 36804 2621
rect 36856 2569 36859 2621
rect 36801 2562 36813 2569
rect 36847 2562 36859 2569
rect 36801 2557 36859 2562
rect 36801 2505 36804 2557
rect 36856 2505 36859 2557
rect 36801 2493 36813 2505
rect 36847 2493 36859 2505
rect 36801 2441 36804 2493
rect 36856 2441 36859 2493
rect 36801 2429 36813 2441
rect 36847 2429 36859 2441
rect 36801 2377 36804 2429
rect 36856 2377 36859 2429
rect 36801 2365 36813 2377
rect 36847 2365 36859 2377
rect 36801 2313 36804 2365
rect 36856 2313 36859 2365
rect 36801 2308 36859 2313
rect 36801 2301 36813 2308
rect 36847 2301 36859 2308
rect 36801 2249 36804 2301
rect 36856 2249 36859 2301
rect 36801 2237 36859 2249
rect 36801 2185 36804 2237
rect 36856 2185 36859 2237
rect 36801 2173 36859 2185
rect 36801 2121 36804 2173
rect 36856 2121 36859 2173
rect 36801 2109 36859 2121
rect 36801 2057 36804 2109
rect 36856 2057 36859 2109
rect 36801 2045 36859 2057
rect 36801 1993 36804 2045
rect 36856 1993 36859 2045
rect 36801 1986 36813 1993
rect 36847 1986 36859 1993
rect 36801 1981 36859 1986
rect 36801 1929 36804 1981
rect 36856 1929 36859 1981
rect 36801 1917 36813 1929
rect 36847 1917 36859 1929
rect 36801 1865 36804 1917
rect 36856 1865 36859 1917
rect 36801 1853 36813 1865
rect 36847 1853 36859 1865
rect 36801 1801 36804 1853
rect 36856 1801 36859 1853
rect 36801 1789 36813 1801
rect 36847 1789 36859 1801
rect 36801 1737 36804 1789
rect 36856 1737 36859 1789
rect 36801 1732 36859 1737
rect 36801 1725 36813 1732
rect 36847 1725 36859 1732
rect 36801 1673 36804 1725
rect 36856 1673 36859 1725
rect 36801 1661 36859 1673
rect 36801 1609 36804 1661
rect 36856 1609 36859 1661
rect 36801 1597 36859 1609
rect 36801 1545 36804 1597
rect 36856 1545 36859 1597
rect 36801 1533 36859 1545
rect 36801 1481 36804 1533
rect 36856 1481 36859 1533
rect 36801 1469 36859 1481
rect 36801 1417 36804 1469
rect 36856 1417 36859 1469
rect 36801 1410 36813 1417
rect 36847 1410 36859 1417
rect 36801 1405 36859 1410
rect 36801 1353 36804 1405
rect 36856 1353 36859 1405
rect 36801 1341 36813 1353
rect 36847 1341 36859 1353
rect 36801 1289 36804 1341
rect 36856 1289 36859 1341
rect 36801 1277 36813 1289
rect 36847 1277 36859 1289
rect 36801 1225 36804 1277
rect 36856 1225 36859 1277
rect 36801 1213 36813 1225
rect 36847 1213 36859 1225
rect 36801 1161 36804 1213
rect 36856 1161 36859 1213
rect 36801 1147 36859 1161
rect 36897 3133 36955 3147
rect 36897 3081 36900 3133
rect 36952 3081 36955 3133
rect 36897 3069 36909 3081
rect 36943 3069 36955 3081
rect 36897 3017 36900 3069
rect 36952 3017 36955 3069
rect 36897 3005 36909 3017
rect 36943 3005 36955 3017
rect 36897 2953 36900 3005
rect 36952 2953 36955 3005
rect 36897 2941 36909 2953
rect 36943 2941 36955 2953
rect 36897 2889 36900 2941
rect 36952 2889 36955 2941
rect 36897 2884 36955 2889
rect 36897 2877 36909 2884
rect 36943 2877 36955 2884
rect 36897 2825 36900 2877
rect 36952 2825 36955 2877
rect 36897 2813 36955 2825
rect 36897 2761 36900 2813
rect 36952 2761 36955 2813
rect 36897 2749 36955 2761
rect 36897 2697 36900 2749
rect 36952 2697 36955 2749
rect 36897 2685 36955 2697
rect 36897 2633 36900 2685
rect 36952 2633 36955 2685
rect 36897 2621 36955 2633
rect 36897 2569 36900 2621
rect 36952 2569 36955 2621
rect 36897 2562 36909 2569
rect 36943 2562 36955 2569
rect 36897 2557 36955 2562
rect 36897 2505 36900 2557
rect 36952 2505 36955 2557
rect 36897 2493 36909 2505
rect 36943 2493 36955 2505
rect 36897 2441 36900 2493
rect 36952 2441 36955 2493
rect 36897 2429 36909 2441
rect 36943 2429 36955 2441
rect 36897 2377 36900 2429
rect 36952 2377 36955 2429
rect 36897 2365 36909 2377
rect 36943 2365 36955 2377
rect 36897 2313 36900 2365
rect 36952 2313 36955 2365
rect 36897 2308 36955 2313
rect 36897 2301 36909 2308
rect 36943 2301 36955 2308
rect 36897 2249 36900 2301
rect 36952 2249 36955 2301
rect 36897 2237 36955 2249
rect 36897 2185 36900 2237
rect 36952 2185 36955 2237
rect 36897 2173 36955 2185
rect 36897 2121 36900 2173
rect 36952 2121 36955 2173
rect 36897 2109 36955 2121
rect 36897 2057 36900 2109
rect 36952 2057 36955 2109
rect 36897 2045 36955 2057
rect 36897 1993 36900 2045
rect 36952 1993 36955 2045
rect 36897 1986 36909 1993
rect 36943 1986 36955 1993
rect 36897 1981 36955 1986
rect 36897 1929 36900 1981
rect 36952 1929 36955 1981
rect 36897 1917 36909 1929
rect 36943 1917 36955 1929
rect 36897 1865 36900 1917
rect 36952 1865 36955 1917
rect 36897 1853 36909 1865
rect 36943 1853 36955 1865
rect 36897 1801 36900 1853
rect 36952 1801 36955 1853
rect 36897 1789 36909 1801
rect 36943 1789 36955 1801
rect 36897 1737 36900 1789
rect 36952 1737 36955 1789
rect 36897 1732 36955 1737
rect 36897 1725 36909 1732
rect 36943 1725 36955 1732
rect 36897 1673 36900 1725
rect 36952 1673 36955 1725
rect 36897 1661 36955 1673
rect 36897 1609 36900 1661
rect 36952 1609 36955 1661
rect 36897 1597 36955 1609
rect 36897 1545 36900 1597
rect 36952 1545 36955 1597
rect 36897 1533 36955 1545
rect 36897 1481 36900 1533
rect 36952 1481 36955 1533
rect 36897 1469 36955 1481
rect 36897 1417 36900 1469
rect 36952 1417 36955 1469
rect 36897 1410 36909 1417
rect 36943 1410 36955 1417
rect 36897 1405 36955 1410
rect 36897 1353 36900 1405
rect 36952 1353 36955 1405
rect 36897 1341 36909 1353
rect 36943 1341 36955 1353
rect 36897 1289 36900 1341
rect 36952 1289 36955 1341
rect 36897 1277 36909 1289
rect 36943 1277 36955 1289
rect 36897 1225 36900 1277
rect 36952 1225 36955 1277
rect 36897 1213 36909 1225
rect 36943 1213 36955 1225
rect 36897 1161 36900 1213
rect 36952 1161 36955 1213
rect 36897 1147 36955 1161
rect 36996 3133 37048 3147
rect 36996 3069 37005 3081
rect 37039 3069 37048 3081
rect 36996 3005 37005 3017
rect 37039 3005 37048 3017
rect 36996 2941 37005 2953
rect 37039 2941 37048 2953
rect 36996 2884 37048 2889
rect 36996 2877 37005 2884
rect 37039 2877 37048 2884
rect 36996 2813 37048 2825
rect 36996 2749 37048 2761
rect 36996 2685 37048 2697
rect 36996 2621 37048 2633
rect 36996 2562 37005 2569
rect 37039 2562 37048 2569
rect 36996 2557 37048 2562
rect 36996 2493 37005 2505
rect 37039 2493 37048 2505
rect 36996 2429 37005 2441
rect 37039 2429 37048 2441
rect 36996 2365 37005 2377
rect 37039 2365 37048 2377
rect 36996 2308 37048 2313
rect 36996 2301 37005 2308
rect 37039 2301 37048 2308
rect 36996 2237 37048 2249
rect 36996 2173 37048 2185
rect 36996 2109 37048 2121
rect 36996 2045 37048 2057
rect 36996 1986 37005 1993
rect 37039 1986 37048 1993
rect 36996 1981 37048 1986
rect 36996 1917 37005 1929
rect 37039 1917 37048 1929
rect 36996 1853 37005 1865
rect 37039 1853 37048 1865
rect 36996 1789 37005 1801
rect 37039 1789 37048 1801
rect 36996 1732 37048 1737
rect 36996 1725 37005 1732
rect 37039 1725 37048 1732
rect 36996 1661 37048 1673
rect 36996 1597 37048 1609
rect 36996 1533 37048 1545
rect 36996 1469 37048 1481
rect 36996 1410 37005 1417
rect 37039 1410 37048 1417
rect 36996 1405 37048 1410
rect 36996 1341 37005 1353
rect 37039 1341 37048 1353
rect 36996 1277 37005 1289
rect 37039 1277 37048 1289
rect 36996 1213 37005 1225
rect 37039 1213 37048 1225
rect 36996 1147 37048 1161
rect 37089 3133 37147 3147
rect 37089 3081 37092 3133
rect 37144 3081 37147 3133
rect 37089 3069 37101 3081
rect 37135 3069 37147 3081
rect 37089 3017 37092 3069
rect 37144 3017 37147 3069
rect 37089 3005 37101 3017
rect 37135 3005 37147 3017
rect 37089 2953 37092 3005
rect 37144 2953 37147 3005
rect 37089 2941 37101 2953
rect 37135 2941 37147 2953
rect 37089 2889 37092 2941
rect 37144 2889 37147 2941
rect 37089 2884 37147 2889
rect 37089 2877 37101 2884
rect 37135 2877 37147 2884
rect 37089 2825 37092 2877
rect 37144 2825 37147 2877
rect 37089 2813 37147 2825
rect 37089 2761 37092 2813
rect 37144 2761 37147 2813
rect 37089 2749 37147 2761
rect 37089 2697 37092 2749
rect 37144 2697 37147 2749
rect 37089 2685 37147 2697
rect 37089 2633 37092 2685
rect 37144 2633 37147 2685
rect 37089 2621 37147 2633
rect 37089 2569 37092 2621
rect 37144 2569 37147 2621
rect 37089 2562 37101 2569
rect 37135 2562 37147 2569
rect 37089 2557 37147 2562
rect 37089 2505 37092 2557
rect 37144 2505 37147 2557
rect 37089 2493 37101 2505
rect 37135 2493 37147 2505
rect 37089 2441 37092 2493
rect 37144 2441 37147 2493
rect 37089 2429 37101 2441
rect 37135 2429 37147 2441
rect 37089 2377 37092 2429
rect 37144 2377 37147 2429
rect 37089 2365 37101 2377
rect 37135 2365 37147 2377
rect 37089 2313 37092 2365
rect 37144 2313 37147 2365
rect 37089 2308 37147 2313
rect 37089 2301 37101 2308
rect 37135 2301 37147 2308
rect 37089 2249 37092 2301
rect 37144 2249 37147 2301
rect 37089 2237 37147 2249
rect 37089 2185 37092 2237
rect 37144 2185 37147 2237
rect 37089 2173 37147 2185
rect 37089 2121 37092 2173
rect 37144 2121 37147 2173
rect 37089 2109 37147 2121
rect 37089 2057 37092 2109
rect 37144 2057 37147 2109
rect 37089 2045 37147 2057
rect 37089 1993 37092 2045
rect 37144 1993 37147 2045
rect 37089 1986 37101 1993
rect 37135 1986 37147 1993
rect 37089 1981 37147 1986
rect 37089 1929 37092 1981
rect 37144 1929 37147 1981
rect 37089 1917 37101 1929
rect 37135 1917 37147 1929
rect 37089 1865 37092 1917
rect 37144 1865 37147 1917
rect 37089 1853 37101 1865
rect 37135 1853 37147 1865
rect 37089 1801 37092 1853
rect 37144 1801 37147 1853
rect 37089 1789 37101 1801
rect 37135 1789 37147 1801
rect 37089 1737 37092 1789
rect 37144 1737 37147 1789
rect 37089 1732 37147 1737
rect 37089 1725 37101 1732
rect 37135 1725 37147 1732
rect 37089 1673 37092 1725
rect 37144 1673 37147 1725
rect 37089 1661 37147 1673
rect 37089 1609 37092 1661
rect 37144 1609 37147 1661
rect 37089 1597 37147 1609
rect 37089 1545 37092 1597
rect 37144 1545 37147 1597
rect 37089 1533 37147 1545
rect 37089 1481 37092 1533
rect 37144 1481 37147 1533
rect 37089 1469 37147 1481
rect 37089 1417 37092 1469
rect 37144 1417 37147 1469
rect 37089 1410 37101 1417
rect 37135 1410 37147 1417
rect 37089 1405 37147 1410
rect 37089 1353 37092 1405
rect 37144 1353 37147 1405
rect 37089 1341 37101 1353
rect 37135 1341 37147 1353
rect 37089 1289 37092 1341
rect 37144 1289 37147 1341
rect 37089 1277 37101 1289
rect 37135 1277 37147 1289
rect 37089 1225 37092 1277
rect 37144 1225 37147 1277
rect 37089 1213 37101 1225
rect 37135 1213 37147 1225
rect 37089 1161 37092 1213
rect 37144 1161 37147 1213
rect 37089 1147 37147 1161
rect 37185 3133 37243 3147
rect 37185 3081 37188 3133
rect 37240 3081 37243 3133
rect 37185 3069 37197 3081
rect 37231 3069 37243 3081
rect 37185 3017 37188 3069
rect 37240 3017 37243 3069
rect 37185 3005 37197 3017
rect 37231 3005 37243 3017
rect 37185 2953 37188 3005
rect 37240 2953 37243 3005
rect 37185 2941 37197 2953
rect 37231 2941 37243 2953
rect 37185 2889 37188 2941
rect 37240 2889 37243 2941
rect 37185 2884 37243 2889
rect 37185 2877 37197 2884
rect 37231 2877 37243 2884
rect 37185 2825 37188 2877
rect 37240 2825 37243 2877
rect 37185 2813 37243 2825
rect 37185 2761 37188 2813
rect 37240 2761 37243 2813
rect 37185 2749 37243 2761
rect 37185 2697 37188 2749
rect 37240 2697 37243 2749
rect 37185 2685 37243 2697
rect 37185 2633 37188 2685
rect 37240 2633 37243 2685
rect 37185 2621 37243 2633
rect 37185 2569 37188 2621
rect 37240 2569 37243 2621
rect 37185 2562 37197 2569
rect 37231 2562 37243 2569
rect 37185 2557 37243 2562
rect 37185 2505 37188 2557
rect 37240 2505 37243 2557
rect 37185 2493 37197 2505
rect 37231 2493 37243 2505
rect 37185 2441 37188 2493
rect 37240 2441 37243 2493
rect 37185 2429 37197 2441
rect 37231 2429 37243 2441
rect 37185 2377 37188 2429
rect 37240 2377 37243 2429
rect 37185 2365 37197 2377
rect 37231 2365 37243 2377
rect 37185 2313 37188 2365
rect 37240 2313 37243 2365
rect 37185 2308 37243 2313
rect 37185 2301 37197 2308
rect 37231 2301 37243 2308
rect 37185 2249 37188 2301
rect 37240 2249 37243 2301
rect 37185 2237 37243 2249
rect 37185 2185 37188 2237
rect 37240 2185 37243 2237
rect 37185 2173 37243 2185
rect 37185 2121 37188 2173
rect 37240 2121 37243 2173
rect 37185 2109 37243 2121
rect 37185 2057 37188 2109
rect 37240 2057 37243 2109
rect 37185 2045 37243 2057
rect 37185 1993 37188 2045
rect 37240 1993 37243 2045
rect 37185 1986 37197 1993
rect 37231 1986 37243 1993
rect 37185 1981 37243 1986
rect 37185 1929 37188 1981
rect 37240 1929 37243 1981
rect 37185 1917 37197 1929
rect 37231 1917 37243 1929
rect 37185 1865 37188 1917
rect 37240 1865 37243 1917
rect 37185 1853 37197 1865
rect 37231 1853 37243 1865
rect 37185 1801 37188 1853
rect 37240 1801 37243 1853
rect 37185 1789 37197 1801
rect 37231 1789 37243 1801
rect 37185 1737 37188 1789
rect 37240 1737 37243 1789
rect 37185 1732 37243 1737
rect 37185 1725 37197 1732
rect 37231 1725 37243 1732
rect 37185 1673 37188 1725
rect 37240 1673 37243 1725
rect 37185 1661 37243 1673
rect 37185 1609 37188 1661
rect 37240 1609 37243 1661
rect 37185 1597 37243 1609
rect 37185 1545 37188 1597
rect 37240 1545 37243 1597
rect 37185 1533 37243 1545
rect 37185 1481 37188 1533
rect 37240 1481 37243 1533
rect 37185 1469 37243 1481
rect 37185 1417 37188 1469
rect 37240 1417 37243 1469
rect 37185 1410 37197 1417
rect 37231 1410 37243 1417
rect 37185 1405 37243 1410
rect 37185 1353 37188 1405
rect 37240 1353 37243 1405
rect 37185 1341 37197 1353
rect 37231 1341 37243 1353
rect 37185 1289 37188 1341
rect 37240 1289 37243 1341
rect 37185 1277 37197 1289
rect 37231 1277 37243 1289
rect 37185 1225 37188 1277
rect 37240 1225 37243 1277
rect 37185 1213 37197 1225
rect 37231 1213 37243 1225
rect 37185 1161 37188 1213
rect 37240 1161 37243 1213
rect 37185 1147 37243 1161
rect 37281 3133 37339 3147
rect 37281 3081 37284 3133
rect 37336 3081 37339 3133
rect 37281 3069 37293 3081
rect 37327 3069 37339 3081
rect 37281 3017 37284 3069
rect 37336 3017 37339 3069
rect 37281 3005 37293 3017
rect 37327 3005 37339 3017
rect 37281 2953 37284 3005
rect 37336 2953 37339 3005
rect 37281 2941 37293 2953
rect 37327 2941 37339 2953
rect 37281 2889 37284 2941
rect 37336 2889 37339 2941
rect 37281 2884 37339 2889
rect 37281 2877 37293 2884
rect 37327 2877 37339 2884
rect 37281 2825 37284 2877
rect 37336 2825 37339 2877
rect 37281 2813 37339 2825
rect 37281 2761 37284 2813
rect 37336 2761 37339 2813
rect 37281 2749 37339 2761
rect 37281 2697 37284 2749
rect 37336 2697 37339 2749
rect 37281 2685 37339 2697
rect 37281 2633 37284 2685
rect 37336 2633 37339 2685
rect 37281 2621 37339 2633
rect 37281 2569 37284 2621
rect 37336 2569 37339 2621
rect 37281 2562 37293 2569
rect 37327 2562 37339 2569
rect 37281 2557 37339 2562
rect 37281 2505 37284 2557
rect 37336 2505 37339 2557
rect 37281 2493 37293 2505
rect 37327 2493 37339 2505
rect 37281 2441 37284 2493
rect 37336 2441 37339 2493
rect 37281 2429 37293 2441
rect 37327 2429 37339 2441
rect 37281 2377 37284 2429
rect 37336 2377 37339 2429
rect 37281 2365 37293 2377
rect 37327 2365 37339 2377
rect 37281 2313 37284 2365
rect 37336 2313 37339 2365
rect 37281 2308 37339 2313
rect 37281 2301 37293 2308
rect 37327 2301 37339 2308
rect 37281 2249 37284 2301
rect 37336 2249 37339 2301
rect 37281 2237 37339 2249
rect 37281 2185 37284 2237
rect 37336 2185 37339 2237
rect 37281 2173 37339 2185
rect 37281 2121 37284 2173
rect 37336 2121 37339 2173
rect 37281 2109 37339 2121
rect 37281 2057 37284 2109
rect 37336 2057 37339 2109
rect 37281 2045 37339 2057
rect 37281 1993 37284 2045
rect 37336 1993 37339 2045
rect 37281 1986 37293 1993
rect 37327 1986 37339 1993
rect 37281 1981 37339 1986
rect 37281 1929 37284 1981
rect 37336 1929 37339 1981
rect 37281 1917 37293 1929
rect 37327 1917 37339 1929
rect 37281 1865 37284 1917
rect 37336 1865 37339 1917
rect 37281 1853 37293 1865
rect 37327 1853 37339 1865
rect 37281 1801 37284 1853
rect 37336 1801 37339 1853
rect 37281 1789 37293 1801
rect 37327 1789 37339 1801
rect 37281 1737 37284 1789
rect 37336 1737 37339 1789
rect 37281 1732 37339 1737
rect 37281 1725 37293 1732
rect 37327 1725 37339 1732
rect 37281 1673 37284 1725
rect 37336 1673 37339 1725
rect 37281 1661 37339 1673
rect 37281 1609 37284 1661
rect 37336 1609 37339 1661
rect 37281 1597 37339 1609
rect 37281 1545 37284 1597
rect 37336 1545 37339 1597
rect 37281 1533 37339 1545
rect 37281 1481 37284 1533
rect 37336 1481 37339 1533
rect 37281 1469 37339 1481
rect 37281 1417 37284 1469
rect 37336 1417 37339 1469
rect 37281 1410 37293 1417
rect 37327 1410 37339 1417
rect 37281 1405 37339 1410
rect 37281 1353 37284 1405
rect 37336 1353 37339 1405
rect 37281 1341 37293 1353
rect 37327 1341 37339 1353
rect 37281 1289 37284 1341
rect 37336 1289 37339 1341
rect 37281 1277 37293 1289
rect 37327 1277 37339 1289
rect 37281 1225 37284 1277
rect 37336 1225 37339 1277
rect 37281 1213 37293 1225
rect 37327 1213 37339 1225
rect 37281 1161 37284 1213
rect 37336 1161 37339 1213
rect 37281 1147 37339 1161
rect 37380 3133 37432 3147
rect 37380 3069 37389 3081
rect 37423 3069 37432 3081
rect 37380 3005 37389 3017
rect 37423 3005 37432 3017
rect 37380 2941 37389 2953
rect 37423 2941 37432 2953
rect 37380 2884 37432 2889
rect 37380 2877 37389 2884
rect 37423 2877 37432 2884
rect 37380 2813 37432 2825
rect 37380 2749 37432 2761
rect 37380 2685 37432 2697
rect 37380 2621 37432 2633
rect 37380 2562 37389 2569
rect 37423 2562 37432 2569
rect 37380 2557 37432 2562
rect 37380 2493 37389 2505
rect 37423 2493 37432 2505
rect 37380 2429 37389 2441
rect 37423 2429 37432 2441
rect 37380 2365 37389 2377
rect 37423 2365 37432 2377
rect 37380 2308 37432 2313
rect 37380 2301 37389 2308
rect 37423 2301 37432 2308
rect 37380 2237 37432 2249
rect 37380 2173 37432 2185
rect 37380 2109 37432 2121
rect 37380 2045 37432 2057
rect 37380 1986 37389 1993
rect 37423 1986 37432 1993
rect 37380 1981 37432 1986
rect 37380 1917 37389 1929
rect 37423 1917 37432 1929
rect 37380 1853 37389 1865
rect 37423 1853 37432 1865
rect 37380 1789 37389 1801
rect 37423 1789 37432 1801
rect 37380 1732 37432 1737
rect 37380 1725 37389 1732
rect 37423 1725 37432 1732
rect 37380 1661 37432 1673
rect 37380 1597 37432 1609
rect 37380 1533 37432 1545
rect 37380 1469 37432 1481
rect 37380 1410 37389 1417
rect 37423 1410 37432 1417
rect 37380 1405 37432 1410
rect 37380 1341 37389 1353
rect 37423 1341 37432 1353
rect 37380 1277 37389 1289
rect 37423 1277 37432 1289
rect 37380 1213 37389 1225
rect 37423 1213 37432 1225
rect 37380 1147 37432 1161
rect 37473 3133 37531 3147
rect 37473 3081 37476 3133
rect 37528 3081 37531 3133
rect 37473 3069 37485 3081
rect 37519 3069 37531 3081
rect 37473 3017 37476 3069
rect 37528 3017 37531 3069
rect 37473 3005 37485 3017
rect 37519 3005 37531 3017
rect 37473 2953 37476 3005
rect 37528 2953 37531 3005
rect 37473 2941 37485 2953
rect 37519 2941 37531 2953
rect 37473 2889 37476 2941
rect 37528 2889 37531 2941
rect 37473 2884 37531 2889
rect 37473 2877 37485 2884
rect 37519 2877 37531 2884
rect 37473 2825 37476 2877
rect 37528 2825 37531 2877
rect 37473 2813 37531 2825
rect 37473 2761 37476 2813
rect 37528 2761 37531 2813
rect 37473 2749 37531 2761
rect 37473 2697 37476 2749
rect 37528 2697 37531 2749
rect 37473 2685 37531 2697
rect 37473 2633 37476 2685
rect 37528 2633 37531 2685
rect 37473 2621 37531 2633
rect 37473 2569 37476 2621
rect 37528 2569 37531 2621
rect 37473 2562 37485 2569
rect 37519 2562 37531 2569
rect 37473 2557 37531 2562
rect 37473 2505 37476 2557
rect 37528 2505 37531 2557
rect 37473 2493 37485 2505
rect 37519 2493 37531 2505
rect 37473 2441 37476 2493
rect 37528 2441 37531 2493
rect 37473 2429 37485 2441
rect 37519 2429 37531 2441
rect 37473 2377 37476 2429
rect 37528 2377 37531 2429
rect 37473 2365 37485 2377
rect 37519 2365 37531 2377
rect 37473 2313 37476 2365
rect 37528 2313 37531 2365
rect 37473 2308 37531 2313
rect 37473 2301 37485 2308
rect 37519 2301 37531 2308
rect 37473 2249 37476 2301
rect 37528 2249 37531 2301
rect 37473 2237 37531 2249
rect 37473 2185 37476 2237
rect 37528 2185 37531 2237
rect 37473 2173 37531 2185
rect 37473 2121 37476 2173
rect 37528 2121 37531 2173
rect 37473 2109 37531 2121
rect 37473 2057 37476 2109
rect 37528 2057 37531 2109
rect 37473 2045 37531 2057
rect 37473 1993 37476 2045
rect 37528 1993 37531 2045
rect 37473 1986 37485 1993
rect 37519 1986 37531 1993
rect 37473 1981 37531 1986
rect 37473 1929 37476 1981
rect 37528 1929 37531 1981
rect 37473 1917 37485 1929
rect 37519 1917 37531 1929
rect 37473 1865 37476 1917
rect 37528 1865 37531 1917
rect 37473 1853 37485 1865
rect 37519 1853 37531 1865
rect 37473 1801 37476 1853
rect 37528 1801 37531 1853
rect 37473 1789 37485 1801
rect 37519 1789 37531 1801
rect 37473 1737 37476 1789
rect 37528 1737 37531 1789
rect 37473 1732 37531 1737
rect 37473 1725 37485 1732
rect 37519 1725 37531 1732
rect 37473 1673 37476 1725
rect 37528 1673 37531 1725
rect 37473 1661 37531 1673
rect 37473 1609 37476 1661
rect 37528 1609 37531 1661
rect 37473 1597 37531 1609
rect 37473 1545 37476 1597
rect 37528 1545 37531 1597
rect 37473 1533 37531 1545
rect 37473 1481 37476 1533
rect 37528 1481 37531 1533
rect 37473 1469 37531 1481
rect 37473 1417 37476 1469
rect 37528 1417 37531 1469
rect 37473 1410 37485 1417
rect 37519 1410 37531 1417
rect 37473 1405 37531 1410
rect 37473 1353 37476 1405
rect 37528 1353 37531 1405
rect 37473 1341 37485 1353
rect 37519 1341 37531 1353
rect 37473 1289 37476 1341
rect 37528 1289 37531 1341
rect 37473 1277 37485 1289
rect 37519 1277 37531 1289
rect 37473 1225 37476 1277
rect 37528 1225 37531 1277
rect 37473 1213 37485 1225
rect 37519 1213 37531 1225
rect 37473 1161 37476 1213
rect 37528 1161 37531 1213
rect 37473 1147 37531 1161
rect 37569 3133 37627 3147
rect 37569 3081 37572 3133
rect 37624 3081 37627 3133
rect 37569 3069 37581 3081
rect 37615 3069 37627 3081
rect 37569 3017 37572 3069
rect 37624 3017 37627 3069
rect 37569 3005 37581 3017
rect 37615 3005 37627 3017
rect 37569 2953 37572 3005
rect 37624 2953 37627 3005
rect 37569 2941 37581 2953
rect 37615 2941 37627 2953
rect 37569 2889 37572 2941
rect 37624 2889 37627 2941
rect 37569 2884 37627 2889
rect 37569 2877 37581 2884
rect 37615 2877 37627 2884
rect 37569 2825 37572 2877
rect 37624 2825 37627 2877
rect 37569 2813 37627 2825
rect 37569 2761 37572 2813
rect 37624 2761 37627 2813
rect 37569 2749 37627 2761
rect 37569 2697 37572 2749
rect 37624 2697 37627 2749
rect 37569 2685 37627 2697
rect 37569 2633 37572 2685
rect 37624 2633 37627 2685
rect 37569 2621 37627 2633
rect 37569 2569 37572 2621
rect 37624 2569 37627 2621
rect 37569 2562 37581 2569
rect 37615 2562 37627 2569
rect 37569 2557 37627 2562
rect 37569 2505 37572 2557
rect 37624 2505 37627 2557
rect 37569 2493 37581 2505
rect 37615 2493 37627 2505
rect 37569 2441 37572 2493
rect 37624 2441 37627 2493
rect 37569 2429 37581 2441
rect 37615 2429 37627 2441
rect 37569 2377 37572 2429
rect 37624 2377 37627 2429
rect 37569 2365 37581 2377
rect 37615 2365 37627 2377
rect 37569 2313 37572 2365
rect 37624 2313 37627 2365
rect 37569 2308 37627 2313
rect 37569 2301 37581 2308
rect 37615 2301 37627 2308
rect 37569 2249 37572 2301
rect 37624 2249 37627 2301
rect 37569 2237 37627 2249
rect 37569 2185 37572 2237
rect 37624 2185 37627 2237
rect 37569 2173 37627 2185
rect 37569 2121 37572 2173
rect 37624 2121 37627 2173
rect 37569 2109 37627 2121
rect 37569 2057 37572 2109
rect 37624 2057 37627 2109
rect 37569 2045 37627 2057
rect 37569 1993 37572 2045
rect 37624 1993 37627 2045
rect 37569 1986 37581 1993
rect 37615 1986 37627 1993
rect 37569 1981 37627 1986
rect 37569 1929 37572 1981
rect 37624 1929 37627 1981
rect 37569 1917 37581 1929
rect 37615 1917 37627 1929
rect 37569 1865 37572 1917
rect 37624 1865 37627 1917
rect 37569 1853 37581 1865
rect 37615 1853 37627 1865
rect 37569 1801 37572 1853
rect 37624 1801 37627 1853
rect 37569 1789 37581 1801
rect 37615 1789 37627 1801
rect 37569 1737 37572 1789
rect 37624 1737 37627 1789
rect 37569 1732 37627 1737
rect 37569 1725 37581 1732
rect 37615 1725 37627 1732
rect 37569 1673 37572 1725
rect 37624 1673 37627 1725
rect 37569 1661 37627 1673
rect 37569 1609 37572 1661
rect 37624 1609 37627 1661
rect 37569 1597 37627 1609
rect 37569 1545 37572 1597
rect 37624 1545 37627 1597
rect 37569 1533 37627 1545
rect 37569 1481 37572 1533
rect 37624 1481 37627 1533
rect 37569 1469 37627 1481
rect 37569 1417 37572 1469
rect 37624 1417 37627 1469
rect 37569 1410 37581 1417
rect 37615 1410 37627 1417
rect 37569 1405 37627 1410
rect 37569 1353 37572 1405
rect 37624 1353 37627 1405
rect 37569 1341 37581 1353
rect 37615 1341 37627 1353
rect 37569 1289 37572 1341
rect 37624 1289 37627 1341
rect 37569 1277 37581 1289
rect 37615 1277 37627 1289
rect 37569 1225 37572 1277
rect 37624 1225 37627 1277
rect 37569 1213 37581 1225
rect 37615 1213 37627 1225
rect 37569 1161 37572 1213
rect 37624 1161 37627 1213
rect 37569 1147 37627 1161
rect 37665 3133 37723 3147
rect 37665 3081 37668 3133
rect 37720 3081 37723 3133
rect 37665 3069 37677 3081
rect 37711 3069 37723 3081
rect 37665 3017 37668 3069
rect 37720 3017 37723 3069
rect 37665 3005 37677 3017
rect 37711 3005 37723 3017
rect 37665 2953 37668 3005
rect 37720 2953 37723 3005
rect 37665 2941 37677 2953
rect 37711 2941 37723 2953
rect 37665 2889 37668 2941
rect 37720 2889 37723 2941
rect 37665 2884 37723 2889
rect 37665 2877 37677 2884
rect 37711 2877 37723 2884
rect 37665 2825 37668 2877
rect 37720 2825 37723 2877
rect 37665 2813 37723 2825
rect 37665 2761 37668 2813
rect 37720 2761 37723 2813
rect 37665 2749 37723 2761
rect 37665 2697 37668 2749
rect 37720 2697 37723 2749
rect 37665 2685 37723 2697
rect 37665 2633 37668 2685
rect 37720 2633 37723 2685
rect 37665 2621 37723 2633
rect 37665 2569 37668 2621
rect 37720 2569 37723 2621
rect 37665 2562 37677 2569
rect 37711 2562 37723 2569
rect 37665 2557 37723 2562
rect 37665 2505 37668 2557
rect 37720 2505 37723 2557
rect 37665 2493 37677 2505
rect 37711 2493 37723 2505
rect 37665 2441 37668 2493
rect 37720 2441 37723 2493
rect 37665 2429 37677 2441
rect 37711 2429 37723 2441
rect 37665 2377 37668 2429
rect 37720 2377 37723 2429
rect 37665 2365 37677 2377
rect 37711 2365 37723 2377
rect 37665 2313 37668 2365
rect 37720 2313 37723 2365
rect 37665 2308 37723 2313
rect 37665 2301 37677 2308
rect 37711 2301 37723 2308
rect 37665 2249 37668 2301
rect 37720 2249 37723 2301
rect 37665 2237 37723 2249
rect 37665 2185 37668 2237
rect 37720 2185 37723 2237
rect 37665 2173 37723 2185
rect 37665 2121 37668 2173
rect 37720 2121 37723 2173
rect 37665 2109 37723 2121
rect 37665 2057 37668 2109
rect 37720 2057 37723 2109
rect 37665 2045 37723 2057
rect 37665 1993 37668 2045
rect 37720 1993 37723 2045
rect 37665 1986 37677 1993
rect 37711 1986 37723 1993
rect 37665 1981 37723 1986
rect 37665 1929 37668 1981
rect 37720 1929 37723 1981
rect 37665 1917 37677 1929
rect 37711 1917 37723 1929
rect 37665 1865 37668 1917
rect 37720 1865 37723 1917
rect 37665 1853 37677 1865
rect 37711 1853 37723 1865
rect 37665 1801 37668 1853
rect 37720 1801 37723 1853
rect 37665 1789 37677 1801
rect 37711 1789 37723 1801
rect 37665 1737 37668 1789
rect 37720 1737 37723 1789
rect 37665 1732 37723 1737
rect 37665 1725 37677 1732
rect 37711 1725 37723 1732
rect 37665 1673 37668 1725
rect 37720 1673 37723 1725
rect 37665 1661 37723 1673
rect 37665 1609 37668 1661
rect 37720 1609 37723 1661
rect 37665 1597 37723 1609
rect 37665 1545 37668 1597
rect 37720 1545 37723 1597
rect 37665 1533 37723 1545
rect 37665 1481 37668 1533
rect 37720 1481 37723 1533
rect 37665 1469 37723 1481
rect 37665 1417 37668 1469
rect 37720 1417 37723 1469
rect 37665 1410 37677 1417
rect 37711 1410 37723 1417
rect 37665 1405 37723 1410
rect 37665 1353 37668 1405
rect 37720 1353 37723 1405
rect 37665 1341 37677 1353
rect 37711 1341 37723 1353
rect 37665 1289 37668 1341
rect 37720 1289 37723 1341
rect 37665 1277 37677 1289
rect 37711 1277 37723 1289
rect 37665 1225 37668 1277
rect 37720 1225 37723 1277
rect 37665 1213 37677 1225
rect 37711 1213 37723 1225
rect 37665 1161 37668 1213
rect 37720 1161 37723 1213
rect 37665 1147 37723 1161
rect 37764 3133 37816 3147
rect 37764 3069 37773 3081
rect 37807 3069 37816 3081
rect 37764 3005 37773 3017
rect 37807 3005 37816 3017
rect 37764 2941 37773 2953
rect 37807 2941 37816 2953
rect 37764 2884 37816 2889
rect 37764 2877 37773 2884
rect 37807 2877 37816 2884
rect 37764 2813 37816 2825
rect 37764 2749 37816 2761
rect 37764 2685 37816 2697
rect 37764 2621 37816 2633
rect 37764 2562 37773 2569
rect 37807 2562 37816 2569
rect 37764 2557 37816 2562
rect 37764 2493 37773 2505
rect 37807 2493 37816 2505
rect 37764 2429 37773 2441
rect 37807 2429 37816 2441
rect 37764 2365 37773 2377
rect 37807 2365 37816 2377
rect 37764 2308 37816 2313
rect 37764 2301 37773 2308
rect 37807 2301 37816 2308
rect 37764 2237 37816 2249
rect 37764 2173 37816 2185
rect 37764 2109 37816 2121
rect 37764 2045 37816 2057
rect 37764 1986 37773 1993
rect 37807 1986 37816 1993
rect 37764 1981 37816 1986
rect 37764 1917 37773 1929
rect 37807 1917 37816 1929
rect 37764 1853 37773 1865
rect 37807 1853 37816 1865
rect 37764 1789 37773 1801
rect 37807 1789 37816 1801
rect 37764 1732 37816 1737
rect 37764 1725 37773 1732
rect 37807 1725 37816 1732
rect 37764 1661 37816 1673
rect 37764 1597 37816 1609
rect 37764 1533 37816 1545
rect 37764 1469 37816 1481
rect 37764 1410 37773 1417
rect 37807 1410 37816 1417
rect 37764 1405 37816 1410
rect 37764 1341 37773 1353
rect 37807 1341 37816 1353
rect 37764 1277 37773 1289
rect 37807 1277 37816 1289
rect 37764 1213 37773 1225
rect 37807 1213 37816 1225
rect 37764 1147 37816 1161
rect 37857 3133 37915 3147
rect 37857 3081 37860 3133
rect 37912 3081 37915 3133
rect 37857 3069 37869 3081
rect 37903 3069 37915 3081
rect 37857 3017 37860 3069
rect 37912 3017 37915 3069
rect 37857 3005 37869 3017
rect 37903 3005 37915 3017
rect 37857 2953 37860 3005
rect 37912 2953 37915 3005
rect 37857 2941 37869 2953
rect 37903 2941 37915 2953
rect 37857 2889 37860 2941
rect 37912 2889 37915 2941
rect 37857 2884 37915 2889
rect 37857 2877 37869 2884
rect 37903 2877 37915 2884
rect 37857 2825 37860 2877
rect 37912 2825 37915 2877
rect 37857 2813 37915 2825
rect 37857 2761 37860 2813
rect 37912 2761 37915 2813
rect 37857 2749 37915 2761
rect 37857 2697 37860 2749
rect 37912 2697 37915 2749
rect 37857 2685 37915 2697
rect 37857 2633 37860 2685
rect 37912 2633 37915 2685
rect 37857 2621 37915 2633
rect 37857 2569 37860 2621
rect 37912 2569 37915 2621
rect 37857 2562 37869 2569
rect 37903 2562 37915 2569
rect 37857 2557 37915 2562
rect 37857 2505 37860 2557
rect 37912 2505 37915 2557
rect 37857 2493 37869 2505
rect 37903 2493 37915 2505
rect 37857 2441 37860 2493
rect 37912 2441 37915 2493
rect 37857 2429 37869 2441
rect 37903 2429 37915 2441
rect 37857 2377 37860 2429
rect 37912 2377 37915 2429
rect 37857 2365 37869 2377
rect 37903 2365 37915 2377
rect 37857 2313 37860 2365
rect 37912 2313 37915 2365
rect 37857 2308 37915 2313
rect 37857 2301 37869 2308
rect 37903 2301 37915 2308
rect 37857 2249 37860 2301
rect 37912 2249 37915 2301
rect 37857 2237 37915 2249
rect 37857 2185 37860 2237
rect 37912 2185 37915 2237
rect 37857 2173 37915 2185
rect 37857 2121 37860 2173
rect 37912 2121 37915 2173
rect 37857 2109 37915 2121
rect 37857 2057 37860 2109
rect 37912 2057 37915 2109
rect 37857 2045 37915 2057
rect 37857 1993 37860 2045
rect 37912 1993 37915 2045
rect 37857 1986 37869 1993
rect 37903 1986 37915 1993
rect 37857 1981 37915 1986
rect 37857 1929 37860 1981
rect 37912 1929 37915 1981
rect 37857 1917 37869 1929
rect 37903 1917 37915 1929
rect 37857 1865 37860 1917
rect 37912 1865 37915 1917
rect 37857 1853 37869 1865
rect 37903 1853 37915 1865
rect 37857 1801 37860 1853
rect 37912 1801 37915 1853
rect 37857 1789 37869 1801
rect 37903 1789 37915 1801
rect 37857 1737 37860 1789
rect 37912 1737 37915 1789
rect 37857 1732 37915 1737
rect 37857 1725 37869 1732
rect 37903 1725 37915 1732
rect 37857 1673 37860 1725
rect 37912 1673 37915 1725
rect 37857 1661 37915 1673
rect 37857 1609 37860 1661
rect 37912 1609 37915 1661
rect 37857 1597 37915 1609
rect 37857 1545 37860 1597
rect 37912 1545 37915 1597
rect 37857 1533 37915 1545
rect 37857 1481 37860 1533
rect 37912 1481 37915 1533
rect 37857 1469 37915 1481
rect 37857 1417 37860 1469
rect 37912 1417 37915 1469
rect 37857 1410 37869 1417
rect 37903 1410 37915 1417
rect 37857 1405 37915 1410
rect 37857 1353 37860 1405
rect 37912 1353 37915 1405
rect 37857 1341 37869 1353
rect 37903 1341 37915 1353
rect 37857 1289 37860 1341
rect 37912 1289 37915 1341
rect 37857 1277 37869 1289
rect 37903 1277 37915 1289
rect 37857 1225 37860 1277
rect 37912 1225 37915 1277
rect 37857 1213 37869 1225
rect 37903 1213 37915 1225
rect 37857 1161 37860 1213
rect 37912 1161 37915 1213
rect 37857 1147 37915 1161
rect 37953 3133 38011 3147
rect 37953 3081 37956 3133
rect 38008 3081 38011 3133
rect 37953 3069 37965 3081
rect 37999 3069 38011 3081
rect 37953 3017 37956 3069
rect 38008 3017 38011 3069
rect 37953 3005 37965 3017
rect 37999 3005 38011 3017
rect 37953 2953 37956 3005
rect 38008 2953 38011 3005
rect 37953 2941 37965 2953
rect 37999 2941 38011 2953
rect 37953 2889 37956 2941
rect 38008 2889 38011 2941
rect 37953 2884 38011 2889
rect 37953 2877 37965 2884
rect 37999 2877 38011 2884
rect 37953 2825 37956 2877
rect 38008 2825 38011 2877
rect 37953 2813 38011 2825
rect 37953 2761 37956 2813
rect 38008 2761 38011 2813
rect 37953 2749 38011 2761
rect 37953 2697 37956 2749
rect 38008 2697 38011 2749
rect 37953 2685 38011 2697
rect 37953 2633 37956 2685
rect 38008 2633 38011 2685
rect 37953 2621 38011 2633
rect 37953 2569 37956 2621
rect 38008 2569 38011 2621
rect 37953 2562 37965 2569
rect 37999 2562 38011 2569
rect 37953 2557 38011 2562
rect 37953 2505 37956 2557
rect 38008 2505 38011 2557
rect 37953 2493 37965 2505
rect 37999 2493 38011 2505
rect 37953 2441 37956 2493
rect 38008 2441 38011 2493
rect 37953 2429 37965 2441
rect 37999 2429 38011 2441
rect 37953 2377 37956 2429
rect 38008 2377 38011 2429
rect 37953 2365 37965 2377
rect 37999 2365 38011 2377
rect 37953 2313 37956 2365
rect 38008 2313 38011 2365
rect 37953 2308 38011 2313
rect 37953 2301 37965 2308
rect 37999 2301 38011 2308
rect 37953 2249 37956 2301
rect 38008 2249 38011 2301
rect 37953 2237 38011 2249
rect 37953 2185 37956 2237
rect 38008 2185 38011 2237
rect 37953 2173 38011 2185
rect 37953 2121 37956 2173
rect 38008 2121 38011 2173
rect 37953 2109 38011 2121
rect 37953 2057 37956 2109
rect 38008 2057 38011 2109
rect 37953 2045 38011 2057
rect 37953 1993 37956 2045
rect 38008 1993 38011 2045
rect 37953 1986 37965 1993
rect 37999 1986 38011 1993
rect 37953 1981 38011 1986
rect 37953 1929 37956 1981
rect 38008 1929 38011 1981
rect 37953 1917 37965 1929
rect 37999 1917 38011 1929
rect 37953 1865 37956 1917
rect 38008 1865 38011 1917
rect 37953 1853 37965 1865
rect 37999 1853 38011 1865
rect 37953 1801 37956 1853
rect 38008 1801 38011 1853
rect 37953 1789 37965 1801
rect 37999 1789 38011 1801
rect 37953 1737 37956 1789
rect 38008 1737 38011 1789
rect 37953 1732 38011 1737
rect 37953 1725 37965 1732
rect 37999 1725 38011 1732
rect 37953 1673 37956 1725
rect 38008 1673 38011 1725
rect 37953 1661 38011 1673
rect 37953 1609 37956 1661
rect 38008 1609 38011 1661
rect 37953 1597 38011 1609
rect 37953 1545 37956 1597
rect 38008 1545 38011 1597
rect 37953 1533 38011 1545
rect 37953 1481 37956 1533
rect 38008 1481 38011 1533
rect 37953 1469 38011 1481
rect 37953 1417 37956 1469
rect 38008 1417 38011 1469
rect 37953 1410 37965 1417
rect 37999 1410 38011 1417
rect 37953 1405 38011 1410
rect 37953 1353 37956 1405
rect 38008 1353 38011 1405
rect 37953 1341 37965 1353
rect 37999 1341 38011 1353
rect 37953 1289 37956 1341
rect 38008 1289 38011 1341
rect 37953 1277 37965 1289
rect 37999 1277 38011 1289
rect 37953 1225 37956 1277
rect 38008 1225 38011 1277
rect 37953 1213 37965 1225
rect 37999 1213 38011 1225
rect 37953 1161 37956 1213
rect 38008 1161 38011 1213
rect 37953 1147 38011 1161
rect 38049 3133 38107 3147
rect 38049 3081 38052 3133
rect 38104 3081 38107 3133
rect 38049 3069 38061 3081
rect 38095 3069 38107 3081
rect 38049 3017 38052 3069
rect 38104 3017 38107 3069
rect 38049 3005 38061 3017
rect 38095 3005 38107 3017
rect 38049 2953 38052 3005
rect 38104 2953 38107 3005
rect 38049 2941 38061 2953
rect 38095 2941 38107 2953
rect 38049 2889 38052 2941
rect 38104 2889 38107 2941
rect 38049 2884 38107 2889
rect 38049 2877 38061 2884
rect 38095 2877 38107 2884
rect 38049 2825 38052 2877
rect 38104 2825 38107 2877
rect 38049 2813 38107 2825
rect 38049 2761 38052 2813
rect 38104 2761 38107 2813
rect 38049 2749 38107 2761
rect 38049 2697 38052 2749
rect 38104 2697 38107 2749
rect 38049 2685 38107 2697
rect 38049 2633 38052 2685
rect 38104 2633 38107 2685
rect 38049 2621 38107 2633
rect 38049 2569 38052 2621
rect 38104 2569 38107 2621
rect 38049 2562 38061 2569
rect 38095 2562 38107 2569
rect 38049 2557 38107 2562
rect 38049 2505 38052 2557
rect 38104 2505 38107 2557
rect 38049 2493 38061 2505
rect 38095 2493 38107 2505
rect 38049 2441 38052 2493
rect 38104 2441 38107 2493
rect 38049 2429 38061 2441
rect 38095 2429 38107 2441
rect 38049 2377 38052 2429
rect 38104 2377 38107 2429
rect 38049 2365 38061 2377
rect 38095 2365 38107 2377
rect 38049 2313 38052 2365
rect 38104 2313 38107 2365
rect 38049 2308 38107 2313
rect 38049 2301 38061 2308
rect 38095 2301 38107 2308
rect 38049 2249 38052 2301
rect 38104 2249 38107 2301
rect 38049 2237 38107 2249
rect 38049 2185 38052 2237
rect 38104 2185 38107 2237
rect 38049 2173 38107 2185
rect 38049 2121 38052 2173
rect 38104 2121 38107 2173
rect 38049 2109 38107 2121
rect 38049 2057 38052 2109
rect 38104 2057 38107 2109
rect 38049 2045 38107 2057
rect 38049 1993 38052 2045
rect 38104 1993 38107 2045
rect 38049 1986 38061 1993
rect 38095 1986 38107 1993
rect 38049 1981 38107 1986
rect 38049 1929 38052 1981
rect 38104 1929 38107 1981
rect 38049 1917 38061 1929
rect 38095 1917 38107 1929
rect 38049 1865 38052 1917
rect 38104 1865 38107 1917
rect 38049 1853 38061 1865
rect 38095 1853 38107 1865
rect 38049 1801 38052 1853
rect 38104 1801 38107 1853
rect 38049 1789 38061 1801
rect 38095 1789 38107 1801
rect 38049 1737 38052 1789
rect 38104 1737 38107 1789
rect 38049 1732 38107 1737
rect 38049 1725 38061 1732
rect 38095 1725 38107 1732
rect 38049 1673 38052 1725
rect 38104 1673 38107 1725
rect 38049 1661 38107 1673
rect 38049 1609 38052 1661
rect 38104 1609 38107 1661
rect 38049 1597 38107 1609
rect 38049 1545 38052 1597
rect 38104 1545 38107 1597
rect 38049 1533 38107 1545
rect 38049 1481 38052 1533
rect 38104 1481 38107 1533
rect 38049 1469 38107 1481
rect 38049 1417 38052 1469
rect 38104 1417 38107 1469
rect 38049 1410 38061 1417
rect 38095 1410 38107 1417
rect 38049 1405 38107 1410
rect 38049 1353 38052 1405
rect 38104 1353 38107 1405
rect 38049 1341 38061 1353
rect 38095 1341 38107 1353
rect 38049 1289 38052 1341
rect 38104 1289 38107 1341
rect 38049 1277 38061 1289
rect 38095 1277 38107 1289
rect 38049 1225 38052 1277
rect 38104 1225 38107 1277
rect 38049 1213 38061 1225
rect 38095 1213 38107 1225
rect 38049 1161 38052 1213
rect 38104 1161 38107 1213
rect 38049 1147 38107 1161
rect 38148 3133 38200 3147
rect 38148 3069 38157 3081
rect 38191 3069 38200 3081
rect 38148 3005 38157 3017
rect 38191 3005 38200 3017
rect 38148 2941 38157 2953
rect 38191 2941 38200 2953
rect 38148 2884 38200 2889
rect 38148 2877 38157 2884
rect 38191 2877 38200 2884
rect 38148 2813 38200 2825
rect 38148 2749 38200 2761
rect 38148 2685 38200 2697
rect 38148 2621 38200 2633
rect 38148 2562 38157 2569
rect 38191 2562 38200 2569
rect 38148 2557 38200 2562
rect 38148 2493 38157 2505
rect 38191 2493 38200 2505
rect 38148 2429 38157 2441
rect 38191 2429 38200 2441
rect 38148 2365 38157 2377
rect 38191 2365 38200 2377
rect 38148 2308 38200 2313
rect 38148 2301 38157 2308
rect 38191 2301 38200 2308
rect 38148 2237 38200 2249
rect 38148 2173 38200 2185
rect 38148 2109 38200 2121
rect 38148 2045 38200 2057
rect 38148 1986 38157 1993
rect 38191 1986 38200 1993
rect 38148 1981 38200 1986
rect 38148 1917 38157 1929
rect 38191 1917 38200 1929
rect 38148 1853 38157 1865
rect 38191 1853 38200 1865
rect 38148 1789 38157 1801
rect 38191 1789 38200 1801
rect 38148 1732 38200 1737
rect 38148 1725 38157 1732
rect 38191 1725 38200 1732
rect 38148 1661 38200 1673
rect 38148 1597 38200 1609
rect 38148 1533 38200 1545
rect 38148 1469 38200 1481
rect 38148 1410 38157 1417
rect 38191 1410 38200 1417
rect 38148 1405 38200 1410
rect 38148 1341 38157 1353
rect 38191 1341 38200 1353
rect 38148 1277 38157 1289
rect 38191 1277 38200 1289
rect 38148 1213 38157 1225
rect 38191 1213 38200 1225
rect 38148 1147 38200 1161
rect 38241 3133 38299 3147
rect 38241 3081 38244 3133
rect 38296 3081 38299 3133
rect 38241 3069 38253 3081
rect 38287 3069 38299 3081
rect 38241 3017 38244 3069
rect 38296 3017 38299 3069
rect 38241 3005 38253 3017
rect 38287 3005 38299 3017
rect 38241 2953 38244 3005
rect 38296 2953 38299 3005
rect 38241 2941 38253 2953
rect 38287 2941 38299 2953
rect 38241 2889 38244 2941
rect 38296 2889 38299 2941
rect 38241 2884 38299 2889
rect 38241 2877 38253 2884
rect 38287 2877 38299 2884
rect 38241 2825 38244 2877
rect 38296 2825 38299 2877
rect 38241 2813 38299 2825
rect 38241 2761 38244 2813
rect 38296 2761 38299 2813
rect 38241 2749 38299 2761
rect 38241 2697 38244 2749
rect 38296 2697 38299 2749
rect 38241 2685 38299 2697
rect 38241 2633 38244 2685
rect 38296 2633 38299 2685
rect 38241 2621 38299 2633
rect 38241 2569 38244 2621
rect 38296 2569 38299 2621
rect 38241 2562 38253 2569
rect 38287 2562 38299 2569
rect 38241 2557 38299 2562
rect 38241 2505 38244 2557
rect 38296 2505 38299 2557
rect 38241 2493 38253 2505
rect 38287 2493 38299 2505
rect 38241 2441 38244 2493
rect 38296 2441 38299 2493
rect 38241 2429 38253 2441
rect 38287 2429 38299 2441
rect 38241 2377 38244 2429
rect 38296 2377 38299 2429
rect 38241 2365 38253 2377
rect 38287 2365 38299 2377
rect 38241 2313 38244 2365
rect 38296 2313 38299 2365
rect 38241 2308 38299 2313
rect 38241 2301 38253 2308
rect 38287 2301 38299 2308
rect 38241 2249 38244 2301
rect 38296 2249 38299 2301
rect 38241 2237 38299 2249
rect 38241 2185 38244 2237
rect 38296 2185 38299 2237
rect 38241 2173 38299 2185
rect 38241 2121 38244 2173
rect 38296 2121 38299 2173
rect 38241 2109 38299 2121
rect 38241 2057 38244 2109
rect 38296 2057 38299 2109
rect 38241 2045 38299 2057
rect 38241 1993 38244 2045
rect 38296 1993 38299 2045
rect 38241 1986 38253 1993
rect 38287 1986 38299 1993
rect 38241 1981 38299 1986
rect 38241 1929 38244 1981
rect 38296 1929 38299 1981
rect 38241 1917 38253 1929
rect 38287 1917 38299 1929
rect 38241 1865 38244 1917
rect 38296 1865 38299 1917
rect 38241 1853 38253 1865
rect 38287 1853 38299 1865
rect 38241 1801 38244 1853
rect 38296 1801 38299 1853
rect 38241 1789 38253 1801
rect 38287 1789 38299 1801
rect 38241 1737 38244 1789
rect 38296 1737 38299 1789
rect 38241 1732 38299 1737
rect 38241 1725 38253 1732
rect 38287 1725 38299 1732
rect 38241 1673 38244 1725
rect 38296 1673 38299 1725
rect 38241 1661 38299 1673
rect 38241 1609 38244 1661
rect 38296 1609 38299 1661
rect 38241 1597 38299 1609
rect 38241 1545 38244 1597
rect 38296 1545 38299 1597
rect 38241 1533 38299 1545
rect 38241 1481 38244 1533
rect 38296 1481 38299 1533
rect 38241 1469 38299 1481
rect 38241 1417 38244 1469
rect 38296 1417 38299 1469
rect 38241 1410 38253 1417
rect 38287 1410 38299 1417
rect 38241 1405 38299 1410
rect 38241 1353 38244 1405
rect 38296 1353 38299 1405
rect 38241 1341 38253 1353
rect 38287 1341 38299 1353
rect 38241 1289 38244 1341
rect 38296 1289 38299 1341
rect 38241 1277 38253 1289
rect 38287 1277 38299 1289
rect 38241 1225 38244 1277
rect 38296 1225 38299 1277
rect 38241 1213 38253 1225
rect 38287 1213 38299 1225
rect 38241 1161 38244 1213
rect 38296 1161 38299 1213
rect 38241 1147 38299 1161
rect 38337 3133 38395 3147
rect 38337 3081 38340 3133
rect 38392 3081 38395 3133
rect 38337 3069 38349 3081
rect 38383 3069 38395 3081
rect 38337 3017 38340 3069
rect 38392 3017 38395 3069
rect 38337 3005 38349 3017
rect 38383 3005 38395 3017
rect 38337 2953 38340 3005
rect 38392 2953 38395 3005
rect 38337 2941 38349 2953
rect 38383 2941 38395 2953
rect 38337 2889 38340 2941
rect 38392 2889 38395 2941
rect 38337 2884 38395 2889
rect 38337 2877 38349 2884
rect 38383 2877 38395 2884
rect 38337 2825 38340 2877
rect 38392 2825 38395 2877
rect 38337 2813 38395 2825
rect 38337 2761 38340 2813
rect 38392 2761 38395 2813
rect 38337 2749 38395 2761
rect 38337 2697 38340 2749
rect 38392 2697 38395 2749
rect 38337 2685 38395 2697
rect 38337 2633 38340 2685
rect 38392 2633 38395 2685
rect 38337 2621 38395 2633
rect 38337 2569 38340 2621
rect 38392 2569 38395 2621
rect 38337 2562 38349 2569
rect 38383 2562 38395 2569
rect 38337 2557 38395 2562
rect 38337 2505 38340 2557
rect 38392 2505 38395 2557
rect 38337 2493 38349 2505
rect 38383 2493 38395 2505
rect 38337 2441 38340 2493
rect 38392 2441 38395 2493
rect 38337 2429 38349 2441
rect 38383 2429 38395 2441
rect 38337 2377 38340 2429
rect 38392 2377 38395 2429
rect 38337 2365 38349 2377
rect 38383 2365 38395 2377
rect 38337 2313 38340 2365
rect 38392 2313 38395 2365
rect 38337 2308 38395 2313
rect 38337 2301 38349 2308
rect 38383 2301 38395 2308
rect 38337 2249 38340 2301
rect 38392 2249 38395 2301
rect 38337 2237 38395 2249
rect 38337 2185 38340 2237
rect 38392 2185 38395 2237
rect 38337 2173 38395 2185
rect 38337 2121 38340 2173
rect 38392 2121 38395 2173
rect 38337 2109 38395 2121
rect 38337 2057 38340 2109
rect 38392 2057 38395 2109
rect 38337 2045 38395 2057
rect 38337 1993 38340 2045
rect 38392 1993 38395 2045
rect 38337 1986 38349 1993
rect 38383 1986 38395 1993
rect 38337 1981 38395 1986
rect 38337 1929 38340 1981
rect 38392 1929 38395 1981
rect 38337 1917 38349 1929
rect 38383 1917 38395 1929
rect 38337 1865 38340 1917
rect 38392 1865 38395 1917
rect 38337 1853 38349 1865
rect 38383 1853 38395 1865
rect 38337 1801 38340 1853
rect 38392 1801 38395 1853
rect 38337 1789 38349 1801
rect 38383 1789 38395 1801
rect 38337 1737 38340 1789
rect 38392 1737 38395 1789
rect 38337 1732 38395 1737
rect 38337 1725 38349 1732
rect 38383 1725 38395 1732
rect 38337 1673 38340 1725
rect 38392 1673 38395 1725
rect 38337 1661 38395 1673
rect 38337 1609 38340 1661
rect 38392 1609 38395 1661
rect 38337 1597 38395 1609
rect 38337 1545 38340 1597
rect 38392 1545 38395 1597
rect 38337 1533 38395 1545
rect 38337 1481 38340 1533
rect 38392 1481 38395 1533
rect 38337 1469 38395 1481
rect 38337 1417 38340 1469
rect 38392 1417 38395 1469
rect 38337 1410 38349 1417
rect 38383 1410 38395 1417
rect 38337 1405 38395 1410
rect 38337 1353 38340 1405
rect 38392 1353 38395 1405
rect 38337 1341 38349 1353
rect 38383 1341 38395 1353
rect 38337 1289 38340 1341
rect 38392 1289 38395 1341
rect 38337 1277 38349 1289
rect 38383 1277 38395 1289
rect 38337 1225 38340 1277
rect 38392 1225 38395 1277
rect 38337 1213 38349 1225
rect 38383 1213 38395 1225
rect 38337 1161 38340 1213
rect 38392 1161 38395 1213
rect 38337 1147 38395 1161
rect 38433 3133 38491 3147
rect 38433 3081 38436 3133
rect 38488 3081 38491 3133
rect 38433 3069 38445 3081
rect 38479 3069 38491 3081
rect 38433 3017 38436 3069
rect 38488 3017 38491 3069
rect 38433 3005 38445 3017
rect 38479 3005 38491 3017
rect 38433 2953 38436 3005
rect 38488 2953 38491 3005
rect 38433 2941 38445 2953
rect 38479 2941 38491 2953
rect 38433 2889 38436 2941
rect 38488 2889 38491 2941
rect 38433 2884 38491 2889
rect 38433 2877 38445 2884
rect 38479 2877 38491 2884
rect 38433 2825 38436 2877
rect 38488 2825 38491 2877
rect 38433 2813 38491 2825
rect 38433 2761 38436 2813
rect 38488 2761 38491 2813
rect 38433 2749 38491 2761
rect 38433 2697 38436 2749
rect 38488 2697 38491 2749
rect 38433 2685 38491 2697
rect 38433 2633 38436 2685
rect 38488 2633 38491 2685
rect 38433 2621 38491 2633
rect 38433 2569 38436 2621
rect 38488 2569 38491 2621
rect 38433 2562 38445 2569
rect 38479 2562 38491 2569
rect 38433 2557 38491 2562
rect 38433 2505 38436 2557
rect 38488 2505 38491 2557
rect 38433 2493 38445 2505
rect 38479 2493 38491 2505
rect 38433 2441 38436 2493
rect 38488 2441 38491 2493
rect 38433 2429 38445 2441
rect 38479 2429 38491 2441
rect 38433 2377 38436 2429
rect 38488 2377 38491 2429
rect 38433 2365 38445 2377
rect 38479 2365 38491 2377
rect 38433 2313 38436 2365
rect 38488 2313 38491 2365
rect 38433 2308 38491 2313
rect 38433 2301 38445 2308
rect 38479 2301 38491 2308
rect 38433 2249 38436 2301
rect 38488 2249 38491 2301
rect 38433 2237 38491 2249
rect 38433 2185 38436 2237
rect 38488 2185 38491 2237
rect 38433 2173 38491 2185
rect 38433 2121 38436 2173
rect 38488 2121 38491 2173
rect 38433 2109 38491 2121
rect 38433 2057 38436 2109
rect 38488 2057 38491 2109
rect 38433 2045 38491 2057
rect 38433 1993 38436 2045
rect 38488 1993 38491 2045
rect 38433 1986 38445 1993
rect 38479 1986 38491 1993
rect 38433 1981 38491 1986
rect 38433 1929 38436 1981
rect 38488 1929 38491 1981
rect 38433 1917 38445 1929
rect 38479 1917 38491 1929
rect 38433 1865 38436 1917
rect 38488 1865 38491 1917
rect 38433 1853 38445 1865
rect 38479 1853 38491 1865
rect 38433 1801 38436 1853
rect 38488 1801 38491 1853
rect 38433 1789 38445 1801
rect 38479 1789 38491 1801
rect 38433 1737 38436 1789
rect 38488 1737 38491 1789
rect 38433 1732 38491 1737
rect 38433 1725 38445 1732
rect 38479 1725 38491 1732
rect 38433 1673 38436 1725
rect 38488 1673 38491 1725
rect 38433 1661 38491 1673
rect 38433 1609 38436 1661
rect 38488 1609 38491 1661
rect 38433 1597 38491 1609
rect 38433 1545 38436 1597
rect 38488 1545 38491 1597
rect 38433 1533 38491 1545
rect 38433 1481 38436 1533
rect 38488 1481 38491 1533
rect 38433 1469 38491 1481
rect 38433 1417 38436 1469
rect 38488 1417 38491 1469
rect 38433 1410 38445 1417
rect 38479 1410 38491 1417
rect 38433 1405 38491 1410
rect 38433 1353 38436 1405
rect 38488 1353 38491 1405
rect 38433 1341 38445 1353
rect 38479 1341 38491 1353
rect 38433 1289 38436 1341
rect 38488 1289 38491 1341
rect 38433 1277 38445 1289
rect 38479 1277 38491 1289
rect 38433 1225 38436 1277
rect 38488 1225 38491 1277
rect 38433 1213 38445 1225
rect 38479 1213 38491 1225
rect 38433 1161 38436 1213
rect 38488 1161 38491 1213
rect 38433 1147 38491 1161
rect 38532 3133 38584 3147
rect 38532 3069 38541 3081
rect 38575 3069 38584 3081
rect 38532 3005 38541 3017
rect 38575 3005 38584 3017
rect 38532 2941 38541 2953
rect 38575 2941 38584 2953
rect 38532 2884 38584 2889
rect 38532 2877 38541 2884
rect 38575 2877 38584 2884
rect 38532 2813 38584 2825
rect 38532 2749 38584 2761
rect 38532 2685 38584 2697
rect 38532 2621 38584 2633
rect 38532 2562 38541 2569
rect 38575 2562 38584 2569
rect 38532 2557 38584 2562
rect 38532 2493 38541 2505
rect 38575 2493 38584 2505
rect 38532 2429 38541 2441
rect 38575 2429 38584 2441
rect 38532 2365 38541 2377
rect 38575 2365 38584 2377
rect 38532 2308 38584 2313
rect 38532 2301 38541 2308
rect 38575 2301 38584 2308
rect 38532 2237 38584 2249
rect 38532 2173 38584 2185
rect 38532 2109 38584 2121
rect 38532 2045 38584 2057
rect 38532 1986 38541 1993
rect 38575 1986 38584 1993
rect 38532 1981 38584 1986
rect 38532 1917 38541 1929
rect 38575 1917 38584 1929
rect 38532 1853 38541 1865
rect 38575 1853 38584 1865
rect 38532 1789 38541 1801
rect 38575 1789 38584 1801
rect 38532 1732 38584 1737
rect 38532 1725 38541 1732
rect 38575 1725 38584 1732
rect 38532 1661 38584 1673
rect 38532 1597 38584 1609
rect 38532 1533 38584 1545
rect 38532 1469 38584 1481
rect 38532 1410 38541 1417
rect 38575 1410 38584 1417
rect 38532 1405 38584 1410
rect 38532 1341 38541 1353
rect 38575 1341 38584 1353
rect 38532 1277 38541 1289
rect 38575 1277 38584 1289
rect 38532 1213 38541 1225
rect 38575 1213 38584 1225
rect 38532 1147 38584 1161
rect 38625 3132 38683 3146
rect 38625 3080 38628 3132
rect 38680 3080 38683 3132
rect 38625 3068 38637 3080
rect 38671 3068 38683 3080
rect 38625 3016 38628 3068
rect 38680 3016 38683 3068
rect 38625 3004 38637 3016
rect 38671 3004 38683 3016
rect 38625 2952 38628 3004
rect 38680 2952 38683 3004
rect 38625 2940 38637 2952
rect 38671 2940 38683 2952
rect 38625 2888 38628 2940
rect 38680 2888 38683 2940
rect 38625 2883 38683 2888
rect 38625 2876 38637 2883
rect 38671 2876 38683 2883
rect 38625 2824 38628 2876
rect 38680 2824 38683 2876
rect 38625 2812 38683 2824
rect 38625 2760 38628 2812
rect 38680 2760 38683 2812
rect 38625 2748 38683 2760
rect 38625 2696 38628 2748
rect 38680 2696 38683 2748
rect 38625 2684 38683 2696
rect 38625 2632 38628 2684
rect 38680 2632 38683 2684
rect 38625 2620 38683 2632
rect 38625 2568 38628 2620
rect 38680 2568 38683 2620
rect 38625 2561 38637 2568
rect 38671 2561 38683 2568
rect 38625 2556 38683 2561
rect 38625 2504 38628 2556
rect 38680 2504 38683 2556
rect 38625 2492 38637 2504
rect 38671 2492 38683 2504
rect 38625 2440 38628 2492
rect 38680 2440 38683 2492
rect 38625 2428 38637 2440
rect 38671 2428 38683 2440
rect 38625 2376 38628 2428
rect 38680 2376 38683 2428
rect 38625 2364 38637 2376
rect 38671 2364 38683 2376
rect 38625 2312 38628 2364
rect 38680 2312 38683 2364
rect 38625 2307 38683 2312
rect 38625 2300 38637 2307
rect 38671 2300 38683 2307
rect 38625 2248 38628 2300
rect 38680 2248 38683 2300
rect 38625 2236 38683 2248
rect 38625 2184 38628 2236
rect 38680 2184 38683 2236
rect 38625 2172 38683 2184
rect 38625 2120 38628 2172
rect 38680 2120 38683 2172
rect 38625 2108 38683 2120
rect 38625 2056 38628 2108
rect 38680 2056 38683 2108
rect 38625 2044 38683 2056
rect 38625 1992 38628 2044
rect 38680 1992 38683 2044
rect 38625 1985 38637 1992
rect 38671 1985 38683 1992
rect 38625 1980 38683 1985
rect 38625 1928 38628 1980
rect 38680 1928 38683 1980
rect 38625 1916 38637 1928
rect 38671 1916 38683 1928
rect 38625 1864 38628 1916
rect 38680 1864 38683 1916
rect 38625 1852 38637 1864
rect 38671 1852 38683 1864
rect 38625 1800 38628 1852
rect 38680 1800 38683 1852
rect 38625 1788 38637 1800
rect 38671 1788 38683 1800
rect 38625 1736 38628 1788
rect 38680 1736 38683 1788
rect 38625 1731 38683 1736
rect 38625 1724 38637 1731
rect 38671 1724 38683 1731
rect 38625 1672 38628 1724
rect 38680 1672 38683 1724
rect 38625 1660 38683 1672
rect 38625 1608 38628 1660
rect 38680 1608 38683 1660
rect 38625 1596 38683 1608
rect 38625 1544 38628 1596
rect 38680 1544 38683 1596
rect 38625 1532 38683 1544
rect 38625 1480 38628 1532
rect 38680 1480 38683 1532
rect 38625 1468 38683 1480
rect 38625 1416 38628 1468
rect 38680 1416 38683 1468
rect 38625 1409 38637 1416
rect 38671 1409 38683 1416
rect 38625 1404 38683 1409
rect 38625 1352 38628 1404
rect 38680 1352 38683 1404
rect 38625 1340 38637 1352
rect 38671 1340 38683 1352
rect 38625 1288 38628 1340
rect 38680 1288 38683 1340
rect 38625 1276 38637 1288
rect 38671 1276 38683 1288
rect 38625 1224 38628 1276
rect 38680 1224 38683 1276
rect 38625 1212 38637 1224
rect 38671 1212 38683 1224
rect 38625 1160 38628 1212
rect 38680 1160 38683 1212
rect 38625 1146 38683 1160
rect 38912 1112 38986 3180
rect 29070 1110 38986 1112
rect 29040 1099 38986 1110
rect 29040 1065 29100 1099
rect 29134 1065 29172 1099
rect 29206 1065 29244 1099
rect 29278 1065 29316 1099
rect 29350 1065 29388 1099
rect 29422 1065 29460 1099
rect 29494 1065 29532 1099
rect 29566 1065 29604 1099
rect 29638 1065 29676 1099
rect 29710 1065 29748 1099
rect 29782 1065 29820 1099
rect 29854 1065 29892 1099
rect 29926 1065 29964 1099
rect 29998 1065 30036 1099
rect 30070 1065 30108 1099
rect 30142 1065 30180 1099
rect 30214 1065 30252 1099
rect 30286 1065 30324 1099
rect 30358 1065 30396 1099
rect 30430 1065 30468 1099
rect 30502 1065 30540 1099
rect 30574 1065 30612 1099
rect 30646 1065 30684 1099
rect 30718 1065 30756 1099
rect 30790 1065 30828 1099
rect 30862 1065 30900 1099
rect 30934 1065 30972 1099
rect 31006 1065 31044 1099
rect 31078 1065 31116 1099
rect 31150 1065 31188 1099
rect 31222 1065 31260 1099
rect 31294 1065 31332 1099
rect 31366 1065 31404 1099
rect 31438 1065 31476 1099
rect 31510 1065 31548 1099
rect 31582 1065 31620 1099
rect 31654 1065 31692 1099
rect 31726 1065 31764 1099
rect 31798 1065 31836 1099
rect 31870 1065 31908 1099
rect 31942 1065 31980 1099
rect 32014 1065 32052 1099
rect 32086 1065 32124 1099
rect 32158 1065 32196 1099
rect 32230 1065 32268 1099
rect 32302 1065 32340 1099
rect 32374 1065 32412 1099
rect 32446 1065 32484 1099
rect 32518 1065 32556 1099
rect 32590 1065 32628 1099
rect 32662 1065 32700 1099
rect 32734 1065 32772 1099
rect 32806 1065 32844 1099
rect 32878 1065 32916 1099
rect 32950 1065 32988 1099
rect 33022 1065 33060 1099
rect 33094 1065 33132 1099
rect 33166 1065 33204 1099
rect 33238 1065 33276 1099
rect 33310 1065 33348 1099
rect 33382 1065 33420 1099
rect 33454 1065 33492 1099
rect 33526 1065 33564 1099
rect 33598 1065 33636 1099
rect 33670 1065 33708 1099
rect 33742 1065 33780 1099
rect 33814 1065 33852 1099
rect 33886 1065 33924 1099
rect 33958 1065 33996 1099
rect 34030 1065 34068 1099
rect 34102 1065 34140 1099
rect 34174 1065 34212 1099
rect 34246 1065 34284 1099
rect 34318 1065 34356 1099
rect 34390 1065 34428 1099
rect 34462 1065 34500 1099
rect 34534 1065 34572 1099
rect 34606 1065 34644 1099
rect 34678 1065 34716 1099
rect 34750 1065 34788 1099
rect 34822 1065 34860 1099
rect 34894 1065 34932 1099
rect 34966 1065 35004 1099
rect 35038 1065 35076 1099
rect 35110 1065 35148 1099
rect 35182 1065 35220 1099
rect 35254 1065 35292 1099
rect 35326 1065 35364 1099
rect 35398 1065 35436 1099
rect 35470 1065 35508 1099
rect 35542 1065 35580 1099
rect 35614 1065 35652 1099
rect 35686 1065 35724 1099
rect 35758 1065 35796 1099
rect 35830 1065 35868 1099
rect 35902 1065 35940 1099
rect 35974 1065 36012 1099
rect 36046 1065 36084 1099
rect 36118 1065 36156 1099
rect 36190 1065 36228 1099
rect 36262 1065 36300 1099
rect 36334 1065 36372 1099
rect 36406 1065 36444 1099
rect 36478 1065 36516 1099
rect 36550 1065 36588 1099
rect 36622 1065 36660 1099
rect 36694 1065 36732 1099
rect 36766 1065 36804 1099
rect 36838 1065 36876 1099
rect 36910 1065 36948 1099
rect 36982 1065 37020 1099
rect 37054 1065 37092 1099
rect 37126 1065 37164 1099
rect 37198 1065 37236 1099
rect 37270 1065 37308 1099
rect 37342 1065 37380 1099
rect 37414 1065 37452 1099
rect 37486 1065 37524 1099
rect 37558 1065 37596 1099
rect 37630 1065 37668 1099
rect 37702 1065 37740 1099
rect 37774 1065 37812 1099
rect 37846 1065 37884 1099
rect 37918 1065 37956 1099
rect 37990 1065 38028 1099
rect 38062 1065 38100 1099
rect 38134 1065 38172 1099
rect 38206 1065 38244 1099
rect 38278 1065 38316 1099
rect 38350 1065 38388 1099
rect 38422 1065 38460 1099
rect 38494 1065 38986 1099
rect 29040 1042 38986 1065
<< via1 >>
rect 29028 3100 29080 3133
rect 29028 3081 29037 3100
rect 29037 3081 29071 3100
rect 29071 3081 29080 3100
rect 29028 3066 29037 3069
rect 29037 3066 29071 3069
rect 29071 3066 29080 3069
rect 29028 3028 29080 3066
rect 29028 3017 29037 3028
rect 29037 3017 29071 3028
rect 29071 3017 29080 3028
rect 29028 2994 29037 3005
rect 29037 2994 29071 3005
rect 29071 2994 29080 3005
rect 29028 2956 29080 2994
rect 29028 2953 29037 2956
rect 29037 2953 29071 2956
rect 29071 2953 29080 2956
rect 29028 2922 29037 2941
rect 29037 2922 29071 2941
rect 29071 2922 29080 2941
rect 29028 2889 29080 2922
rect 29028 2850 29037 2877
rect 29037 2850 29071 2877
rect 29071 2850 29080 2877
rect 29028 2825 29080 2850
rect 29028 2812 29080 2813
rect 29028 2778 29037 2812
rect 29037 2778 29071 2812
rect 29071 2778 29080 2812
rect 29028 2761 29080 2778
rect 29028 2740 29080 2749
rect 29028 2706 29037 2740
rect 29037 2706 29071 2740
rect 29071 2706 29080 2740
rect 29028 2697 29080 2706
rect 29028 2668 29080 2685
rect 29028 2634 29037 2668
rect 29037 2634 29071 2668
rect 29071 2634 29080 2668
rect 29028 2633 29080 2634
rect 29028 2596 29080 2621
rect 29028 2569 29037 2596
rect 29037 2569 29071 2596
rect 29071 2569 29080 2596
rect 29028 2524 29080 2557
rect 29028 2505 29037 2524
rect 29037 2505 29071 2524
rect 29071 2505 29080 2524
rect 29028 2490 29037 2493
rect 29037 2490 29071 2493
rect 29071 2490 29080 2493
rect 29028 2452 29080 2490
rect 29028 2441 29037 2452
rect 29037 2441 29071 2452
rect 29071 2441 29080 2452
rect 29028 2418 29037 2429
rect 29037 2418 29071 2429
rect 29071 2418 29080 2429
rect 29028 2380 29080 2418
rect 29028 2377 29037 2380
rect 29037 2377 29071 2380
rect 29071 2377 29080 2380
rect 29028 2346 29037 2365
rect 29037 2346 29071 2365
rect 29071 2346 29080 2365
rect 29028 2313 29080 2346
rect 29028 2274 29037 2301
rect 29037 2274 29071 2301
rect 29071 2274 29080 2301
rect 29028 2249 29080 2274
rect 29028 2236 29080 2237
rect 29028 2202 29037 2236
rect 29037 2202 29071 2236
rect 29071 2202 29080 2236
rect 29028 2185 29080 2202
rect 29028 2164 29080 2173
rect 29028 2130 29037 2164
rect 29037 2130 29071 2164
rect 29071 2130 29080 2164
rect 29028 2121 29080 2130
rect 29028 2092 29080 2109
rect 29028 2058 29037 2092
rect 29037 2058 29071 2092
rect 29071 2058 29080 2092
rect 29028 2057 29080 2058
rect 29028 2020 29080 2045
rect 29028 1993 29037 2020
rect 29037 1993 29071 2020
rect 29071 1993 29080 2020
rect 29028 1948 29080 1981
rect 29028 1929 29037 1948
rect 29037 1929 29071 1948
rect 29071 1929 29080 1948
rect 29028 1914 29037 1917
rect 29037 1914 29071 1917
rect 29071 1914 29080 1917
rect 29028 1876 29080 1914
rect 29028 1865 29037 1876
rect 29037 1865 29071 1876
rect 29071 1865 29080 1876
rect 29028 1842 29037 1853
rect 29037 1842 29071 1853
rect 29071 1842 29080 1853
rect 29028 1804 29080 1842
rect 29028 1801 29037 1804
rect 29037 1801 29071 1804
rect 29071 1801 29080 1804
rect 29028 1770 29037 1789
rect 29037 1770 29071 1789
rect 29071 1770 29080 1789
rect 29028 1737 29080 1770
rect 29028 1698 29037 1725
rect 29037 1698 29071 1725
rect 29071 1698 29080 1725
rect 29028 1673 29080 1698
rect 29028 1660 29080 1661
rect 29028 1626 29037 1660
rect 29037 1626 29071 1660
rect 29071 1626 29080 1660
rect 29028 1609 29080 1626
rect 29028 1588 29080 1597
rect 29028 1554 29037 1588
rect 29037 1554 29071 1588
rect 29071 1554 29080 1588
rect 29028 1545 29080 1554
rect 29028 1516 29080 1533
rect 29028 1482 29037 1516
rect 29037 1482 29071 1516
rect 29071 1482 29080 1516
rect 29028 1481 29080 1482
rect 29028 1444 29080 1469
rect 29028 1417 29037 1444
rect 29037 1417 29071 1444
rect 29071 1417 29080 1444
rect 29028 1372 29080 1405
rect 29028 1353 29037 1372
rect 29037 1353 29071 1372
rect 29071 1353 29080 1372
rect 29028 1338 29037 1341
rect 29037 1338 29071 1341
rect 29071 1338 29080 1341
rect 29028 1300 29080 1338
rect 29028 1289 29037 1300
rect 29037 1289 29071 1300
rect 29071 1289 29080 1300
rect 29028 1266 29037 1277
rect 29037 1266 29071 1277
rect 29071 1266 29080 1277
rect 29028 1228 29080 1266
rect 29028 1225 29037 1228
rect 29037 1225 29071 1228
rect 29071 1225 29080 1228
rect 29028 1194 29037 1213
rect 29037 1194 29071 1213
rect 29071 1194 29080 1213
rect 29028 1161 29080 1194
rect 29124 3100 29176 3133
rect 29124 3081 29133 3100
rect 29133 3081 29167 3100
rect 29167 3081 29176 3100
rect 29124 3066 29133 3069
rect 29133 3066 29167 3069
rect 29167 3066 29176 3069
rect 29124 3028 29176 3066
rect 29124 3017 29133 3028
rect 29133 3017 29167 3028
rect 29167 3017 29176 3028
rect 29124 2994 29133 3005
rect 29133 2994 29167 3005
rect 29167 2994 29176 3005
rect 29124 2956 29176 2994
rect 29124 2953 29133 2956
rect 29133 2953 29167 2956
rect 29167 2953 29176 2956
rect 29124 2922 29133 2941
rect 29133 2922 29167 2941
rect 29167 2922 29176 2941
rect 29124 2889 29176 2922
rect 29124 2850 29133 2877
rect 29133 2850 29167 2877
rect 29167 2850 29176 2877
rect 29124 2825 29176 2850
rect 29124 2812 29176 2813
rect 29124 2778 29133 2812
rect 29133 2778 29167 2812
rect 29167 2778 29176 2812
rect 29124 2761 29176 2778
rect 29124 2740 29176 2749
rect 29124 2706 29133 2740
rect 29133 2706 29167 2740
rect 29167 2706 29176 2740
rect 29124 2697 29176 2706
rect 29124 2668 29176 2685
rect 29124 2634 29133 2668
rect 29133 2634 29167 2668
rect 29167 2634 29176 2668
rect 29124 2633 29176 2634
rect 29124 2596 29176 2621
rect 29124 2569 29133 2596
rect 29133 2569 29167 2596
rect 29167 2569 29176 2596
rect 29124 2524 29176 2557
rect 29124 2505 29133 2524
rect 29133 2505 29167 2524
rect 29167 2505 29176 2524
rect 29124 2490 29133 2493
rect 29133 2490 29167 2493
rect 29167 2490 29176 2493
rect 29124 2452 29176 2490
rect 29124 2441 29133 2452
rect 29133 2441 29167 2452
rect 29167 2441 29176 2452
rect 29124 2418 29133 2429
rect 29133 2418 29167 2429
rect 29167 2418 29176 2429
rect 29124 2380 29176 2418
rect 29124 2377 29133 2380
rect 29133 2377 29167 2380
rect 29167 2377 29176 2380
rect 29124 2346 29133 2365
rect 29133 2346 29167 2365
rect 29167 2346 29176 2365
rect 29124 2313 29176 2346
rect 29124 2274 29133 2301
rect 29133 2274 29167 2301
rect 29167 2274 29176 2301
rect 29124 2249 29176 2274
rect 29124 2236 29176 2237
rect 29124 2202 29133 2236
rect 29133 2202 29167 2236
rect 29167 2202 29176 2236
rect 29124 2185 29176 2202
rect 29124 2164 29176 2173
rect 29124 2130 29133 2164
rect 29133 2130 29167 2164
rect 29167 2130 29176 2164
rect 29124 2121 29176 2130
rect 29124 2092 29176 2109
rect 29124 2058 29133 2092
rect 29133 2058 29167 2092
rect 29167 2058 29176 2092
rect 29124 2057 29176 2058
rect 29124 2020 29176 2045
rect 29124 1993 29133 2020
rect 29133 1993 29167 2020
rect 29167 1993 29176 2020
rect 29124 1948 29176 1981
rect 29124 1929 29133 1948
rect 29133 1929 29167 1948
rect 29167 1929 29176 1948
rect 29124 1914 29133 1917
rect 29133 1914 29167 1917
rect 29167 1914 29176 1917
rect 29124 1876 29176 1914
rect 29124 1865 29133 1876
rect 29133 1865 29167 1876
rect 29167 1865 29176 1876
rect 29124 1842 29133 1853
rect 29133 1842 29167 1853
rect 29167 1842 29176 1853
rect 29124 1804 29176 1842
rect 29124 1801 29133 1804
rect 29133 1801 29167 1804
rect 29167 1801 29176 1804
rect 29124 1770 29133 1789
rect 29133 1770 29167 1789
rect 29167 1770 29176 1789
rect 29124 1737 29176 1770
rect 29124 1698 29133 1725
rect 29133 1698 29167 1725
rect 29167 1698 29176 1725
rect 29124 1673 29176 1698
rect 29124 1660 29176 1661
rect 29124 1626 29133 1660
rect 29133 1626 29167 1660
rect 29167 1626 29176 1660
rect 29124 1609 29176 1626
rect 29124 1588 29176 1597
rect 29124 1554 29133 1588
rect 29133 1554 29167 1588
rect 29167 1554 29176 1588
rect 29124 1545 29176 1554
rect 29124 1516 29176 1533
rect 29124 1482 29133 1516
rect 29133 1482 29167 1516
rect 29167 1482 29176 1516
rect 29124 1481 29176 1482
rect 29124 1444 29176 1469
rect 29124 1417 29133 1444
rect 29133 1417 29167 1444
rect 29167 1417 29176 1444
rect 29124 1372 29176 1405
rect 29124 1353 29133 1372
rect 29133 1353 29167 1372
rect 29167 1353 29176 1372
rect 29124 1338 29133 1341
rect 29133 1338 29167 1341
rect 29167 1338 29176 1341
rect 29124 1300 29176 1338
rect 29124 1289 29133 1300
rect 29133 1289 29167 1300
rect 29167 1289 29176 1300
rect 29124 1266 29133 1277
rect 29133 1266 29167 1277
rect 29167 1266 29176 1277
rect 29124 1228 29176 1266
rect 29124 1225 29133 1228
rect 29133 1225 29167 1228
rect 29167 1225 29176 1228
rect 29124 1194 29133 1213
rect 29133 1194 29167 1213
rect 29167 1194 29176 1213
rect 29124 1161 29176 1194
rect 29220 3100 29272 3133
rect 29220 3081 29229 3100
rect 29229 3081 29263 3100
rect 29263 3081 29272 3100
rect 29220 3066 29229 3069
rect 29229 3066 29263 3069
rect 29263 3066 29272 3069
rect 29220 3028 29272 3066
rect 29220 3017 29229 3028
rect 29229 3017 29263 3028
rect 29263 3017 29272 3028
rect 29220 2994 29229 3005
rect 29229 2994 29263 3005
rect 29263 2994 29272 3005
rect 29220 2956 29272 2994
rect 29220 2953 29229 2956
rect 29229 2953 29263 2956
rect 29263 2953 29272 2956
rect 29220 2922 29229 2941
rect 29229 2922 29263 2941
rect 29263 2922 29272 2941
rect 29220 2889 29272 2922
rect 29220 2850 29229 2877
rect 29229 2850 29263 2877
rect 29263 2850 29272 2877
rect 29220 2825 29272 2850
rect 29220 2812 29272 2813
rect 29220 2778 29229 2812
rect 29229 2778 29263 2812
rect 29263 2778 29272 2812
rect 29220 2761 29272 2778
rect 29220 2740 29272 2749
rect 29220 2706 29229 2740
rect 29229 2706 29263 2740
rect 29263 2706 29272 2740
rect 29220 2697 29272 2706
rect 29220 2668 29272 2685
rect 29220 2634 29229 2668
rect 29229 2634 29263 2668
rect 29263 2634 29272 2668
rect 29220 2633 29272 2634
rect 29220 2596 29272 2621
rect 29220 2569 29229 2596
rect 29229 2569 29263 2596
rect 29263 2569 29272 2596
rect 29220 2524 29272 2557
rect 29220 2505 29229 2524
rect 29229 2505 29263 2524
rect 29263 2505 29272 2524
rect 29220 2490 29229 2493
rect 29229 2490 29263 2493
rect 29263 2490 29272 2493
rect 29220 2452 29272 2490
rect 29220 2441 29229 2452
rect 29229 2441 29263 2452
rect 29263 2441 29272 2452
rect 29220 2418 29229 2429
rect 29229 2418 29263 2429
rect 29263 2418 29272 2429
rect 29220 2380 29272 2418
rect 29220 2377 29229 2380
rect 29229 2377 29263 2380
rect 29263 2377 29272 2380
rect 29220 2346 29229 2365
rect 29229 2346 29263 2365
rect 29263 2346 29272 2365
rect 29220 2313 29272 2346
rect 29220 2274 29229 2301
rect 29229 2274 29263 2301
rect 29263 2274 29272 2301
rect 29220 2249 29272 2274
rect 29220 2236 29272 2237
rect 29220 2202 29229 2236
rect 29229 2202 29263 2236
rect 29263 2202 29272 2236
rect 29220 2185 29272 2202
rect 29220 2164 29272 2173
rect 29220 2130 29229 2164
rect 29229 2130 29263 2164
rect 29263 2130 29272 2164
rect 29220 2121 29272 2130
rect 29220 2092 29272 2109
rect 29220 2058 29229 2092
rect 29229 2058 29263 2092
rect 29263 2058 29272 2092
rect 29220 2057 29272 2058
rect 29220 2020 29272 2045
rect 29220 1993 29229 2020
rect 29229 1993 29263 2020
rect 29263 1993 29272 2020
rect 29220 1948 29272 1981
rect 29220 1929 29229 1948
rect 29229 1929 29263 1948
rect 29263 1929 29272 1948
rect 29220 1914 29229 1917
rect 29229 1914 29263 1917
rect 29263 1914 29272 1917
rect 29220 1876 29272 1914
rect 29220 1865 29229 1876
rect 29229 1865 29263 1876
rect 29263 1865 29272 1876
rect 29220 1842 29229 1853
rect 29229 1842 29263 1853
rect 29263 1842 29272 1853
rect 29220 1804 29272 1842
rect 29220 1801 29229 1804
rect 29229 1801 29263 1804
rect 29263 1801 29272 1804
rect 29220 1770 29229 1789
rect 29229 1770 29263 1789
rect 29263 1770 29272 1789
rect 29220 1737 29272 1770
rect 29220 1698 29229 1725
rect 29229 1698 29263 1725
rect 29263 1698 29272 1725
rect 29220 1673 29272 1698
rect 29220 1660 29272 1661
rect 29220 1626 29229 1660
rect 29229 1626 29263 1660
rect 29263 1626 29272 1660
rect 29220 1609 29272 1626
rect 29220 1588 29272 1597
rect 29220 1554 29229 1588
rect 29229 1554 29263 1588
rect 29263 1554 29272 1588
rect 29220 1545 29272 1554
rect 29220 1516 29272 1533
rect 29220 1482 29229 1516
rect 29229 1482 29263 1516
rect 29263 1482 29272 1516
rect 29220 1481 29272 1482
rect 29220 1444 29272 1469
rect 29220 1417 29229 1444
rect 29229 1417 29263 1444
rect 29263 1417 29272 1444
rect 29220 1372 29272 1405
rect 29220 1353 29229 1372
rect 29229 1353 29263 1372
rect 29263 1353 29272 1372
rect 29220 1338 29229 1341
rect 29229 1338 29263 1341
rect 29263 1338 29272 1341
rect 29220 1300 29272 1338
rect 29220 1289 29229 1300
rect 29229 1289 29263 1300
rect 29263 1289 29272 1300
rect 29220 1266 29229 1277
rect 29229 1266 29263 1277
rect 29263 1266 29272 1277
rect 29220 1228 29272 1266
rect 29220 1225 29229 1228
rect 29229 1225 29263 1228
rect 29263 1225 29272 1228
rect 29220 1194 29229 1213
rect 29229 1194 29263 1213
rect 29263 1194 29272 1213
rect 29220 1161 29272 1194
rect 29316 3100 29368 3133
rect 29316 3081 29325 3100
rect 29325 3081 29359 3100
rect 29359 3081 29368 3100
rect 29316 3066 29325 3069
rect 29325 3066 29359 3069
rect 29359 3066 29368 3069
rect 29316 3028 29368 3066
rect 29316 3017 29325 3028
rect 29325 3017 29359 3028
rect 29359 3017 29368 3028
rect 29316 2994 29325 3005
rect 29325 2994 29359 3005
rect 29359 2994 29368 3005
rect 29316 2956 29368 2994
rect 29316 2953 29325 2956
rect 29325 2953 29359 2956
rect 29359 2953 29368 2956
rect 29316 2922 29325 2941
rect 29325 2922 29359 2941
rect 29359 2922 29368 2941
rect 29316 2889 29368 2922
rect 29316 2850 29325 2877
rect 29325 2850 29359 2877
rect 29359 2850 29368 2877
rect 29316 2825 29368 2850
rect 29316 2812 29368 2813
rect 29316 2778 29325 2812
rect 29325 2778 29359 2812
rect 29359 2778 29368 2812
rect 29316 2761 29368 2778
rect 29316 2740 29368 2749
rect 29316 2706 29325 2740
rect 29325 2706 29359 2740
rect 29359 2706 29368 2740
rect 29316 2697 29368 2706
rect 29316 2668 29368 2685
rect 29316 2634 29325 2668
rect 29325 2634 29359 2668
rect 29359 2634 29368 2668
rect 29316 2633 29368 2634
rect 29316 2596 29368 2621
rect 29316 2569 29325 2596
rect 29325 2569 29359 2596
rect 29359 2569 29368 2596
rect 29316 2524 29368 2557
rect 29316 2505 29325 2524
rect 29325 2505 29359 2524
rect 29359 2505 29368 2524
rect 29316 2490 29325 2493
rect 29325 2490 29359 2493
rect 29359 2490 29368 2493
rect 29316 2452 29368 2490
rect 29316 2441 29325 2452
rect 29325 2441 29359 2452
rect 29359 2441 29368 2452
rect 29316 2418 29325 2429
rect 29325 2418 29359 2429
rect 29359 2418 29368 2429
rect 29316 2380 29368 2418
rect 29316 2377 29325 2380
rect 29325 2377 29359 2380
rect 29359 2377 29368 2380
rect 29316 2346 29325 2365
rect 29325 2346 29359 2365
rect 29359 2346 29368 2365
rect 29316 2313 29368 2346
rect 29316 2274 29325 2301
rect 29325 2274 29359 2301
rect 29359 2274 29368 2301
rect 29316 2249 29368 2274
rect 29316 2236 29368 2237
rect 29316 2202 29325 2236
rect 29325 2202 29359 2236
rect 29359 2202 29368 2236
rect 29316 2185 29368 2202
rect 29316 2164 29368 2173
rect 29316 2130 29325 2164
rect 29325 2130 29359 2164
rect 29359 2130 29368 2164
rect 29316 2121 29368 2130
rect 29316 2092 29368 2109
rect 29316 2058 29325 2092
rect 29325 2058 29359 2092
rect 29359 2058 29368 2092
rect 29316 2057 29368 2058
rect 29316 2020 29368 2045
rect 29316 1993 29325 2020
rect 29325 1993 29359 2020
rect 29359 1993 29368 2020
rect 29316 1948 29368 1981
rect 29316 1929 29325 1948
rect 29325 1929 29359 1948
rect 29359 1929 29368 1948
rect 29316 1914 29325 1917
rect 29325 1914 29359 1917
rect 29359 1914 29368 1917
rect 29316 1876 29368 1914
rect 29316 1865 29325 1876
rect 29325 1865 29359 1876
rect 29359 1865 29368 1876
rect 29316 1842 29325 1853
rect 29325 1842 29359 1853
rect 29359 1842 29368 1853
rect 29316 1804 29368 1842
rect 29316 1801 29325 1804
rect 29325 1801 29359 1804
rect 29359 1801 29368 1804
rect 29316 1770 29325 1789
rect 29325 1770 29359 1789
rect 29359 1770 29368 1789
rect 29316 1737 29368 1770
rect 29316 1698 29325 1725
rect 29325 1698 29359 1725
rect 29359 1698 29368 1725
rect 29316 1673 29368 1698
rect 29316 1660 29368 1661
rect 29316 1626 29325 1660
rect 29325 1626 29359 1660
rect 29359 1626 29368 1660
rect 29316 1609 29368 1626
rect 29316 1588 29368 1597
rect 29316 1554 29325 1588
rect 29325 1554 29359 1588
rect 29359 1554 29368 1588
rect 29316 1545 29368 1554
rect 29316 1516 29368 1533
rect 29316 1482 29325 1516
rect 29325 1482 29359 1516
rect 29359 1482 29368 1516
rect 29316 1481 29368 1482
rect 29316 1444 29368 1469
rect 29316 1417 29325 1444
rect 29325 1417 29359 1444
rect 29359 1417 29368 1444
rect 29316 1372 29368 1405
rect 29316 1353 29325 1372
rect 29325 1353 29359 1372
rect 29359 1353 29368 1372
rect 29316 1338 29325 1341
rect 29325 1338 29359 1341
rect 29359 1338 29368 1341
rect 29316 1300 29368 1338
rect 29316 1289 29325 1300
rect 29325 1289 29359 1300
rect 29359 1289 29368 1300
rect 29316 1266 29325 1277
rect 29325 1266 29359 1277
rect 29359 1266 29368 1277
rect 29316 1228 29368 1266
rect 29316 1225 29325 1228
rect 29325 1225 29359 1228
rect 29359 1225 29368 1228
rect 29316 1194 29325 1213
rect 29325 1194 29359 1213
rect 29359 1194 29368 1213
rect 29316 1161 29368 1194
rect 29412 3100 29464 3133
rect 29412 3081 29421 3100
rect 29421 3081 29455 3100
rect 29455 3081 29464 3100
rect 29412 3066 29421 3069
rect 29421 3066 29455 3069
rect 29455 3066 29464 3069
rect 29412 3028 29464 3066
rect 29412 3017 29421 3028
rect 29421 3017 29455 3028
rect 29455 3017 29464 3028
rect 29412 2994 29421 3005
rect 29421 2994 29455 3005
rect 29455 2994 29464 3005
rect 29412 2956 29464 2994
rect 29412 2953 29421 2956
rect 29421 2953 29455 2956
rect 29455 2953 29464 2956
rect 29412 2922 29421 2941
rect 29421 2922 29455 2941
rect 29455 2922 29464 2941
rect 29412 2889 29464 2922
rect 29412 2850 29421 2877
rect 29421 2850 29455 2877
rect 29455 2850 29464 2877
rect 29412 2825 29464 2850
rect 29412 2812 29464 2813
rect 29412 2778 29421 2812
rect 29421 2778 29455 2812
rect 29455 2778 29464 2812
rect 29412 2761 29464 2778
rect 29412 2740 29464 2749
rect 29412 2706 29421 2740
rect 29421 2706 29455 2740
rect 29455 2706 29464 2740
rect 29412 2697 29464 2706
rect 29412 2668 29464 2685
rect 29412 2634 29421 2668
rect 29421 2634 29455 2668
rect 29455 2634 29464 2668
rect 29412 2633 29464 2634
rect 29412 2596 29464 2621
rect 29412 2569 29421 2596
rect 29421 2569 29455 2596
rect 29455 2569 29464 2596
rect 29412 2524 29464 2557
rect 29412 2505 29421 2524
rect 29421 2505 29455 2524
rect 29455 2505 29464 2524
rect 29412 2490 29421 2493
rect 29421 2490 29455 2493
rect 29455 2490 29464 2493
rect 29412 2452 29464 2490
rect 29412 2441 29421 2452
rect 29421 2441 29455 2452
rect 29455 2441 29464 2452
rect 29412 2418 29421 2429
rect 29421 2418 29455 2429
rect 29455 2418 29464 2429
rect 29412 2380 29464 2418
rect 29412 2377 29421 2380
rect 29421 2377 29455 2380
rect 29455 2377 29464 2380
rect 29412 2346 29421 2365
rect 29421 2346 29455 2365
rect 29455 2346 29464 2365
rect 29412 2313 29464 2346
rect 29412 2274 29421 2301
rect 29421 2274 29455 2301
rect 29455 2274 29464 2301
rect 29412 2249 29464 2274
rect 29412 2236 29464 2237
rect 29412 2202 29421 2236
rect 29421 2202 29455 2236
rect 29455 2202 29464 2236
rect 29412 2185 29464 2202
rect 29412 2164 29464 2173
rect 29412 2130 29421 2164
rect 29421 2130 29455 2164
rect 29455 2130 29464 2164
rect 29412 2121 29464 2130
rect 29412 2092 29464 2109
rect 29412 2058 29421 2092
rect 29421 2058 29455 2092
rect 29455 2058 29464 2092
rect 29412 2057 29464 2058
rect 29412 2020 29464 2045
rect 29412 1993 29421 2020
rect 29421 1993 29455 2020
rect 29455 1993 29464 2020
rect 29412 1948 29464 1981
rect 29412 1929 29421 1948
rect 29421 1929 29455 1948
rect 29455 1929 29464 1948
rect 29412 1914 29421 1917
rect 29421 1914 29455 1917
rect 29455 1914 29464 1917
rect 29412 1876 29464 1914
rect 29412 1865 29421 1876
rect 29421 1865 29455 1876
rect 29455 1865 29464 1876
rect 29412 1842 29421 1853
rect 29421 1842 29455 1853
rect 29455 1842 29464 1853
rect 29412 1804 29464 1842
rect 29412 1801 29421 1804
rect 29421 1801 29455 1804
rect 29455 1801 29464 1804
rect 29412 1770 29421 1789
rect 29421 1770 29455 1789
rect 29455 1770 29464 1789
rect 29412 1737 29464 1770
rect 29412 1698 29421 1725
rect 29421 1698 29455 1725
rect 29455 1698 29464 1725
rect 29412 1673 29464 1698
rect 29412 1660 29464 1661
rect 29412 1626 29421 1660
rect 29421 1626 29455 1660
rect 29455 1626 29464 1660
rect 29412 1609 29464 1626
rect 29412 1588 29464 1597
rect 29412 1554 29421 1588
rect 29421 1554 29455 1588
rect 29455 1554 29464 1588
rect 29412 1545 29464 1554
rect 29412 1516 29464 1533
rect 29412 1482 29421 1516
rect 29421 1482 29455 1516
rect 29455 1482 29464 1516
rect 29412 1481 29464 1482
rect 29412 1444 29464 1469
rect 29412 1417 29421 1444
rect 29421 1417 29455 1444
rect 29455 1417 29464 1444
rect 29412 1372 29464 1405
rect 29412 1353 29421 1372
rect 29421 1353 29455 1372
rect 29455 1353 29464 1372
rect 29412 1338 29421 1341
rect 29421 1338 29455 1341
rect 29455 1338 29464 1341
rect 29412 1300 29464 1338
rect 29412 1289 29421 1300
rect 29421 1289 29455 1300
rect 29455 1289 29464 1300
rect 29412 1266 29421 1277
rect 29421 1266 29455 1277
rect 29455 1266 29464 1277
rect 29412 1228 29464 1266
rect 29412 1225 29421 1228
rect 29421 1225 29455 1228
rect 29455 1225 29464 1228
rect 29412 1194 29421 1213
rect 29421 1194 29455 1213
rect 29455 1194 29464 1213
rect 29412 1161 29464 1194
rect 29508 3100 29560 3133
rect 29508 3081 29517 3100
rect 29517 3081 29551 3100
rect 29551 3081 29560 3100
rect 29508 3066 29517 3069
rect 29517 3066 29551 3069
rect 29551 3066 29560 3069
rect 29508 3028 29560 3066
rect 29508 3017 29517 3028
rect 29517 3017 29551 3028
rect 29551 3017 29560 3028
rect 29508 2994 29517 3005
rect 29517 2994 29551 3005
rect 29551 2994 29560 3005
rect 29508 2956 29560 2994
rect 29508 2953 29517 2956
rect 29517 2953 29551 2956
rect 29551 2953 29560 2956
rect 29508 2922 29517 2941
rect 29517 2922 29551 2941
rect 29551 2922 29560 2941
rect 29508 2889 29560 2922
rect 29508 2850 29517 2877
rect 29517 2850 29551 2877
rect 29551 2850 29560 2877
rect 29508 2825 29560 2850
rect 29508 2812 29560 2813
rect 29508 2778 29517 2812
rect 29517 2778 29551 2812
rect 29551 2778 29560 2812
rect 29508 2761 29560 2778
rect 29508 2740 29560 2749
rect 29508 2706 29517 2740
rect 29517 2706 29551 2740
rect 29551 2706 29560 2740
rect 29508 2697 29560 2706
rect 29508 2668 29560 2685
rect 29508 2634 29517 2668
rect 29517 2634 29551 2668
rect 29551 2634 29560 2668
rect 29508 2633 29560 2634
rect 29508 2596 29560 2621
rect 29508 2569 29517 2596
rect 29517 2569 29551 2596
rect 29551 2569 29560 2596
rect 29508 2524 29560 2557
rect 29508 2505 29517 2524
rect 29517 2505 29551 2524
rect 29551 2505 29560 2524
rect 29508 2490 29517 2493
rect 29517 2490 29551 2493
rect 29551 2490 29560 2493
rect 29508 2452 29560 2490
rect 29508 2441 29517 2452
rect 29517 2441 29551 2452
rect 29551 2441 29560 2452
rect 29508 2418 29517 2429
rect 29517 2418 29551 2429
rect 29551 2418 29560 2429
rect 29508 2380 29560 2418
rect 29508 2377 29517 2380
rect 29517 2377 29551 2380
rect 29551 2377 29560 2380
rect 29508 2346 29517 2365
rect 29517 2346 29551 2365
rect 29551 2346 29560 2365
rect 29508 2313 29560 2346
rect 29508 2274 29517 2301
rect 29517 2274 29551 2301
rect 29551 2274 29560 2301
rect 29508 2249 29560 2274
rect 29508 2236 29560 2237
rect 29508 2202 29517 2236
rect 29517 2202 29551 2236
rect 29551 2202 29560 2236
rect 29508 2185 29560 2202
rect 29508 2164 29560 2173
rect 29508 2130 29517 2164
rect 29517 2130 29551 2164
rect 29551 2130 29560 2164
rect 29508 2121 29560 2130
rect 29508 2092 29560 2109
rect 29508 2058 29517 2092
rect 29517 2058 29551 2092
rect 29551 2058 29560 2092
rect 29508 2057 29560 2058
rect 29508 2020 29560 2045
rect 29508 1993 29517 2020
rect 29517 1993 29551 2020
rect 29551 1993 29560 2020
rect 29508 1948 29560 1981
rect 29508 1929 29517 1948
rect 29517 1929 29551 1948
rect 29551 1929 29560 1948
rect 29508 1914 29517 1917
rect 29517 1914 29551 1917
rect 29551 1914 29560 1917
rect 29508 1876 29560 1914
rect 29508 1865 29517 1876
rect 29517 1865 29551 1876
rect 29551 1865 29560 1876
rect 29508 1842 29517 1853
rect 29517 1842 29551 1853
rect 29551 1842 29560 1853
rect 29508 1804 29560 1842
rect 29508 1801 29517 1804
rect 29517 1801 29551 1804
rect 29551 1801 29560 1804
rect 29508 1770 29517 1789
rect 29517 1770 29551 1789
rect 29551 1770 29560 1789
rect 29508 1737 29560 1770
rect 29508 1698 29517 1725
rect 29517 1698 29551 1725
rect 29551 1698 29560 1725
rect 29508 1673 29560 1698
rect 29508 1660 29560 1661
rect 29508 1626 29517 1660
rect 29517 1626 29551 1660
rect 29551 1626 29560 1660
rect 29508 1609 29560 1626
rect 29508 1588 29560 1597
rect 29508 1554 29517 1588
rect 29517 1554 29551 1588
rect 29551 1554 29560 1588
rect 29508 1545 29560 1554
rect 29508 1516 29560 1533
rect 29508 1482 29517 1516
rect 29517 1482 29551 1516
rect 29551 1482 29560 1516
rect 29508 1481 29560 1482
rect 29508 1444 29560 1469
rect 29508 1417 29517 1444
rect 29517 1417 29551 1444
rect 29551 1417 29560 1444
rect 29508 1372 29560 1405
rect 29508 1353 29517 1372
rect 29517 1353 29551 1372
rect 29551 1353 29560 1372
rect 29508 1338 29517 1341
rect 29517 1338 29551 1341
rect 29551 1338 29560 1341
rect 29508 1300 29560 1338
rect 29508 1289 29517 1300
rect 29517 1289 29551 1300
rect 29551 1289 29560 1300
rect 29508 1266 29517 1277
rect 29517 1266 29551 1277
rect 29551 1266 29560 1277
rect 29508 1228 29560 1266
rect 29508 1225 29517 1228
rect 29517 1225 29551 1228
rect 29551 1225 29560 1228
rect 29508 1194 29517 1213
rect 29517 1194 29551 1213
rect 29551 1194 29560 1213
rect 29508 1161 29560 1194
rect 29604 3100 29656 3133
rect 29604 3081 29613 3100
rect 29613 3081 29647 3100
rect 29647 3081 29656 3100
rect 29604 3066 29613 3069
rect 29613 3066 29647 3069
rect 29647 3066 29656 3069
rect 29604 3028 29656 3066
rect 29604 3017 29613 3028
rect 29613 3017 29647 3028
rect 29647 3017 29656 3028
rect 29604 2994 29613 3005
rect 29613 2994 29647 3005
rect 29647 2994 29656 3005
rect 29604 2956 29656 2994
rect 29604 2953 29613 2956
rect 29613 2953 29647 2956
rect 29647 2953 29656 2956
rect 29604 2922 29613 2941
rect 29613 2922 29647 2941
rect 29647 2922 29656 2941
rect 29604 2889 29656 2922
rect 29604 2850 29613 2877
rect 29613 2850 29647 2877
rect 29647 2850 29656 2877
rect 29604 2825 29656 2850
rect 29604 2812 29656 2813
rect 29604 2778 29613 2812
rect 29613 2778 29647 2812
rect 29647 2778 29656 2812
rect 29604 2761 29656 2778
rect 29604 2740 29656 2749
rect 29604 2706 29613 2740
rect 29613 2706 29647 2740
rect 29647 2706 29656 2740
rect 29604 2697 29656 2706
rect 29604 2668 29656 2685
rect 29604 2634 29613 2668
rect 29613 2634 29647 2668
rect 29647 2634 29656 2668
rect 29604 2633 29656 2634
rect 29604 2596 29656 2621
rect 29604 2569 29613 2596
rect 29613 2569 29647 2596
rect 29647 2569 29656 2596
rect 29604 2524 29656 2557
rect 29604 2505 29613 2524
rect 29613 2505 29647 2524
rect 29647 2505 29656 2524
rect 29604 2490 29613 2493
rect 29613 2490 29647 2493
rect 29647 2490 29656 2493
rect 29604 2452 29656 2490
rect 29604 2441 29613 2452
rect 29613 2441 29647 2452
rect 29647 2441 29656 2452
rect 29604 2418 29613 2429
rect 29613 2418 29647 2429
rect 29647 2418 29656 2429
rect 29604 2380 29656 2418
rect 29604 2377 29613 2380
rect 29613 2377 29647 2380
rect 29647 2377 29656 2380
rect 29604 2346 29613 2365
rect 29613 2346 29647 2365
rect 29647 2346 29656 2365
rect 29604 2313 29656 2346
rect 29604 2274 29613 2301
rect 29613 2274 29647 2301
rect 29647 2274 29656 2301
rect 29604 2249 29656 2274
rect 29604 2236 29656 2237
rect 29604 2202 29613 2236
rect 29613 2202 29647 2236
rect 29647 2202 29656 2236
rect 29604 2185 29656 2202
rect 29604 2164 29656 2173
rect 29604 2130 29613 2164
rect 29613 2130 29647 2164
rect 29647 2130 29656 2164
rect 29604 2121 29656 2130
rect 29604 2092 29656 2109
rect 29604 2058 29613 2092
rect 29613 2058 29647 2092
rect 29647 2058 29656 2092
rect 29604 2057 29656 2058
rect 29604 2020 29656 2045
rect 29604 1993 29613 2020
rect 29613 1993 29647 2020
rect 29647 1993 29656 2020
rect 29604 1948 29656 1981
rect 29604 1929 29613 1948
rect 29613 1929 29647 1948
rect 29647 1929 29656 1948
rect 29604 1914 29613 1917
rect 29613 1914 29647 1917
rect 29647 1914 29656 1917
rect 29604 1876 29656 1914
rect 29604 1865 29613 1876
rect 29613 1865 29647 1876
rect 29647 1865 29656 1876
rect 29604 1842 29613 1853
rect 29613 1842 29647 1853
rect 29647 1842 29656 1853
rect 29604 1804 29656 1842
rect 29604 1801 29613 1804
rect 29613 1801 29647 1804
rect 29647 1801 29656 1804
rect 29604 1770 29613 1789
rect 29613 1770 29647 1789
rect 29647 1770 29656 1789
rect 29604 1737 29656 1770
rect 29604 1698 29613 1725
rect 29613 1698 29647 1725
rect 29647 1698 29656 1725
rect 29604 1673 29656 1698
rect 29604 1660 29656 1661
rect 29604 1626 29613 1660
rect 29613 1626 29647 1660
rect 29647 1626 29656 1660
rect 29604 1609 29656 1626
rect 29604 1588 29656 1597
rect 29604 1554 29613 1588
rect 29613 1554 29647 1588
rect 29647 1554 29656 1588
rect 29604 1545 29656 1554
rect 29604 1516 29656 1533
rect 29604 1482 29613 1516
rect 29613 1482 29647 1516
rect 29647 1482 29656 1516
rect 29604 1481 29656 1482
rect 29604 1444 29656 1469
rect 29604 1417 29613 1444
rect 29613 1417 29647 1444
rect 29647 1417 29656 1444
rect 29604 1372 29656 1405
rect 29604 1353 29613 1372
rect 29613 1353 29647 1372
rect 29647 1353 29656 1372
rect 29604 1338 29613 1341
rect 29613 1338 29647 1341
rect 29647 1338 29656 1341
rect 29604 1300 29656 1338
rect 29604 1289 29613 1300
rect 29613 1289 29647 1300
rect 29647 1289 29656 1300
rect 29604 1266 29613 1277
rect 29613 1266 29647 1277
rect 29647 1266 29656 1277
rect 29604 1228 29656 1266
rect 29604 1225 29613 1228
rect 29613 1225 29647 1228
rect 29647 1225 29656 1228
rect 29604 1194 29613 1213
rect 29613 1194 29647 1213
rect 29647 1194 29656 1213
rect 29604 1161 29656 1194
rect 29700 3100 29752 3133
rect 29700 3081 29709 3100
rect 29709 3081 29743 3100
rect 29743 3081 29752 3100
rect 29700 3066 29709 3069
rect 29709 3066 29743 3069
rect 29743 3066 29752 3069
rect 29700 3028 29752 3066
rect 29700 3017 29709 3028
rect 29709 3017 29743 3028
rect 29743 3017 29752 3028
rect 29700 2994 29709 3005
rect 29709 2994 29743 3005
rect 29743 2994 29752 3005
rect 29700 2956 29752 2994
rect 29700 2953 29709 2956
rect 29709 2953 29743 2956
rect 29743 2953 29752 2956
rect 29700 2922 29709 2941
rect 29709 2922 29743 2941
rect 29743 2922 29752 2941
rect 29700 2889 29752 2922
rect 29700 2850 29709 2877
rect 29709 2850 29743 2877
rect 29743 2850 29752 2877
rect 29700 2825 29752 2850
rect 29700 2812 29752 2813
rect 29700 2778 29709 2812
rect 29709 2778 29743 2812
rect 29743 2778 29752 2812
rect 29700 2761 29752 2778
rect 29700 2740 29752 2749
rect 29700 2706 29709 2740
rect 29709 2706 29743 2740
rect 29743 2706 29752 2740
rect 29700 2697 29752 2706
rect 29700 2668 29752 2685
rect 29700 2634 29709 2668
rect 29709 2634 29743 2668
rect 29743 2634 29752 2668
rect 29700 2633 29752 2634
rect 29700 2596 29752 2621
rect 29700 2569 29709 2596
rect 29709 2569 29743 2596
rect 29743 2569 29752 2596
rect 29700 2524 29752 2557
rect 29700 2505 29709 2524
rect 29709 2505 29743 2524
rect 29743 2505 29752 2524
rect 29700 2490 29709 2493
rect 29709 2490 29743 2493
rect 29743 2490 29752 2493
rect 29700 2452 29752 2490
rect 29700 2441 29709 2452
rect 29709 2441 29743 2452
rect 29743 2441 29752 2452
rect 29700 2418 29709 2429
rect 29709 2418 29743 2429
rect 29743 2418 29752 2429
rect 29700 2380 29752 2418
rect 29700 2377 29709 2380
rect 29709 2377 29743 2380
rect 29743 2377 29752 2380
rect 29700 2346 29709 2365
rect 29709 2346 29743 2365
rect 29743 2346 29752 2365
rect 29700 2313 29752 2346
rect 29700 2274 29709 2301
rect 29709 2274 29743 2301
rect 29743 2274 29752 2301
rect 29700 2249 29752 2274
rect 29700 2236 29752 2237
rect 29700 2202 29709 2236
rect 29709 2202 29743 2236
rect 29743 2202 29752 2236
rect 29700 2185 29752 2202
rect 29700 2164 29752 2173
rect 29700 2130 29709 2164
rect 29709 2130 29743 2164
rect 29743 2130 29752 2164
rect 29700 2121 29752 2130
rect 29700 2092 29752 2109
rect 29700 2058 29709 2092
rect 29709 2058 29743 2092
rect 29743 2058 29752 2092
rect 29700 2057 29752 2058
rect 29700 2020 29752 2045
rect 29700 1993 29709 2020
rect 29709 1993 29743 2020
rect 29743 1993 29752 2020
rect 29700 1948 29752 1981
rect 29700 1929 29709 1948
rect 29709 1929 29743 1948
rect 29743 1929 29752 1948
rect 29700 1914 29709 1917
rect 29709 1914 29743 1917
rect 29743 1914 29752 1917
rect 29700 1876 29752 1914
rect 29700 1865 29709 1876
rect 29709 1865 29743 1876
rect 29743 1865 29752 1876
rect 29700 1842 29709 1853
rect 29709 1842 29743 1853
rect 29743 1842 29752 1853
rect 29700 1804 29752 1842
rect 29700 1801 29709 1804
rect 29709 1801 29743 1804
rect 29743 1801 29752 1804
rect 29700 1770 29709 1789
rect 29709 1770 29743 1789
rect 29743 1770 29752 1789
rect 29700 1737 29752 1770
rect 29700 1698 29709 1725
rect 29709 1698 29743 1725
rect 29743 1698 29752 1725
rect 29700 1673 29752 1698
rect 29700 1660 29752 1661
rect 29700 1626 29709 1660
rect 29709 1626 29743 1660
rect 29743 1626 29752 1660
rect 29700 1609 29752 1626
rect 29700 1588 29752 1597
rect 29700 1554 29709 1588
rect 29709 1554 29743 1588
rect 29743 1554 29752 1588
rect 29700 1545 29752 1554
rect 29700 1516 29752 1533
rect 29700 1482 29709 1516
rect 29709 1482 29743 1516
rect 29743 1482 29752 1516
rect 29700 1481 29752 1482
rect 29700 1444 29752 1469
rect 29700 1417 29709 1444
rect 29709 1417 29743 1444
rect 29743 1417 29752 1444
rect 29700 1372 29752 1405
rect 29700 1353 29709 1372
rect 29709 1353 29743 1372
rect 29743 1353 29752 1372
rect 29700 1338 29709 1341
rect 29709 1338 29743 1341
rect 29743 1338 29752 1341
rect 29700 1300 29752 1338
rect 29700 1289 29709 1300
rect 29709 1289 29743 1300
rect 29743 1289 29752 1300
rect 29700 1266 29709 1277
rect 29709 1266 29743 1277
rect 29743 1266 29752 1277
rect 29700 1228 29752 1266
rect 29700 1225 29709 1228
rect 29709 1225 29743 1228
rect 29743 1225 29752 1228
rect 29700 1194 29709 1213
rect 29709 1194 29743 1213
rect 29743 1194 29752 1213
rect 29700 1161 29752 1194
rect 29796 3100 29848 3133
rect 29796 3081 29805 3100
rect 29805 3081 29839 3100
rect 29839 3081 29848 3100
rect 29796 3066 29805 3069
rect 29805 3066 29839 3069
rect 29839 3066 29848 3069
rect 29796 3028 29848 3066
rect 29796 3017 29805 3028
rect 29805 3017 29839 3028
rect 29839 3017 29848 3028
rect 29796 2994 29805 3005
rect 29805 2994 29839 3005
rect 29839 2994 29848 3005
rect 29796 2956 29848 2994
rect 29796 2953 29805 2956
rect 29805 2953 29839 2956
rect 29839 2953 29848 2956
rect 29796 2922 29805 2941
rect 29805 2922 29839 2941
rect 29839 2922 29848 2941
rect 29796 2889 29848 2922
rect 29796 2850 29805 2877
rect 29805 2850 29839 2877
rect 29839 2850 29848 2877
rect 29796 2825 29848 2850
rect 29796 2812 29848 2813
rect 29796 2778 29805 2812
rect 29805 2778 29839 2812
rect 29839 2778 29848 2812
rect 29796 2761 29848 2778
rect 29796 2740 29848 2749
rect 29796 2706 29805 2740
rect 29805 2706 29839 2740
rect 29839 2706 29848 2740
rect 29796 2697 29848 2706
rect 29796 2668 29848 2685
rect 29796 2634 29805 2668
rect 29805 2634 29839 2668
rect 29839 2634 29848 2668
rect 29796 2633 29848 2634
rect 29796 2596 29848 2621
rect 29796 2569 29805 2596
rect 29805 2569 29839 2596
rect 29839 2569 29848 2596
rect 29796 2524 29848 2557
rect 29796 2505 29805 2524
rect 29805 2505 29839 2524
rect 29839 2505 29848 2524
rect 29796 2490 29805 2493
rect 29805 2490 29839 2493
rect 29839 2490 29848 2493
rect 29796 2452 29848 2490
rect 29796 2441 29805 2452
rect 29805 2441 29839 2452
rect 29839 2441 29848 2452
rect 29796 2418 29805 2429
rect 29805 2418 29839 2429
rect 29839 2418 29848 2429
rect 29796 2380 29848 2418
rect 29796 2377 29805 2380
rect 29805 2377 29839 2380
rect 29839 2377 29848 2380
rect 29796 2346 29805 2365
rect 29805 2346 29839 2365
rect 29839 2346 29848 2365
rect 29796 2313 29848 2346
rect 29796 2274 29805 2301
rect 29805 2274 29839 2301
rect 29839 2274 29848 2301
rect 29796 2249 29848 2274
rect 29796 2236 29848 2237
rect 29796 2202 29805 2236
rect 29805 2202 29839 2236
rect 29839 2202 29848 2236
rect 29796 2185 29848 2202
rect 29796 2164 29848 2173
rect 29796 2130 29805 2164
rect 29805 2130 29839 2164
rect 29839 2130 29848 2164
rect 29796 2121 29848 2130
rect 29796 2092 29848 2109
rect 29796 2058 29805 2092
rect 29805 2058 29839 2092
rect 29839 2058 29848 2092
rect 29796 2057 29848 2058
rect 29796 2020 29848 2045
rect 29796 1993 29805 2020
rect 29805 1993 29839 2020
rect 29839 1993 29848 2020
rect 29796 1948 29848 1981
rect 29796 1929 29805 1948
rect 29805 1929 29839 1948
rect 29839 1929 29848 1948
rect 29796 1914 29805 1917
rect 29805 1914 29839 1917
rect 29839 1914 29848 1917
rect 29796 1876 29848 1914
rect 29796 1865 29805 1876
rect 29805 1865 29839 1876
rect 29839 1865 29848 1876
rect 29796 1842 29805 1853
rect 29805 1842 29839 1853
rect 29839 1842 29848 1853
rect 29796 1804 29848 1842
rect 29796 1801 29805 1804
rect 29805 1801 29839 1804
rect 29839 1801 29848 1804
rect 29796 1770 29805 1789
rect 29805 1770 29839 1789
rect 29839 1770 29848 1789
rect 29796 1737 29848 1770
rect 29796 1698 29805 1725
rect 29805 1698 29839 1725
rect 29839 1698 29848 1725
rect 29796 1673 29848 1698
rect 29796 1660 29848 1661
rect 29796 1626 29805 1660
rect 29805 1626 29839 1660
rect 29839 1626 29848 1660
rect 29796 1609 29848 1626
rect 29796 1588 29848 1597
rect 29796 1554 29805 1588
rect 29805 1554 29839 1588
rect 29839 1554 29848 1588
rect 29796 1545 29848 1554
rect 29796 1516 29848 1533
rect 29796 1482 29805 1516
rect 29805 1482 29839 1516
rect 29839 1482 29848 1516
rect 29796 1481 29848 1482
rect 29796 1444 29848 1469
rect 29796 1417 29805 1444
rect 29805 1417 29839 1444
rect 29839 1417 29848 1444
rect 29796 1372 29848 1405
rect 29796 1353 29805 1372
rect 29805 1353 29839 1372
rect 29839 1353 29848 1372
rect 29796 1338 29805 1341
rect 29805 1338 29839 1341
rect 29839 1338 29848 1341
rect 29796 1300 29848 1338
rect 29796 1289 29805 1300
rect 29805 1289 29839 1300
rect 29839 1289 29848 1300
rect 29796 1266 29805 1277
rect 29805 1266 29839 1277
rect 29839 1266 29848 1277
rect 29796 1228 29848 1266
rect 29796 1225 29805 1228
rect 29805 1225 29839 1228
rect 29839 1225 29848 1228
rect 29796 1194 29805 1213
rect 29805 1194 29839 1213
rect 29839 1194 29848 1213
rect 29796 1161 29848 1194
rect 29892 3100 29944 3133
rect 29892 3081 29901 3100
rect 29901 3081 29935 3100
rect 29935 3081 29944 3100
rect 29892 3066 29901 3069
rect 29901 3066 29935 3069
rect 29935 3066 29944 3069
rect 29892 3028 29944 3066
rect 29892 3017 29901 3028
rect 29901 3017 29935 3028
rect 29935 3017 29944 3028
rect 29892 2994 29901 3005
rect 29901 2994 29935 3005
rect 29935 2994 29944 3005
rect 29892 2956 29944 2994
rect 29892 2953 29901 2956
rect 29901 2953 29935 2956
rect 29935 2953 29944 2956
rect 29892 2922 29901 2941
rect 29901 2922 29935 2941
rect 29935 2922 29944 2941
rect 29892 2889 29944 2922
rect 29892 2850 29901 2877
rect 29901 2850 29935 2877
rect 29935 2850 29944 2877
rect 29892 2825 29944 2850
rect 29892 2812 29944 2813
rect 29892 2778 29901 2812
rect 29901 2778 29935 2812
rect 29935 2778 29944 2812
rect 29892 2761 29944 2778
rect 29892 2740 29944 2749
rect 29892 2706 29901 2740
rect 29901 2706 29935 2740
rect 29935 2706 29944 2740
rect 29892 2697 29944 2706
rect 29892 2668 29944 2685
rect 29892 2634 29901 2668
rect 29901 2634 29935 2668
rect 29935 2634 29944 2668
rect 29892 2633 29944 2634
rect 29892 2596 29944 2621
rect 29892 2569 29901 2596
rect 29901 2569 29935 2596
rect 29935 2569 29944 2596
rect 29892 2524 29944 2557
rect 29892 2505 29901 2524
rect 29901 2505 29935 2524
rect 29935 2505 29944 2524
rect 29892 2490 29901 2493
rect 29901 2490 29935 2493
rect 29935 2490 29944 2493
rect 29892 2452 29944 2490
rect 29892 2441 29901 2452
rect 29901 2441 29935 2452
rect 29935 2441 29944 2452
rect 29892 2418 29901 2429
rect 29901 2418 29935 2429
rect 29935 2418 29944 2429
rect 29892 2380 29944 2418
rect 29892 2377 29901 2380
rect 29901 2377 29935 2380
rect 29935 2377 29944 2380
rect 29892 2346 29901 2365
rect 29901 2346 29935 2365
rect 29935 2346 29944 2365
rect 29892 2313 29944 2346
rect 29892 2274 29901 2301
rect 29901 2274 29935 2301
rect 29935 2274 29944 2301
rect 29892 2249 29944 2274
rect 29892 2236 29944 2237
rect 29892 2202 29901 2236
rect 29901 2202 29935 2236
rect 29935 2202 29944 2236
rect 29892 2185 29944 2202
rect 29892 2164 29944 2173
rect 29892 2130 29901 2164
rect 29901 2130 29935 2164
rect 29935 2130 29944 2164
rect 29892 2121 29944 2130
rect 29892 2092 29944 2109
rect 29892 2058 29901 2092
rect 29901 2058 29935 2092
rect 29935 2058 29944 2092
rect 29892 2057 29944 2058
rect 29892 2020 29944 2045
rect 29892 1993 29901 2020
rect 29901 1993 29935 2020
rect 29935 1993 29944 2020
rect 29892 1948 29944 1981
rect 29892 1929 29901 1948
rect 29901 1929 29935 1948
rect 29935 1929 29944 1948
rect 29892 1914 29901 1917
rect 29901 1914 29935 1917
rect 29935 1914 29944 1917
rect 29892 1876 29944 1914
rect 29892 1865 29901 1876
rect 29901 1865 29935 1876
rect 29935 1865 29944 1876
rect 29892 1842 29901 1853
rect 29901 1842 29935 1853
rect 29935 1842 29944 1853
rect 29892 1804 29944 1842
rect 29892 1801 29901 1804
rect 29901 1801 29935 1804
rect 29935 1801 29944 1804
rect 29892 1770 29901 1789
rect 29901 1770 29935 1789
rect 29935 1770 29944 1789
rect 29892 1737 29944 1770
rect 29892 1698 29901 1725
rect 29901 1698 29935 1725
rect 29935 1698 29944 1725
rect 29892 1673 29944 1698
rect 29892 1660 29944 1661
rect 29892 1626 29901 1660
rect 29901 1626 29935 1660
rect 29935 1626 29944 1660
rect 29892 1609 29944 1626
rect 29892 1588 29944 1597
rect 29892 1554 29901 1588
rect 29901 1554 29935 1588
rect 29935 1554 29944 1588
rect 29892 1545 29944 1554
rect 29892 1516 29944 1533
rect 29892 1482 29901 1516
rect 29901 1482 29935 1516
rect 29935 1482 29944 1516
rect 29892 1481 29944 1482
rect 29892 1444 29944 1469
rect 29892 1417 29901 1444
rect 29901 1417 29935 1444
rect 29935 1417 29944 1444
rect 29892 1372 29944 1405
rect 29892 1353 29901 1372
rect 29901 1353 29935 1372
rect 29935 1353 29944 1372
rect 29892 1338 29901 1341
rect 29901 1338 29935 1341
rect 29935 1338 29944 1341
rect 29892 1300 29944 1338
rect 29892 1289 29901 1300
rect 29901 1289 29935 1300
rect 29935 1289 29944 1300
rect 29892 1266 29901 1277
rect 29901 1266 29935 1277
rect 29935 1266 29944 1277
rect 29892 1228 29944 1266
rect 29892 1225 29901 1228
rect 29901 1225 29935 1228
rect 29935 1225 29944 1228
rect 29892 1194 29901 1213
rect 29901 1194 29935 1213
rect 29935 1194 29944 1213
rect 29892 1161 29944 1194
rect 29988 3100 30040 3133
rect 29988 3081 29997 3100
rect 29997 3081 30031 3100
rect 30031 3081 30040 3100
rect 29988 3066 29997 3069
rect 29997 3066 30031 3069
rect 30031 3066 30040 3069
rect 29988 3028 30040 3066
rect 29988 3017 29997 3028
rect 29997 3017 30031 3028
rect 30031 3017 30040 3028
rect 29988 2994 29997 3005
rect 29997 2994 30031 3005
rect 30031 2994 30040 3005
rect 29988 2956 30040 2994
rect 29988 2953 29997 2956
rect 29997 2953 30031 2956
rect 30031 2953 30040 2956
rect 29988 2922 29997 2941
rect 29997 2922 30031 2941
rect 30031 2922 30040 2941
rect 29988 2889 30040 2922
rect 29988 2850 29997 2877
rect 29997 2850 30031 2877
rect 30031 2850 30040 2877
rect 29988 2825 30040 2850
rect 29988 2812 30040 2813
rect 29988 2778 29997 2812
rect 29997 2778 30031 2812
rect 30031 2778 30040 2812
rect 29988 2761 30040 2778
rect 29988 2740 30040 2749
rect 29988 2706 29997 2740
rect 29997 2706 30031 2740
rect 30031 2706 30040 2740
rect 29988 2697 30040 2706
rect 29988 2668 30040 2685
rect 29988 2634 29997 2668
rect 29997 2634 30031 2668
rect 30031 2634 30040 2668
rect 29988 2633 30040 2634
rect 29988 2596 30040 2621
rect 29988 2569 29997 2596
rect 29997 2569 30031 2596
rect 30031 2569 30040 2596
rect 29988 2524 30040 2557
rect 29988 2505 29997 2524
rect 29997 2505 30031 2524
rect 30031 2505 30040 2524
rect 29988 2490 29997 2493
rect 29997 2490 30031 2493
rect 30031 2490 30040 2493
rect 29988 2452 30040 2490
rect 29988 2441 29997 2452
rect 29997 2441 30031 2452
rect 30031 2441 30040 2452
rect 29988 2418 29997 2429
rect 29997 2418 30031 2429
rect 30031 2418 30040 2429
rect 29988 2380 30040 2418
rect 29988 2377 29997 2380
rect 29997 2377 30031 2380
rect 30031 2377 30040 2380
rect 29988 2346 29997 2365
rect 29997 2346 30031 2365
rect 30031 2346 30040 2365
rect 29988 2313 30040 2346
rect 29988 2274 29997 2301
rect 29997 2274 30031 2301
rect 30031 2274 30040 2301
rect 29988 2249 30040 2274
rect 29988 2236 30040 2237
rect 29988 2202 29997 2236
rect 29997 2202 30031 2236
rect 30031 2202 30040 2236
rect 29988 2185 30040 2202
rect 29988 2164 30040 2173
rect 29988 2130 29997 2164
rect 29997 2130 30031 2164
rect 30031 2130 30040 2164
rect 29988 2121 30040 2130
rect 29988 2092 30040 2109
rect 29988 2058 29997 2092
rect 29997 2058 30031 2092
rect 30031 2058 30040 2092
rect 29988 2057 30040 2058
rect 29988 2020 30040 2045
rect 29988 1993 29997 2020
rect 29997 1993 30031 2020
rect 30031 1993 30040 2020
rect 29988 1948 30040 1981
rect 29988 1929 29997 1948
rect 29997 1929 30031 1948
rect 30031 1929 30040 1948
rect 29988 1914 29997 1917
rect 29997 1914 30031 1917
rect 30031 1914 30040 1917
rect 29988 1876 30040 1914
rect 29988 1865 29997 1876
rect 29997 1865 30031 1876
rect 30031 1865 30040 1876
rect 29988 1842 29997 1853
rect 29997 1842 30031 1853
rect 30031 1842 30040 1853
rect 29988 1804 30040 1842
rect 29988 1801 29997 1804
rect 29997 1801 30031 1804
rect 30031 1801 30040 1804
rect 29988 1770 29997 1789
rect 29997 1770 30031 1789
rect 30031 1770 30040 1789
rect 29988 1737 30040 1770
rect 29988 1698 29997 1725
rect 29997 1698 30031 1725
rect 30031 1698 30040 1725
rect 29988 1673 30040 1698
rect 29988 1660 30040 1661
rect 29988 1626 29997 1660
rect 29997 1626 30031 1660
rect 30031 1626 30040 1660
rect 29988 1609 30040 1626
rect 29988 1588 30040 1597
rect 29988 1554 29997 1588
rect 29997 1554 30031 1588
rect 30031 1554 30040 1588
rect 29988 1545 30040 1554
rect 29988 1516 30040 1533
rect 29988 1482 29997 1516
rect 29997 1482 30031 1516
rect 30031 1482 30040 1516
rect 29988 1481 30040 1482
rect 29988 1444 30040 1469
rect 29988 1417 29997 1444
rect 29997 1417 30031 1444
rect 30031 1417 30040 1444
rect 29988 1372 30040 1405
rect 29988 1353 29997 1372
rect 29997 1353 30031 1372
rect 30031 1353 30040 1372
rect 29988 1338 29997 1341
rect 29997 1338 30031 1341
rect 30031 1338 30040 1341
rect 29988 1300 30040 1338
rect 29988 1289 29997 1300
rect 29997 1289 30031 1300
rect 30031 1289 30040 1300
rect 29988 1266 29997 1277
rect 29997 1266 30031 1277
rect 30031 1266 30040 1277
rect 29988 1228 30040 1266
rect 29988 1225 29997 1228
rect 29997 1225 30031 1228
rect 30031 1225 30040 1228
rect 29988 1194 29997 1213
rect 29997 1194 30031 1213
rect 30031 1194 30040 1213
rect 29988 1161 30040 1194
rect 30084 3100 30136 3133
rect 30084 3081 30093 3100
rect 30093 3081 30127 3100
rect 30127 3081 30136 3100
rect 30084 3066 30093 3069
rect 30093 3066 30127 3069
rect 30127 3066 30136 3069
rect 30084 3028 30136 3066
rect 30084 3017 30093 3028
rect 30093 3017 30127 3028
rect 30127 3017 30136 3028
rect 30084 2994 30093 3005
rect 30093 2994 30127 3005
rect 30127 2994 30136 3005
rect 30084 2956 30136 2994
rect 30084 2953 30093 2956
rect 30093 2953 30127 2956
rect 30127 2953 30136 2956
rect 30084 2922 30093 2941
rect 30093 2922 30127 2941
rect 30127 2922 30136 2941
rect 30084 2889 30136 2922
rect 30084 2850 30093 2877
rect 30093 2850 30127 2877
rect 30127 2850 30136 2877
rect 30084 2825 30136 2850
rect 30084 2812 30136 2813
rect 30084 2778 30093 2812
rect 30093 2778 30127 2812
rect 30127 2778 30136 2812
rect 30084 2761 30136 2778
rect 30084 2740 30136 2749
rect 30084 2706 30093 2740
rect 30093 2706 30127 2740
rect 30127 2706 30136 2740
rect 30084 2697 30136 2706
rect 30084 2668 30136 2685
rect 30084 2634 30093 2668
rect 30093 2634 30127 2668
rect 30127 2634 30136 2668
rect 30084 2633 30136 2634
rect 30084 2596 30136 2621
rect 30084 2569 30093 2596
rect 30093 2569 30127 2596
rect 30127 2569 30136 2596
rect 30084 2524 30136 2557
rect 30084 2505 30093 2524
rect 30093 2505 30127 2524
rect 30127 2505 30136 2524
rect 30084 2490 30093 2493
rect 30093 2490 30127 2493
rect 30127 2490 30136 2493
rect 30084 2452 30136 2490
rect 30084 2441 30093 2452
rect 30093 2441 30127 2452
rect 30127 2441 30136 2452
rect 30084 2418 30093 2429
rect 30093 2418 30127 2429
rect 30127 2418 30136 2429
rect 30084 2380 30136 2418
rect 30084 2377 30093 2380
rect 30093 2377 30127 2380
rect 30127 2377 30136 2380
rect 30084 2346 30093 2365
rect 30093 2346 30127 2365
rect 30127 2346 30136 2365
rect 30084 2313 30136 2346
rect 30084 2274 30093 2301
rect 30093 2274 30127 2301
rect 30127 2274 30136 2301
rect 30084 2249 30136 2274
rect 30084 2236 30136 2237
rect 30084 2202 30093 2236
rect 30093 2202 30127 2236
rect 30127 2202 30136 2236
rect 30084 2185 30136 2202
rect 30084 2164 30136 2173
rect 30084 2130 30093 2164
rect 30093 2130 30127 2164
rect 30127 2130 30136 2164
rect 30084 2121 30136 2130
rect 30084 2092 30136 2109
rect 30084 2058 30093 2092
rect 30093 2058 30127 2092
rect 30127 2058 30136 2092
rect 30084 2057 30136 2058
rect 30084 2020 30136 2045
rect 30084 1993 30093 2020
rect 30093 1993 30127 2020
rect 30127 1993 30136 2020
rect 30084 1948 30136 1981
rect 30084 1929 30093 1948
rect 30093 1929 30127 1948
rect 30127 1929 30136 1948
rect 30084 1914 30093 1917
rect 30093 1914 30127 1917
rect 30127 1914 30136 1917
rect 30084 1876 30136 1914
rect 30084 1865 30093 1876
rect 30093 1865 30127 1876
rect 30127 1865 30136 1876
rect 30084 1842 30093 1853
rect 30093 1842 30127 1853
rect 30127 1842 30136 1853
rect 30084 1804 30136 1842
rect 30084 1801 30093 1804
rect 30093 1801 30127 1804
rect 30127 1801 30136 1804
rect 30084 1770 30093 1789
rect 30093 1770 30127 1789
rect 30127 1770 30136 1789
rect 30084 1737 30136 1770
rect 30084 1698 30093 1725
rect 30093 1698 30127 1725
rect 30127 1698 30136 1725
rect 30084 1673 30136 1698
rect 30084 1660 30136 1661
rect 30084 1626 30093 1660
rect 30093 1626 30127 1660
rect 30127 1626 30136 1660
rect 30084 1609 30136 1626
rect 30084 1588 30136 1597
rect 30084 1554 30093 1588
rect 30093 1554 30127 1588
rect 30127 1554 30136 1588
rect 30084 1545 30136 1554
rect 30084 1516 30136 1533
rect 30084 1482 30093 1516
rect 30093 1482 30127 1516
rect 30127 1482 30136 1516
rect 30084 1481 30136 1482
rect 30084 1444 30136 1469
rect 30084 1417 30093 1444
rect 30093 1417 30127 1444
rect 30127 1417 30136 1444
rect 30084 1372 30136 1405
rect 30084 1353 30093 1372
rect 30093 1353 30127 1372
rect 30127 1353 30136 1372
rect 30084 1338 30093 1341
rect 30093 1338 30127 1341
rect 30127 1338 30136 1341
rect 30084 1300 30136 1338
rect 30084 1289 30093 1300
rect 30093 1289 30127 1300
rect 30127 1289 30136 1300
rect 30084 1266 30093 1277
rect 30093 1266 30127 1277
rect 30127 1266 30136 1277
rect 30084 1228 30136 1266
rect 30084 1225 30093 1228
rect 30093 1225 30127 1228
rect 30127 1225 30136 1228
rect 30084 1194 30093 1213
rect 30093 1194 30127 1213
rect 30127 1194 30136 1213
rect 30084 1161 30136 1194
rect 30180 3100 30232 3133
rect 30180 3081 30189 3100
rect 30189 3081 30223 3100
rect 30223 3081 30232 3100
rect 30180 3066 30189 3069
rect 30189 3066 30223 3069
rect 30223 3066 30232 3069
rect 30180 3028 30232 3066
rect 30180 3017 30189 3028
rect 30189 3017 30223 3028
rect 30223 3017 30232 3028
rect 30180 2994 30189 3005
rect 30189 2994 30223 3005
rect 30223 2994 30232 3005
rect 30180 2956 30232 2994
rect 30180 2953 30189 2956
rect 30189 2953 30223 2956
rect 30223 2953 30232 2956
rect 30180 2922 30189 2941
rect 30189 2922 30223 2941
rect 30223 2922 30232 2941
rect 30180 2889 30232 2922
rect 30180 2850 30189 2877
rect 30189 2850 30223 2877
rect 30223 2850 30232 2877
rect 30180 2825 30232 2850
rect 30180 2812 30232 2813
rect 30180 2778 30189 2812
rect 30189 2778 30223 2812
rect 30223 2778 30232 2812
rect 30180 2761 30232 2778
rect 30180 2740 30232 2749
rect 30180 2706 30189 2740
rect 30189 2706 30223 2740
rect 30223 2706 30232 2740
rect 30180 2697 30232 2706
rect 30180 2668 30232 2685
rect 30180 2634 30189 2668
rect 30189 2634 30223 2668
rect 30223 2634 30232 2668
rect 30180 2633 30232 2634
rect 30180 2596 30232 2621
rect 30180 2569 30189 2596
rect 30189 2569 30223 2596
rect 30223 2569 30232 2596
rect 30180 2524 30232 2557
rect 30180 2505 30189 2524
rect 30189 2505 30223 2524
rect 30223 2505 30232 2524
rect 30180 2490 30189 2493
rect 30189 2490 30223 2493
rect 30223 2490 30232 2493
rect 30180 2452 30232 2490
rect 30180 2441 30189 2452
rect 30189 2441 30223 2452
rect 30223 2441 30232 2452
rect 30180 2418 30189 2429
rect 30189 2418 30223 2429
rect 30223 2418 30232 2429
rect 30180 2380 30232 2418
rect 30180 2377 30189 2380
rect 30189 2377 30223 2380
rect 30223 2377 30232 2380
rect 30180 2346 30189 2365
rect 30189 2346 30223 2365
rect 30223 2346 30232 2365
rect 30180 2313 30232 2346
rect 30180 2274 30189 2301
rect 30189 2274 30223 2301
rect 30223 2274 30232 2301
rect 30180 2249 30232 2274
rect 30180 2236 30232 2237
rect 30180 2202 30189 2236
rect 30189 2202 30223 2236
rect 30223 2202 30232 2236
rect 30180 2185 30232 2202
rect 30180 2164 30232 2173
rect 30180 2130 30189 2164
rect 30189 2130 30223 2164
rect 30223 2130 30232 2164
rect 30180 2121 30232 2130
rect 30180 2092 30232 2109
rect 30180 2058 30189 2092
rect 30189 2058 30223 2092
rect 30223 2058 30232 2092
rect 30180 2057 30232 2058
rect 30180 2020 30232 2045
rect 30180 1993 30189 2020
rect 30189 1993 30223 2020
rect 30223 1993 30232 2020
rect 30180 1948 30232 1981
rect 30180 1929 30189 1948
rect 30189 1929 30223 1948
rect 30223 1929 30232 1948
rect 30180 1914 30189 1917
rect 30189 1914 30223 1917
rect 30223 1914 30232 1917
rect 30180 1876 30232 1914
rect 30180 1865 30189 1876
rect 30189 1865 30223 1876
rect 30223 1865 30232 1876
rect 30180 1842 30189 1853
rect 30189 1842 30223 1853
rect 30223 1842 30232 1853
rect 30180 1804 30232 1842
rect 30180 1801 30189 1804
rect 30189 1801 30223 1804
rect 30223 1801 30232 1804
rect 30180 1770 30189 1789
rect 30189 1770 30223 1789
rect 30223 1770 30232 1789
rect 30180 1737 30232 1770
rect 30180 1698 30189 1725
rect 30189 1698 30223 1725
rect 30223 1698 30232 1725
rect 30180 1673 30232 1698
rect 30180 1660 30232 1661
rect 30180 1626 30189 1660
rect 30189 1626 30223 1660
rect 30223 1626 30232 1660
rect 30180 1609 30232 1626
rect 30180 1588 30232 1597
rect 30180 1554 30189 1588
rect 30189 1554 30223 1588
rect 30223 1554 30232 1588
rect 30180 1545 30232 1554
rect 30180 1516 30232 1533
rect 30180 1482 30189 1516
rect 30189 1482 30223 1516
rect 30223 1482 30232 1516
rect 30180 1481 30232 1482
rect 30180 1444 30232 1469
rect 30180 1417 30189 1444
rect 30189 1417 30223 1444
rect 30223 1417 30232 1444
rect 30180 1372 30232 1405
rect 30180 1353 30189 1372
rect 30189 1353 30223 1372
rect 30223 1353 30232 1372
rect 30180 1338 30189 1341
rect 30189 1338 30223 1341
rect 30223 1338 30232 1341
rect 30180 1300 30232 1338
rect 30180 1289 30189 1300
rect 30189 1289 30223 1300
rect 30223 1289 30232 1300
rect 30180 1266 30189 1277
rect 30189 1266 30223 1277
rect 30223 1266 30232 1277
rect 30180 1228 30232 1266
rect 30180 1225 30189 1228
rect 30189 1225 30223 1228
rect 30223 1225 30232 1228
rect 30180 1194 30189 1213
rect 30189 1194 30223 1213
rect 30223 1194 30232 1213
rect 30180 1161 30232 1194
rect 30276 3100 30328 3133
rect 30276 3081 30285 3100
rect 30285 3081 30319 3100
rect 30319 3081 30328 3100
rect 30276 3066 30285 3069
rect 30285 3066 30319 3069
rect 30319 3066 30328 3069
rect 30276 3028 30328 3066
rect 30276 3017 30285 3028
rect 30285 3017 30319 3028
rect 30319 3017 30328 3028
rect 30276 2994 30285 3005
rect 30285 2994 30319 3005
rect 30319 2994 30328 3005
rect 30276 2956 30328 2994
rect 30276 2953 30285 2956
rect 30285 2953 30319 2956
rect 30319 2953 30328 2956
rect 30276 2922 30285 2941
rect 30285 2922 30319 2941
rect 30319 2922 30328 2941
rect 30276 2889 30328 2922
rect 30276 2850 30285 2877
rect 30285 2850 30319 2877
rect 30319 2850 30328 2877
rect 30276 2825 30328 2850
rect 30276 2812 30328 2813
rect 30276 2778 30285 2812
rect 30285 2778 30319 2812
rect 30319 2778 30328 2812
rect 30276 2761 30328 2778
rect 30276 2740 30328 2749
rect 30276 2706 30285 2740
rect 30285 2706 30319 2740
rect 30319 2706 30328 2740
rect 30276 2697 30328 2706
rect 30276 2668 30328 2685
rect 30276 2634 30285 2668
rect 30285 2634 30319 2668
rect 30319 2634 30328 2668
rect 30276 2633 30328 2634
rect 30276 2596 30328 2621
rect 30276 2569 30285 2596
rect 30285 2569 30319 2596
rect 30319 2569 30328 2596
rect 30276 2524 30328 2557
rect 30276 2505 30285 2524
rect 30285 2505 30319 2524
rect 30319 2505 30328 2524
rect 30276 2490 30285 2493
rect 30285 2490 30319 2493
rect 30319 2490 30328 2493
rect 30276 2452 30328 2490
rect 30276 2441 30285 2452
rect 30285 2441 30319 2452
rect 30319 2441 30328 2452
rect 30276 2418 30285 2429
rect 30285 2418 30319 2429
rect 30319 2418 30328 2429
rect 30276 2380 30328 2418
rect 30276 2377 30285 2380
rect 30285 2377 30319 2380
rect 30319 2377 30328 2380
rect 30276 2346 30285 2365
rect 30285 2346 30319 2365
rect 30319 2346 30328 2365
rect 30276 2313 30328 2346
rect 30276 2274 30285 2301
rect 30285 2274 30319 2301
rect 30319 2274 30328 2301
rect 30276 2249 30328 2274
rect 30276 2236 30328 2237
rect 30276 2202 30285 2236
rect 30285 2202 30319 2236
rect 30319 2202 30328 2236
rect 30276 2185 30328 2202
rect 30276 2164 30328 2173
rect 30276 2130 30285 2164
rect 30285 2130 30319 2164
rect 30319 2130 30328 2164
rect 30276 2121 30328 2130
rect 30276 2092 30328 2109
rect 30276 2058 30285 2092
rect 30285 2058 30319 2092
rect 30319 2058 30328 2092
rect 30276 2057 30328 2058
rect 30276 2020 30328 2045
rect 30276 1993 30285 2020
rect 30285 1993 30319 2020
rect 30319 1993 30328 2020
rect 30276 1948 30328 1981
rect 30276 1929 30285 1948
rect 30285 1929 30319 1948
rect 30319 1929 30328 1948
rect 30276 1914 30285 1917
rect 30285 1914 30319 1917
rect 30319 1914 30328 1917
rect 30276 1876 30328 1914
rect 30276 1865 30285 1876
rect 30285 1865 30319 1876
rect 30319 1865 30328 1876
rect 30276 1842 30285 1853
rect 30285 1842 30319 1853
rect 30319 1842 30328 1853
rect 30276 1804 30328 1842
rect 30276 1801 30285 1804
rect 30285 1801 30319 1804
rect 30319 1801 30328 1804
rect 30276 1770 30285 1789
rect 30285 1770 30319 1789
rect 30319 1770 30328 1789
rect 30276 1737 30328 1770
rect 30276 1698 30285 1725
rect 30285 1698 30319 1725
rect 30319 1698 30328 1725
rect 30276 1673 30328 1698
rect 30276 1660 30328 1661
rect 30276 1626 30285 1660
rect 30285 1626 30319 1660
rect 30319 1626 30328 1660
rect 30276 1609 30328 1626
rect 30276 1588 30328 1597
rect 30276 1554 30285 1588
rect 30285 1554 30319 1588
rect 30319 1554 30328 1588
rect 30276 1545 30328 1554
rect 30276 1516 30328 1533
rect 30276 1482 30285 1516
rect 30285 1482 30319 1516
rect 30319 1482 30328 1516
rect 30276 1481 30328 1482
rect 30276 1444 30328 1469
rect 30276 1417 30285 1444
rect 30285 1417 30319 1444
rect 30319 1417 30328 1444
rect 30276 1372 30328 1405
rect 30276 1353 30285 1372
rect 30285 1353 30319 1372
rect 30319 1353 30328 1372
rect 30276 1338 30285 1341
rect 30285 1338 30319 1341
rect 30319 1338 30328 1341
rect 30276 1300 30328 1338
rect 30276 1289 30285 1300
rect 30285 1289 30319 1300
rect 30319 1289 30328 1300
rect 30276 1266 30285 1277
rect 30285 1266 30319 1277
rect 30319 1266 30328 1277
rect 30276 1228 30328 1266
rect 30276 1225 30285 1228
rect 30285 1225 30319 1228
rect 30319 1225 30328 1228
rect 30276 1194 30285 1213
rect 30285 1194 30319 1213
rect 30319 1194 30328 1213
rect 30276 1161 30328 1194
rect 30372 3100 30424 3133
rect 30372 3081 30381 3100
rect 30381 3081 30415 3100
rect 30415 3081 30424 3100
rect 30372 3066 30381 3069
rect 30381 3066 30415 3069
rect 30415 3066 30424 3069
rect 30372 3028 30424 3066
rect 30372 3017 30381 3028
rect 30381 3017 30415 3028
rect 30415 3017 30424 3028
rect 30372 2994 30381 3005
rect 30381 2994 30415 3005
rect 30415 2994 30424 3005
rect 30372 2956 30424 2994
rect 30372 2953 30381 2956
rect 30381 2953 30415 2956
rect 30415 2953 30424 2956
rect 30372 2922 30381 2941
rect 30381 2922 30415 2941
rect 30415 2922 30424 2941
rect 30372 2889 30424 2922
rect 30372 2850 30381 2877
rect 30381 2850 30415 2877
rect 30415 2850 30424 2877
rect 30372 2825 30424 2850
rect 30372 2812 30424 2813
rect 30372 2778 30381 2812
rect 30381 2778 30415 2812
rect 30415 2778 30424 2812
rect 30372 2761 30424 2778
rect 30372 2740 30424 2749
rect 30372 2706 30381 2740
rect 30381 2706 30415 2740
rect 30415 2706 30424 2740
rect 30372 2697 30424 2706
rect 30372 2668 30424 2685
rect 30372 2634 30381 2668
rect 30381 2634 30415 2668
rect 30415 2634 30424 2668
rect 30372 2633 30424 2634
rect 30372 2596 30424 2621
rect 30372 2569 30381 2596
rect 30381 2569 30415 2596
rect 30415 2569 30424 2596
rect 30372 2524 30424 2557
rect 30372 2505 30381 2524
rect 30381 2505 30415 2524
rect 30415 2505 30424 2524
rect 30372 2490 30381 2493
rect 30381 2490 30415 2493
rect 30415 2490 30424 2493
rect 30372 2452 30424 2490
rect 30372 2441 30381 2452
rect 30381 2441 30415 2452
rect 30415 2441 30424 2452
rect 30372 2418 30381 2429
rect 30381 2418 30415 2429
rect 30415 2418 30424 2429
rect 30372 2380 30424 2418
rect 30372 2377 30381 2380
rect 30381 2377 30415 2380
rect 30415 2377 30424 2380
rect 30372 2346 30381 2365
rect 30381 2346 30415 2365
rect 30415 2346 30424 2365
rect 30372 2313 30424 2346
rect 30372 2274 30381 2301
rect 30381 2274 30415 2301
rect 30415 2274 30424 2301
rect 30372 2249 30424 2274
rect 30372 2236 30424 2237
rect 30372 2202 30381 2236
rect 30381 2202 30415 2236
rect 30415 2202 30424 2236
rect 30372 2185 30424 2202
rect 30372 2164 30424 2173
rect 30372 2130 30381 2164
rect 30381 2130 30415 2164
rect 30415 2130 30424 2164
rect 30372 2121 30424 2130
rect 30372 2092 30424 2109
rect 30372 2058 30381 2092
rect 30381 2058 30415 2092
rect 30415 2058 30424 2092
rect 30372 2057 30424 2058
rect 30372 2020 30424 2045
rect 30372 1993 30381 2020
rect 30381 1993 30415 2020
rect 30415 1993 30424 2020
rect 30372 1948 30424 1981
rect 30372 1929 30381 1948
rect 30381 1929 30415 1948
rect 30415 1929 30424 1948
rect 30372 1914 30381 1917
rect 30381 1914 30415 1917
rect 30415 1914 30424 1917
rect 30372 1876 30424 1914
rect 30372 1865 30381 1876
rect 30381 1865 30415 1876
rect 30415 1865 30424 1876
rect 30372 1842 30381 1853
rect 30381 1842 30415 1853
rect 30415 1842 30424 1853
rect 30372 1804 30424 1842
rect 30372 1801 30381 1804
rect 30381 1801 30415 1804
rect 30415 1801 30424 1804
rect 30372 1770 30381 1789
rect 30381 1770 30415 1789
rect 30415 1770 30424 1789
rect 30372 1737 30424 1770
rect 30372 1698 30381 1725
rect 30381 1698 30415 1725
rect 30415 1698 30424 1725
rect 30372 1673 30424 1698
rect 30372 1660 30424 1661
rect 30372 1626 30381 1660
rect 30381 1626 30415 1660
rect 30415 1626 30424 1660
rect 30372 1609 30424 1626
rect 30372 1588 30424 1597
rect 30372 1554 30381 1588
rect 30381 1554 30415 1588
rect 30415 1554 30424 1588
rect 30372 1545 30424 1554
rect 30372 1516 30424 1533
rect 30372 1482 30381 1516
rect 30381 1482 30415 1516
rect 30415 1482 30424 1516
rect 30372 1481 30424 1482
rect 30372 1444 30424 1469
rect 30372 1417 30381 1444
rect 30381 1417 30415 1444
rect 30415 1417 30424 1444
rect 30372 1372 30424 1405
rect 30372 1353 30381 1372
rect 30381 1353 30415 1372
rect 30415 1353 30424 1372
rect 30372 1338 30381 1341
rect 30381 1338 30415 1341
rect 30415 1338 30424 1341
rect 30372 1300 30424 1338
rect 30372 1289 30381 1300
rect 30381 1289 30415 1300
rect 30415 1289 30424 1300
rect 30372 1266 30381 1277
rect 30381 1266 30415 1277
rect 30415 1266 30424 1277
rect 30372 1228 30424 1266
rect 30372 1225 30381 1228
rect 30381 1225 30415 1228
rect 30415 1225 30424 1228
rect 30372 1194 30381 1213
rect 30381 1194 30415 1213
rect 30415 1194 30424 1213
rect 30372 1161 30424 1194
rect 30468 3100 30520 3133
rect 30468 3081 30477 3100
rect 30477 3081 30511 3100
rect 30511 3081 30520 3100
rect 30468 3066 30477 3069
rect 30477 3066 30511 3069
rect 30511 3066 30520 3069
rect 30468 3028 30520 3066
rect 30468 3017 30477 3028
rect 30477 3017 30511 3028
rect 30511 3017 30520 3028
rect 30468 2994 30477 3005
rect 30477 2994 30511 3005
rect 30511 2994 30520 3005
rect 30468 2956 30520 2994
rect 30468 2953 30477 2956
rect 30477 2953 30511 2956
rect 30511 2953 30520 2956
rect 30468 2922 30477 2941
rect 30477 2922 30511 2941
rect 30511 2922 30520 2941
rect 30468 2889 30520 2922
rect 30468 2850 30477 2877
rect 30477 2850 30511 2877
rect 30511 2850 30520 2877
rect 30468 2825 30520 2850
rect 30468 2812 30520 2813
rect 30468 2778 30477 2812
rect 30477 2778 30511 2812
rect 30511 2778 30520 2812
rect 30468 2761 30520 2778
rect 30468 2740 30520 2749
rect 30468 2706 30477 2740
rect 30477 2706 30511 2740
rect 30511 2706 30520 2740
rect 30468 2697 30520 2706
rect 30468 2668 30520 2685
rect 30468 2634 30477 2668
rect 30477 2634 30511 2668
rect 30511 2634 30520 2668
rect 30468 2633 30520 2634
rect 30468 2596 30520 2621
rect 30468 2569 30477 2596
rect 30477 2569 30511 2596
rect 30511 2569 30520 2596
rect 30468 2524 30520 2557
rect 30468 2505 30477 2524
rect 30477 2505 30511 2524
rect 30511 2505 30520 2524
rect 30468 2490 30477 2493
rect 30477 2490 30511 2493
rect 30511 2490 30520 2493
rect 30468 2452 30520 2490
rect 30468 2441 30477 2452
rect 30477 2441 30511 2452
rect 30511 2441 30520 2452
rect 30468 2418 30477 2429
rect 30477 2418 30511 2429
rect 30511 2418 30520 2429
rect 30468 2380 30520 2418
rect 30468 2377 30477 2380
rect 30477 2377 30511 2380
rect 30511 2377 30520 2380
rect 30468 2346 30477 2365
rect 30477 2346 30511 2365
rect 30511 2346 30520 2365
rect 30468 2313 30520 2346
rect 30468 2274 30477 2301
rect 30477 2274 30511 2301
rect 30511 2274 30520 2301
rect 30468 2249 30520 2274
rect 30468 2236 30520 2237
rect 30468 2202 30477 2236
rect 30477 2202 30511 2236
rect 30511 2202 30520 2236
rect 30468 2185 30520 2202
rect 30468 2164 30520 2173
rect 30468 2130 30477 2164
rect 30477 2130 30511 2164
rect 30511 2130 30520 2164
rect 30468 2121 30520 2130
rect 30468 2092 30520 2109
rect 30468 2058 30477 2092
rect 30477 2058 30511 2092
rect 30511 2058 30520 2092
rect 30468 2057 30520 2058
rect 30468 2020 30520 2045
rect 30468 1993 30477 2020
rect 30477 1993 30511 2020
rect 30511 1993 30520 2020
rect 30468 1948 30520 1981
rect 30468 1929 30477 1948
rect 30477 1929 30511 1948
rect 30511 1929 30520 1948
rect 30468 1914 30477 1917
rect 30477 1914 30511 1917
rect 30511 1914 30520 1917
rect 30468 1876 30520 1914
rect 30468 1865 30477 1876
rect 30477 1865 30511 1876
rect 30511 1865 30520 1876
rect 30468 1842 30477 1853
rect 30477 1842 30511 1853
rect 30511 1842 30520 1853
rect 30468 1804 30520 1842
rect 30468 1801 30477 1804
rect 30477 1801 30511 1804
rect 30511 1801 30520 1804
rect 30468 1770 30477 1789
rect 30477 1770 30511 1789
rect 30511 1770 30520 1789
rect 30468 1737 30520 1770
rect 30468 1698 30477 1725
rect 30477 1698 30511 1725
rect 30511 1698 30520 1725
rect 30468 1673 30520 1698
rect 30468 1660 30520 1661
rect 30468 1626 30477 1660
rect 30477 1626 30511 1660
rect 30511 1626 30520 1660
rect 30468 1609 30520 1626
rect 30468 1588 30520 1597
rect 30468 1554 30477 1588
rect 30477 1554 30511 1588
rect 30511 1554 30520 1588
rect 30468 1545 30520 1554
rect 30468 1516 30520 1533
rect 30468 1482 30477 1516
rect 30477 1482 30511 1516
rect 30511 1482 30520 1516
rect 30468 1481 30520 1482
rect 30468 1444 30520 1469
rect 30468 1417 30477 1444
rect 30477 1417 30511 1444
rect 30511 1417 30520 1444
rect 30468 1372 30520 1405
rect 30468 1353 30477 1372
rect 30477 1353 30511 1372
rect 30511 1353 30520 1372
rect 30468 1338 30477 1341
rect 30477 1338 30511 1341
rect 30511 1338 30520 1341
rect 30468 1300 30520 1338
rect 30468 1289 30477 1300
rect 30477 1289 30511 1300
rect 30511 1289 30520 1300
rect 30468 1266 30477 1277
rect 30477 1266 30511 1277
rect 30511 1266 30520 1277
rect 30468 1228 30520 1266
rect 30468 1225 30477 1228
rect 30477 1225 30511 1228
rect 30511 1225 30520 1228
rect 30468 1194 30477 1213
rect 30477 1194 30511 1213
rect 30511 1194 30520 1213
rect 30468 1161 30520 1194
rect 30564 3100 30616 3133
rect 30564 3081 30573 3100
rect 30573 3081 30607 3100
rect 30607 3081 30616 3100
rect 30564 3066 30573 3069
rect 30573 3066 30607 3069
rect 30607 3066 30616 3069
rect 30564 3028 30616 3066
rect 30564 3017 30573 3028
rect 30573 3017 30607 3028
rect 30607 3017 30616 3028
rect 30564 2994 30573 3005
rect 30573 2994 30607 3005
rect 30607 2994 30616 3005
rect 30564 2956 30616 2994
rect 30564 2953 30573 2956
rect 30573 2953 30607 2956
rect 30607 2953 30616 2956
rect 30564 2922 30573 2941
rect 30573 2922 30607 2941
rect 30607 2922 30616 2941
rect 30564 2889 30616 2922
rect 30564 2850 30573 2877
rect 30573 2850 30607 2877
rect 30607 2850 30616 2877
rect 30564 2825 30616 2850
rect 30564 2812 30616 2813
rect 30564 2778 30573 2812
rect 30573 2778 30607 2812
rect 30607 2778 30616 2812
rect 30564 2761 30616 2778
rect 30564 2740 30616 2749
rect 30564 2706 30573 2740
rect 30573 2706 30607 2740
rect 30607 2706 30616 2740
rect 30564 2697 30616 2706
rect 30564 2668 30616 2685
rect 30564 2634 30573 2668
rect 30573 2634 30607 2668
rect 30607 2634 30616 2668
rect 30564 2633 30616 2634
rect 30564 2596 30616 2621
rect 30564 2569 30573 2596
rect 30573 2569 30607 2596
rect 30607 2569 30616 2596
rect 30564 2524 30616 2557
rect 30564 2505 30573 2524
rect 30573 2505 30607 2524
rect 30607 2505 30616 2524
rect 30564 2490 30573 2493
rect 30573 2490 30607 2493
rect 30607 2490 30616 2493
rect 30564 2452 30616 2490
rect 30564 2441 30573 2452
rect 30573 2441 30607 2452
rect 30607 2441 30616 2452
rect 30564 2418 30573 2429
rect 30573 2418 30607 2429
rect 30607 2418 30616 2429
rect 30564 2380 30616 2418
rect 30564 2377 30573 2380
rect 30573 2377 30607 2380
rect 30607 2377 30616 2380
rect 30564 2346 30573 2365
rect 30573 2346 30607 2365
rect 30607 2346 30616 2365
rect 30564 2313 30616 2346
rect 30564 2274 30573 2301
rect 30573 2274 30607 2301
rect 30607 2274 30616 2301
rect 30564 2249 30616 2274
rect 30564 2236 30616 2237
rect 30564 2202 30573 2236
rect 30573 2202 30607 2236
rect 30607 2202 30616 2236
rect 30564 2185 30616 2202
rect 30564 2164 30616 2173
rect 30564 2130 30573 2164
rect 30573 2130 30607 2164
rect 30607 2130 30616 2164
rect 30564 2121 30616 2130
rect 30564 2092 30616 2109
rect 30564 2058 30573 2092
rect 30573 2058 30607 2092
rect 30607 2058 30616 2092
rect 30564 2057 30616 2058
rect 30564 2020 30616 2045
rect 30564 1993 30573 2020
rect 30573 1993 30607 2020
rect 30607 1993 30616 2020
rect 30564 1948 30616 1981
rect 30564 1929 30573 1948
rect 30573 1929 30607 1948
rect 30607 1929 30616 1948
rect 30564 1914 30573 1917
rect 30573 1914 30607 1917
rect 30607 1914 30616 1917
rect 30564 1876 30616 1914
rect 30564 1865 30573 1876
rect 30573 1865 30607 1876
rect 30607 1865 30616 1876
rect 30564 1842 30573 1853
rect 30573 1842 30607 1853
rect 30607 1842 30616 1853
rect 30564 1804 30616 1842
rect 30564 1801 30573 1804
rect 30573 1801 30607 1804
rect 30607 1801 30616 1804
rect 30564 1770 30573 1789
rect 30573 1770 30607 1789
rect 30607 1770 30616 1789
rect 30564 1737 30616 1770
rect 30564 1698 30573 1725
rect 30573 1698 30607 1725
rect 30607 1698 30616 1725
rect 30564 1673 30616 1698
rect 30564 1660 30616 1661
rect 30564 1626 30573 1660
rect 30573 1626 30607 1660
rect 30607 1626 30616 1660
rect 30564 1609 30616 1626
rect 30564 1588 30616 1597
rect 30564 1554 30573 1588
rect 30573 1554 30607 1588
rect 30607 1554 30616 1588
rect 30564 1545 30616 1554
rect 30564 1516 30616 1533
rect 30564 1482 30573 1516
rect 30573 1482 30607 1516
rect 30607 1482 30616 1516
rect 30564 1481 30616 1482
rect 30564 1444 30616 1469
rect 30564 1417 30573 1444
rect 30573 1417 30607 1444
rect 30607 1417 30616 1444
rect 30564 1372 30616 1405
rect 30564 1353 30573 1372
rect 30573 1353 30607 1372
rect 30607 1353 30616 1372
rect 30564 1338 30573 1341
rect 30573 1338 30607 1341
rect 30607 1338 30616 1341
rect 30564 1300 30616 1338
rect 30564 1289 30573 1300
rect 30573 1289 30607 1300
rect 30607 1289 30616 1300
rect 30564 1266 30573 1277
rect 30573 1266 30607 1277
rect 30607 1266 30616 1277
rect 30564 1228 30616 1266
rect 30564 1225 30573 1228
rect 30573 1225 30607 1228
rect 30607 1225 30616 1228
rect 30564 1194 30573 1213
rect 30573 1194 30607 1213
rect 30607 1194 30616 1213
rect 30564 1161 30616 1194
rect 30660 3100 30712 3133
rect 30660 3081 30669 3100
rect 30669 3081 30703 3100
rect 30703 3081 30712 3100
rect 30660 3066 30669 3069
rect 30669 3066 30703 3069
rect 30703 3066 30712 3069
rect 30660 3028 30712 3066
rect 30660 3017 30669 3028
rect 30669 3017 30703 3028
rect 30703 3017 30712 3028
rect 30660 2994 30669 3005
rect 30669 2994 30703 3005
rect 30703 2994 30712 3005
rect 30660 2956 30712 2994
rect 30660 2953 30669 2956
rect 30669 2953 30703 2956
rect 30703 2953 30712 2956
rect 30660 2922 30669 2941
rect 30669 2922 30703 2941
rect 30703 2922 30712 2941
rect 30660 2889 30712 2922
rect 30660 2850 30669 2877
rect 30669 2850 30703 2877
rect 30703 2850 30712 2877
rect 30660 2825 30712 2850
rect 30660 2812 30712 2813
rect 30660 2778 30669 2812
rect 30669 2778 30703 2812
rect 30703 2778 30712 2812
rect 30660 2761 30712 2778
rect 30660 2740 30712 2749
rect 30660 2706 30669 2740
rect 30669 2706 30703 2740
rect 30703 2706 30712 2740
rect 30660 2697 30712 2706
rect 30660 2668 30712 2685
rect 30660 2634 30669 2668
rect 30669 2634 30703 2668
rect 30703 2634 30712 2668
rect 30660 2633 30712 2634
rect 30660 2596 30712 2621
rect 30660 2569 30669 2596
rect 30669 2569 30703 2596
rect 30703 2569 30712 2596
rect 30660 2524 30712 2557
rect 30660 2505 30669 2524
rect 30669 2505 30703 2524
rect 30703 2505 30712 2524
rect 30660 2490 30669 2493
rect 30669 2490 30703 2493
rect 30703 2490 30712 2493
rect 30660 2452 30712 2490
rect 30660 2441 30669 2452
rect 30669 2441 30703 2452
rect 30703 2441 30712 2452
rect 30660 2418 30669 2429
rect 30669 2418 30703 2429
rect 30703 2418 30712 2429
rect 30660 2380 30712 2418
rect 30660 2377 30669 2380
rect 30669 2377 30703 2380
rect 30703 2377 30712 2380
rect 30660 2346 30669 2365
rect 30669 2346 30703 2365
rect 30703 2346 30712 2365
rect 30660 2313 30712 2346
rect 30660 2274 30669 2301
rect 30669 2274 30703 2301
rect 30703 2274 30712 2301
rect 30660 2249 30712 2274
rect 30660 2236 30712 2237
rect 30660 2202 30669 2236
rect 30669 2202 30703 2236
rect 30703 2202 30712 2236
rect 30660 2185 30712 2202
rect 30660 2164 30712 2173
rect 30660 2130 30669 2164
rect 30669 2130 30703 2164
rect 30703 2130 30712 2164
rect 30660 2121 30712 2130
rect 30660 2092 30712 2109
rect 30660 2058 30669 2092
rect 30669 2058 30703 2092
rect 30703 2058 30712 2092
rect 30660 2057 30712 2058
rect 30660 2020 30712 2045
rect 30660 1993 30669 2020
rect 30669 1993 30703 2020
rect 30703 1993 30712 2020
rect 30660 1948 30712 1981
rect 30660 1929 30669 1948
rect 30669 1929 30703 1948
rect 30703 1929 30712 1948
rect 30660 1914 30669 1917
rect 30669 1914 30703 1917
rect 30703 1914 30712 1917
rect 30660 1876 30712 1914
rect 30660 1865 30669 1876
rect 30669 1865 30703 1876
rect 30703 1865 30712 1876
rect 30660 1842 30669 1853
rect 30669 1842 30703 1853
rect 30703 1842 30712 1853
rect 30660 1804 30712 1842
rect 30660 1801 30669 1804
rect 30669 1801 30703 1804
rect 30703 1801 30712 1804
rect 30660 1770 30669 1789
rect 30669 1770 30703 1789
rect 30703 1770 30712 1789
rect 30660 1737 30712 1770
rect 30660 1698 30669 1725
rect 30669 1698 30703 1725
rect 30703 1698 30712 1725
rect 30660 1673 30712 1698
rect 30660 1660 30712 1661
rect 30660 1626 30669 1660
rect 30669 1626 30703 1660
rect 30703 1626 30712 1660
rect 30660 1609 30712 1626
rect 30660 1588 30712 1597
rect 30660 1554 30669 1588
rect 30669 1554 30703 1588
rect 30703 1554 30712 1588
rect 30660 1545 30712 1554
rect 30660 1516 30712 1533
rect 30660 1482 30669 1516
rect 30669 1482 30703 1516
rect 30703 1482 30712 1516
rect 30660 1481 30712 1482
rect 30660 1444 30712 1469
rect 30660 1417 30669 1444
rect 30669 1417 30703 1444
rect 30703 1417 30712 1444
rect 30660 1372 30712 1405
rect 30660 1353 30669 1372
rect 30669 1353 30703 1372
rect 30703 1353 30712 1372
rect 30660 1338 30669 1341
rect 30669 1338 30703 1341
rect 30703 1338 30712 1341
rect 30660 1300 30712 1338
rect 30660 1289 30669 1300
rect 30669 1289 30703 1300
rect 30703 1289 30712 1300
rect 30660 1266 30669 1277
rect 30669 1266 30703 1277
rect 30703 1266 30712 1277
rect 30660 1228 30712 1266
rect 30660 1225 30669 1228
rect 30669 1225 30703 1228
rect 30703 1225 30712 1228
rect 30660 1194 30669 1213
rect 30669 1194 30703 1213
rect 30703 1194 30712 1213
rect 30660 1161 30712 1194
rect 30756 3100 30808 3133
rect 30756 3081 30765 3100
rect 30765 3081 30799 3100
rect 30799 3081 30808 3100
rect 30756 3066 30765 3069
rect 30765 3066 30799 3069
rect 30799 3066 30808 3069
rect 30756 3028 30808 3066
rect 30756 3017 30765 3028
rect 30765 3017 30799 3028
rect 30799 3017 30808 3028
rect 30756 2994 30765 3005
rect 30765 2994 30799 3005
rect 30799 2994 30808 3005
rect 30756 2956 30808 2994
rect 30756 2953 30765 2956
rect 30765 2953 30799 2956
rect 30799 2953 30808 2956
rect 30756 2922 30765 2941
rect 30765 2922 30799 2941
rect 30799 2922 30808 2941
rect 30756 2889 30808 2922
rect 30756 2850 30765 2877
rect 30765 2850 30799 2877
rect 30799 2850 30808 2877
rect 30756 2825 30808 2850
rect 30756 2812 30808 2813
rect 30756 2778 30765 2812
rect 30765 2778 30799 2812
rect 30799 2778 30808 2812
rect 30756 2761 30808 2778
rect 30756 2740 30808 2749
rect 30756 2706 30765 2740
rect 30765 2706 30799 2740
rect 30799 2706 30808 2740
rect 30756 2697 30808 2706
rect 30756 2668 30808 2685
rect 30756 2634 30765 2668
rect 30765 2634 30799 2668
rect 30799 2634 30808 2668
rect 30756 2633 30808 2634
rect 30756 2596 30808 2621
rect 30756 2569 30765 2596
rect 30765 2569 30799 2596
rect 30799 2569 30808 2596
rect 30756 2524 30808 2557
rect 30756 2505 30765 2524
rect 30765 2505 30799 2524
rect 30799 2505 30808 2524
rect 30756 2490 30765 2493
rect 30765 2490 30799 2493
rect 30799 2490 30808 2493
rect 30756 2452 30808 2490
rect 30756 2441 30765 2452
rect 30765 2441 30799 2452
rect 30799 2441 30808 2452
rect 30756 2418 30765 2429
rect 30765 2418 30799 2429
rect 30799 2418 30808 2429
rect 30756 2380 30808 2418
rect 30756 2377 30765 2380
rect 30765 2377 30799 2380
rect 30799 2377 30808 2380
rect 30756 2346 30765 2365
rect 30765 2346 30799 2365
rect 30799 2346 30808 2365
rect 30756 2313 30808 2346
rect 30756 2274 30765 2301
rect 30765 2274 30799 2301
rect 30799 2274 30808 2301
rect 30756 2249 30808 2274
rect 30756 2236 30808 2237
rect 30756 2202 30765 2236
rect 30765 2202 30799 2236
rect 30799 2202 30808 2236
rect 30756 2185 30808 2202
rect 30756 2164 30808 2173
rect 30756 2130 30765 2164
rect 30765 2130 30799 2164
rect 30799 2130 30808 2164
rect 30756 2121 30808 2130
rect 30756 2092 30808 2109
rect 30756 2058 30765 2092
rect 30765 2058 30799 2092
rect 30799 2058 30808 2092
rect 30756 2057 30808 2058
rect 30756 2020 30808 2045
rect 30756 1993 30765 2020
rect 30765 1993 30799 2020
rect 30799 1993 30808 2020
rect 30756 1948 30808 1981
rect 30756 1929 30765 1948
rect 30765 1929 30799 1948
rect 30799 1929 30808 1948
rect 30756 1914 30765 1917
rect 30765 1914 30799 1917
rect 30799 1914 30808 1917
rect 30756 1876 30808 1914
rect 30756 1865 30765 1876
rect 30765 1865 30799 1876
rect 30799 1865 30808 1876
rect 30756 1842 30765 1853
rect 30765 1842 30799 1853
rect 30799 1842 30808 1853
rect 30756 1804 30808 1842
rect 30756 1801 30765 1804
rect 30765 1801 30799 1804
rect 30799 1801 30808 1804
rect 30756 1770 30765 1789
rect 30765 1770 30799 1789
rect 30799 1770 30808 1789
rect 30756 1737 30808 1770
rect 30756 1698 30765 1725
rect 30765 1698 30799 1725
rect 30799 1698 30808 1725
rect 30756 1673 30808 1698
rect 30756 1660 30808 1661
rect 30756 1626 30765 1660
rect 30765 1626 30799 1660
rect 30799 1626 30808 1660
rect 30756 1609 30808 1626
rect 30756 1588 30808 1597
rect 30756 1554 30765 1588
rect 30765 1554 30799 1588
rect 30799 1554 30808 1588
rect 30756 1545 30808 1554
rect 30756 1516 30808 1533
rect 30756 1482 30765 1516
rect 30765 1482 30799 1516
rect 30799 1482 30808 1516
rect 30756 1481 30808 1482
rect 30756 1444 30808 1469
rect 30756 1417 30765 1444
rect 30765 1417 30799 1444
rect 30799 1417 30808 1444
rect 30756 1372 30808 1405
rect 30756 1353 30765 1372
rect 30765 1353 30799 1372
rect 30799 1353 30808 1372
rect 30756 1338 30765 1341
rect 30765 1338 30799 1341
rect 30799 1338 30808 1341
rect 30756 1300 30808 1338
rect 30756 1289 30765 1300
rect 30765 1289 30799 1300
rect 30799 1289 30808 1300
rect 30756 1266 30765 1277
rect 30765 1266 30799 1277
rect 30799 1266 30808 1277
rect 30756 1228 30808 1266
rect 30756 1225 30765 1228
rect 30765 1225 30799 1228
rect 30799 1225 30808 1228
rect 30756 1194 30765 1213
rect 30765 1194 30799 1213
rect 30799 1194 30808 1213
rect 30756 1161 30808 1194
rect 30852 3100 30904 3133
rect 30852 3081 30861 3100
rect 30861 3081 30895 3100
rect 30895 3081 30904 3100
rect 30852 3066 30861 3069
rect 30861 3066 30895 3069
rect 30895 3066 30904 3069
rect 30852 3028 30904 3066
rect 30852 3017 30861 3028
rect 30861 3017 30895 3028
rect 30895 3017 30904 3028
rect 30852 2994 30861 3005
rect 30861 2994 30895 3005
rect 30895 2994 30904 3005
rect 30852 2956 30904 2994
rect 30852 2953 30861 2956
rect 30861 2953 30895 2956
rect 30895 2953 30904 2956
rect 30852 2922 30861 2941
rect 30861 2922 30895 2941
rect 30895 2922 30904 2941
rect 30852 2889 30904 2922
rect 30852 2850 30861 2877
rect 30861 2850 30895 2877
rect 30895 2850 30904 2877
rect 30852 2825 30904 2850
rect 30852 2812 30904 2813
rect 30852 2778 30861 2812
rect 30861 2778 30895 2812
rect 30895 2778 30904 2812
rect 30852 2761 30904 2778
rect 30852 2740 30904 2749
rect 30852 2706 30861 2740
rect 30861 2706 30895 2740
rect 30895 2706 30904 2740
rect 30852 2697 30904 2706
rect 30852 2668 30904 2685
rect 30852 2634 30861 2668
rect 30861 2634 30895 2668
rect 30895 2634 30904 2668
rect 30852 2633 30904 2634
rect 30852 2596 30904 2621
rect 30852 2569 30861 2596
rect 30861 2569 30895 2596
rect 30895 2569 30904 2596
rect 30852 2524 30904 2557
rect 30852 2505 30861 2524
rect 30861 2505 30895 2524
rect 30895 2505 30904 2524
rect 30852 2490 30861 2493
rect 30861 2490 30895 2493
rect 30895 2490 30904 2493
rect 30852 2452 30904 2490
rect 30852 2441 30861 2452
rect 30861 2441 30895 2452
rect 30895 2441 30904 2452
rect 30852 2418 30861 2429
rect 30861 2418 30895 2429
rect 30895 2418 30904 2429
rect 30852 2380 30904 2418
rect 30852 2377 30861 2380
rect 30861 2377 30895 2380
rect 30895 2377 30904 2380
rect 30852 2346 30861 2365
rect 30861 2346 30895 2365
rect 30895 2346 30904 2365
rect 30852 2313 30904 2346
rect 30852 2274 30861 2301
rect 30861 2274 30895 2301
rect 30895 2274 30904 2301
rect 30852 2249 30904 2274
rect 30852 2236 30904 2237
rect 30852 2202 30861 2236
rect 30861 2202 30895 2236
rect 30895 2202 30904 2236
rect 30852 2185 30904 2202
rect 30852 2164 30904 2173
rect 30852 2130 30861 2164
rect 30861 2130 30895 2164
rect 30895 2130 30904 2164
rect 30852 2121 30904 2130
rect 30852 2092 30904 2109
rect 30852 2058 30861 2092
rect 30861 2058 30895 2092
rect 30895 2058 30904 2092
rect 30852 2057 30904 2058
rect 30852 2020 30904 2045
rect 30852 1993 30861 2020
rect 30861 1993 30895 2020
rect 30895 1993 30904 2020
rect 30852 1948 30904 1981
rect 30852 1929 30861 1948
rect 30861 1929 30895 1948
rect 30895 1929 30904 1948
rect 30852 1914 30861 1917
rect 30861 1914 30895 1917
rect 30895 1914 30904 1917
rect 30852 1876 30904 1914
rect 30852 1865 30861 1876
rect 30861 1865 30895 1876
rect 30895 1865 30904 1876
rect 30852 1842 30861 1853
rect 30861 1842 30895 1853
rect 30895 1842 30904 1853
rect 30852 1804 30904 1842
rect 30852 1801 30861 1804
rect 30861 1801 30895 1804
rect 30895 1801 30904 1804
rect 30852 1770 30861 1789
rect 30861 1770 30895 1789
rect 30895 1770 30904 1789
rect 30852 1737 30904 1770
rect 30852 1698 30861 1725
rect 30861 1698 30895 1725
rect 30895 1698 30904 1725
rect 30852 1673 30904 1698
rect 30852 1660 30904 1661
rect 30852 1626 30861 1660
rect 30861 1626 30895 1660
rect 30895 1626 30904 1660
rect 30852 1609 30904 1626
rect 30852 1588 30904 1597
rect 30852 1554 30861 1588
rect 30861 1554 30895 1588
rect 30895 1554 30904 1588
rect 30852 1545 30904 1554
rect 30852 1516 30904 1533
rect 30852 1482 30861 1516
rect 30861 1482 30895 1516
rect 30895 1482 30904 1516
rect 30852 1481 30904 1482
rect 30852 1444 30904 1469
rect 30852 1417 30861 1444
rect 30861 1417 30895 1444
rect 30895 1417 30904 1444
rect 30852 1372 30904 1405
rect 30852 1353 30861 1372
rect 30861 1353 30895 1372
rect 30895 1353 30904 1372
rect 30852 1338 30861 1341
rect 30861 1338 30895 1341
rect 30895 1338 30904 1341
rect 30852 1300 30904 1338
rect 30852 1289 30861 1300
rect 30861 1289 30895 1300
rect 30895 1289 30904 1300
rect 30852 1266 30861 1277
rect 30861 1266 30895 1277
rect 30895 1266 30904 1277
rect 30852 1228 30904 1266
rect 30852 1225 30861 1228
rect 30861 1225 30895 1228
rect 30895 1225 30904 1228
rect 30852 1194 30861 1213
rect 30861 1194 30895 1213
rect 30895 1194 30904 1213
rect 30852 1161 30904 1194
rect 30948 3100 31000 3133
rect 30948 3081 30957 3100
rect 30957 3081 30991 3100
rect 30991 3081 31000 3100
rect 30948 3066 30957 3069
rect 30957 3066 30991 3069
rect 30991 3066 31000 3069
rect 30948 3028 31000 3066
rect 30948 3017 30957 3028
rect 30957 3017 30991 3028
rect 30991 3017 31000 3028
rect 30948 2994 30957 3005
rect 30957 2994 30991 3005
rect 30991 2994 31000 3005
rect 30948 2956 31000 2994
rect 30948 2953 30957 2956
rect 30957 2953 30991 2956
rect 30991 2953 31000 2956
rect 30948 2922 30957 2941
rect 30957 2922 30991 2941
rect 30991 2922 31000 2941
rect 30948 2889 31000 2922
rect 30948 2850 30957 2877
rect 30957 2850 30991 2877
rect 30991 2850 31000 2877
rect 30948 2825 31000 2850
rect 30948 2812 31000 2813
rect 30948 2778 30957 2812
rect 30957 2778 30991 2812
rect 30991 2778 31000 2812
rect 30948 2761 31000 2778
rect 30948 2740 31000 2749
rect 30948 2706 30957 2740
rect 30957 2706 30991 2740
rect 30991 2706 31000 2740
rect 30948 2697 31000 2706
rect 30948 2668 31000 2685
rect 30948 2634 30957 2668
rect 30957 2634 30991 2668
rect 30991 2634 31000 2668
rect 30948 2633 31000 2634
rect 30948 2596 31000 2621
rect 30948 2569 30957 2596
rect 30957 2569 30991 2596
rect 30991 2569 31000 2596
rect 30948 2524 31000 2557
rect 30948 2505 30957 2524
rect 30957 2505 30991 2524
rect 30991 2505 31000 2524
rect 30948 2490 30957 2493
rect 30957 2490 30991 2493
rect 30991 2490 31000 2493
rect 30948 2452 31000 2490
rect 30948 2441 30957 2452
rect 30957 2441 30991 2452
rect 30991 2441 31000 2452
rect 30948 2418 30957 2429
rect 30957 2418 30991 2429
rect 30991 2418 31000 2429
rect 30948 2380 31000 2418
rect 30948 2377 30957 2380
rect 30957 2377 30991 2380
rect 30991 2377 31000 2380
rect 30948 2346 30957 2365
rect 30957 2346 30991 2365
rect 30991 2346 31000 2365
rect 30948 2313 31000 2346
rect 30948 2274 30957 2301
rect 30957 2274 30991 2301
rect 30991 2274 31000 2301
rect 30948 2249 31000 2274
rect 30948 2236 31000 2237
rect 30948 2202 30957 2236
rect 30957 2202 30991 2236
rect 30991 2202 31000 2236
rect 30948 2185 31000 2202
rect 30948 2164 31000 2173
rect 30948 2130 30957 2164
rect 30957 2130 30991 2164
rect 30991 2130 31000 2164
rect 30948 2121 31000 2130
rect 30948 2092 31000 2109
rect 30948 2058 30957 2092
rect 30957 2058 30991 2092
rect 30991 2058 31000 2092
rect 30948 2057 31000 2058
rect 30948 2020 31000 2045
rect 30948 1993 30957 2020
rect 30957 1993 30991 2020
rect 30991 1993 31000 2020
rect 30948 1948 31000 1981
rect 30948 1929 30957 1948
rect 30957 1929 30991 1948
rect 30991 1929 31000 1948
rect 30948 1914 30957 1917
rect 30957 1914 30991 1917
rect 30991 1914 31000 1917
rect 30948 1876 31000 1914
rect 30948 1865 30957 1876
rect 30957 1865 30991 1876
rect 30991 1865 31000 1876
rect 30948 1842 30957 1853
rect 30957 1842 30991 1853
rect 30991 1842 31000 1853
rect 30948 1804 31000 1842
rect 30948 1801 30957 1804
rect 30957 1801 30991 1804
rect 30991 1801 31000 1804
rect 30948 1770 30957 1789
rect 30957 1770 30991 1789
rect 30991 1770 31000 1789
rect 30948 1737 31000 1770
rect 30948 1698 30957 1725
rect 30957 1698 30991 1725
rect 30991 1698 31000 1725
rect 30948 1673 31000 1698
rect 30948 1660 31000 1661
rect 30948 1626 30957 1660
rect 30957 1626 30991 1660
rect 30991 1626 31000 1660
rect 30948 1609 31000 1626
rect 30948 1588 31000 1597
rect 30948 1554 30957 1588
rect 30957 1554 30991 1588
rect 30991 1554 31000 1588
rect 30948 1545 31000 1554
rect 30948 1516 31000 1533
rect 30948 1482 30957 1516
rect 30957 1482 30991 1516
rect 30991 1482 31000 1516
rect 30948 1481 31000 1482
rect 30948 1444 31000 1469
rect 30948 1417 30957 1444
rect 30957 1417 30991 1444
rect 30991 1417 31000 1444
rect 30948 1372 31000 1405
rect 30948 1353 30957 1372
rect 30957 1353 30991 1372
rect 30991 1353 31000 1372
rect 30948 1338 30957 1341
rect 30957 1338 30991 1341
rect 30991 1338 31000 1341
rect 30948 1300 31000 1338
rect 30948 1289 30957 1300
rect 30957 1289 30991 1300
rect 30991 1289 31000 1300
rect 30948 1266 30957 1277
rect 30957 1266 30991 1277
rect 30991 1266 31000 1277
rect 30948 1228 31000 1266
rect 30948 1225 30957 1228
rect 30957 1225 30991 1228
rect 30991 1225 31000 1228
rect 30948 1194 30957 1213
rect 30957 1194 30991 1213
rect 30991 1194 31000 1213
rect 30948 1161 31000 1194
rect 31044 3100 31096 3133
rect 31044 3081 31053 3100
rect 31053 3081 31087 3100
rect 31087 3081 31096 3100
rect 31044 3066 31053 3069
rect 31053 3066 31087 3069
rect 31087 3066 31096 3069
rect 31044 3028 31096 3066
rect 31044 3017 31053 3028
rect 31053 3017 31087 3028
rect 31087 3017 31096 3028
rect 31044 2994 31053 3005
rect 31053 2994 31087 3005
rect 31087 2994 31096 3005
rect 31044 2956 31096 2994
rect 31044 2953 31053 2956
rect 31053 2953 31087 2956
rect 31087 2953 31096 2956
rect 31044 2922 31053 2941
rect 31053 2922 31087 2941
rect 31087 2922 31096 2941
rect 31044 2889 31096 2922
rect 31044 2850 31053 2877
rect 31053 2850 31087 2877
rect 31087 2850 31096 2877
rect 31044 2825 31096 2850
rect 31044 2812 31096 2813
rect 31044 2778 31053 2812
rect 31053 2778 31087 2812
rect 31087 2778 31096 2812
rect 31044 2761 31096 2778
rect 31044 2740 31096 2749
rect 31044 2706 31053 2740
rect 31053 2706 31087 2740
rect 31087 2706 31096 2740
rect 31044 2697 31096 2706
rect 31044 2668 31096 2685
rect 31044 2634 31053 2668
rect 31053 2634 31087 2668
rect 31087 2634 31096 2668
rect 31044 2633 31096 2634
rect 31044 2596 31096 2621
rect 31044 2569 31053 2596
rect 31053 2569 31087 2596
rect 31087 2569 31096 2596
rect 31044 2524 31096 2557
rect 31044 2505 31053 2524
rect 31053 2505 31087 2524
rect 31087 2505 31096 2524
rect 31044 2490 31053 2493
rect 31053 2490 31087 2493
rect 31087 2490 31096 2493
rect 31044 2452 31096 2490
rect 31044 2441 31053 2452
rect 31053 2441 31087 2452
rect 31087 2441 31096 2452
rect 31044 2418 31053 2429
rect 31053 2418 31087 2429
rect 31087 2418 31096 2429
rect 31044 2380 31096 2418
rect 31044 2377 31053 2380
rect 31053 2377 31087 2380
rect 31087 2377 31096 2380
rect 31044 2346 31053 2365
rect 31053 2346 31087 2365
rect 31087 2346 31096 2365
rect 31044 2313 31096 2346
rect 31044 2274 31053 2301
rect 31053 2274 31087 2301
rect 31087 2274 31096 2301
rect 31044 2249 31096 2274
rect 31044 2236 31096 2237
rect 31044 2202 31053 2236
rect 31053 2202 31087 2236
rect 31087 2202 31096 2236
rect 31044 2185 31096 2202
rect 31044 2164 31096 2173
rect 31044 2130 31053 2164
rect 31053 2130 31087 2164
rect 31087 2130 31096 2164
rect 31044 2121 31096 2130
rect 31044 2092 31096 2109
rect 31044 2058 31053 2092
rect 31053 2058 31087 2092
rect 31087 2058 31096 2092
rect 31044 2057 31096 2058
rect 31044 2020 31096 2045
rect 31044 1993 31053 2020
rect 31053 1993 31087 2020
rect 31087 1993 31096 2020
rect 31044 1948 31096 1981
rect 31044 1929 31053 1948
rect 31053 1929 31087 1948
rect 31087 1929 31096 1948
rect 31044 1914 31053 1917
rect 31053 1914 31087 1917
rect 31087 1914 31096 1917
rect 31044 1876 31096 1914
rect 31044 1865 31053 1876
rect 31053 1865 31087 1876
rect 31087 1865 31096 1876
rect 31044 1842 31053 1853
rect 31053 1842 31087 1853
rect 31087 1842 31096 1853
rect 31044 1804 31096 1842
rect 31044 1801 31053 1804
rect 31053 1801 31087 1804
rect 31087 1801 31096 1804
rect 31044 1770 31053 1789
rect 31053 1770 31087 1789
rect 31087 1770 31096 1789
rect 31044 1737 31096 1770
rect 31044 1698 31053 1725
rect 31053 1698 31087 1725
rect 31087 1698 31096 1725
rect 31044 1673 31096 1698
rect 31044 1660 31096 1661
rect 31044 1626 31053 1660
rect 31053 1626 31087 1660
rect 31087 1626 31096 1660
rect 31044 1609 31096 1626
rect 31044 1588 31096 1597
rect 31044 1554 31053 1588
rect 31053 1554 31087 1588
rect 31087 1554 31096 1588
rect 31044 1545 31096 1554
rect 31044 1516 31096 1533
rect 31044 1482 31053 1516
rect 31053 1482 31087 1516
rect 31087 1482 31096 1516
rect 31044 1481 31096 1482
rect 31044 1444 31096 1469
rect 31044 1417 31053 1444
rect 31053 1417 31087 1444
rect 31087 1417 31096 1444
rect 31044 1372 31096 1405
rect 31044 1353 31053 1372
rect 31053 1353 31087 1372
rect 31087 1353 31096 1372
rect 31044 1338 31053 1341
rect 31053 1338 31087 1341
rect 31087 1338 31096 1341
rect 31044 1300 31096 1338
rect 31044 1289 31053 1300
rect 31053 1289 31087 1300
rect 31087 1289 31096 1300
rect 31044 1266 31053 1277
rect 31053 1266 31087 1277
rect 31087 1266 31096 1277
rect 31044 1228 31096 1266
rect 31044 1225 31053 1228
rect 31053 1225 31087 1228
rect 31087 1225 31096 1228
rect 31044 1194 31053 1213
rect 31053 1194 31087 1213
rect 31087 1194 31096 1213
rect 31044 1161 31096 1194
rect 31140 3100 31192 3133
rect 31140 3081 31149 3100
rect 31149 3081 31183 3100
rect 31183 3081 31192 3100
rect 31140 3066 31149 3069
rect 31149 3066 31183 3069
rect 31183 3066 31192 3069
rect 31140 3028 31192 3066
rect 31140 3017 31149 3028
rect 31149 3017 31183 3028
rect 31183 3017 31192 3028
rect 31140 2994 31149 3005
rect 31149 2994 31183 3005
rect 31183 2994 31192 3005
rect 31140 2956 31192 2994
rect 31140 2953 31149 2956
rect 31149 2953 31183 2956
rect 31183 2953 31192 2956
rect 31140 2922 31149 2941
rect 31149 2922 31183 2941
rect 31183 2922 31192 2941
rect 31140 2889 31192 2922
rect 31140 2850 31149 2877
rect 31149 2850 31183 2877
rect 31183 2850 31192 2877
rect 31140 2825 31192 2850
rect 31140 2812 31192 2813
rect 31140 2778 31149 2812
rect 31149 2778 31183 2812
rect 31183 2778 31192 2812
rect 31140 2761 31192 2778
rect 31140 2740 31192 2749
rect 31140 2706 31149 2740
rect 31149 2706 31183 2740
rect 31183 2706 31192 2740
rect 31140 2697 31192 2706
rect 31140 2668 31192 2685
rect 31140 2634 31149 2668
rect 31149 2634 31183 2668
rect 31183 2634 31192 2668
rect 31140 2633 31192 2634
rect 31140 2596 31192 2621
rect 31140 2569 31149 2596
rect 31149 2569 31183 2596
rect 31183 2569 31192 2596
rect 31140 2524 31192 2557
rect 31140 2505 31149 2524
rect 31149 2505 31183 2524
rect 31183 2505 31192 2524
rect 31140 2490 31149 2493
rect 31149 2490 31183 2493
rect 31183 2490 31192 2493
rect 31140 2452 31192 2490
rect 31140 2441 31149 2452
rect 31149 2441 31183 2452
rect 31183 2441 31192 2452
rect 31140 2418 31149 2429
rect 31149 2418 31183 2429
rect 31183 2418 31192 2429
rect 31140 2380 31192 2418
rect 31140 2377 31149 2380
rect 31149 2377 31183 2380
rect 31183 2377 31192 2380
rect 31140 2346 31149 2365
rect 31149 2346 31183 2365
rect 31183 2346 31192 2365
rect 31140 2313 31192 2346
rect 31140 2274 31149 2301
rect 31149 2274 31183 2301
rect 31183 2274 31192 2301
rect 31140 2249 31192 2274
rect 31140 2236 31192 2237
rect 31140 2202 31149 2236
rect 31149 2202 31183 2236
rect 31183 2202 31192 2236
rect 31140 2185 31192 2202
rect 31140 2164 31192 2173
rect 31140 2130 31149 2164
rect 31149 2130 31183 2164
rect 31183 2130 31192 2164
rect 31140 2121 31192 2130
rect 31140 2092 31192 2109
rect 31140 2058 31149 2092
rect 31149 2058 31183 2092
rect 31183 2058 31192 2092
rect 31140 2057 31192 2058
rect 31140 2020 31192 2045
rect 31140 1993 31149 2020
rect 31149 1993 31183 2020
rect 31183 1993 31192 2020
rect 31140 1948 31192 1981
rect 31140 1929 31149 1948
rect 31149 1929 31183 1948
rect 31183 1929 31192 1948
rect 31140 1914 31149 1917
rect 31149 1914 31183 1917
rect 31183 1914 31192 1917
rect 31140 1876 31192 1914
rect 31140 1865 31149 1876
rect 31149 1865 31183 1876
rect 31183 1865 31192 1876
rect 31140 1842 31149 1853
rect 31149 1842 31183 1853
rect 31183 1842 31192 1853
rect 31140 1804 31192 1842
rect 31140 1801 31149 1804
rect 31149 1801 31183 1804
rect 31183 1801 31192 1804
rect 31140 1770 31149 1789
rect 31149 1770 31183 1789
rect 31183 1770 31192 1789
rect 31140 1737 31192 1770
rect 31140 1698 31149 1725
rect 31149 1698 31183 1725
rect 31183 1698 31192 1725
rect 31140 1673 31192 1698
rect 31140 1660 31192 1661
rect 31140 1626 31149 1660
rect 31149 1626 31183 1660
rect 31183 1626 31192 1660
rect 31140 1609 31192 1626
rect 31140 1588 31192 1597
rect 31140 1554 31149 1588
rect 31149 1554 31183 1588
rect 31183 1554 31192 1588
rect 31140 1545 31192 1554
rect 31140 1516 31192 1533
rect 31140 1482 31149 1516
rect 31149 1482 31183 1516
rect 31183 1482 31192 1516
rect 31140 1481 31192 1482
rect 31140 1444 31192 1469
rect 31140 1417 31149 1444
rect 31149 1417 31183 1444
rect 31183 1417 31192 1444
rect 31140 1372 31192 1405
rect 31140 1353 31149 1372
rect 31149 1353 31183 1372
rect 31183 1353 31192 1372
rect 31140 1338 31149 1341
rect 31149 1338 31183 1341
rect 31183 1338 31192 1341
rect 31140 1300 31192 1338
rect 31140 1289 31149 1300
rect 31149 1289 31183 1300
rect 31183 1289 31192 1300
rect 31140 1266 31149 1277
rect 31149 1266 31183 1277
rect 31183 1266 31192 1277
rect 31140 1228 31192 1266
rect 31140 1225 31149 1228
rect 31149 1225 31183 1228
rect 31183 1225 31192 1228
rect 31140 1194 31149 1213
rect 31149 1194 31183 1213
rect 31183 1194 31192 1213
rect 31140 1161 31192 1194
rect 31236 3100 31288 3133
rect 31236 3081 31245 3100
rect 31245 3081 31279 3100
rect 31279 3081 31288 3100
rect 31236 3066 31245 3069
rect 31245 3066 31279 3069
rect 31279 3066 31288 3069
rect 31236 3028 31288 3066
rect 31236 3017 31245 3028
rect 31245 3017 31279 3028
rect 31279 3017 31288 3028
rect 31236 2994 31245 3005
rect 31245 2994 31279 3005
rect 31279 2994 31288 3005
rect 31236 2956 31288 2994
rect 31236 2953 31245 2956
rect 31245 2953 31279 2956
rect 31279 2953 31288 2956
rect 31236 2922 31245 2941
rect 31245 2922 31279 2941
rect 31279 2922 31288 2941
rect 31236 2889 31288 2922
rect 31236 2850 31245 2877
rect 31245 2850 31279 2877
rect 31279 2850 31288 2877
rect 31236 2825 31288 2850
rect 31236 2812 31288 2813
rect 31236 2778 31245 2812
rect 31245 2778 31279 2812
rect 31279 2778 31288 2812
rect 31236 2761 31288 2778
rect 31236 2740 31288 2749
rect 31236 2706 31245 2740
rect 31245 2706 31279 2740
rect 31279 2706 31288 2740
rect 31236 2697 31288 2706
rect 31236 2668 31288 2685
rect 31236 2634 31245 2668
rect 31245 2634 31279 2668
rect 31279 2634 31288 2668
rect 31236 2633 31288 2634
rect 31236 2596 31288 2621
rect 31236 2569 31245 2596
rect 31245 2569 31279 2596
rect 31279 2569 31288 2596
rect 31236 2524 31288 2557
rect 31236 2505 31245 2524
rect 31245 2505 31279 2524
rect 31279 2505 31288 2524
rect 31236 2490 31245 2493
rect 31245 2490 31279 2493
rect 31279 2490 31288 2493
rect 31236 2452 31288 2490
rect 31236 2441 31245 2452
rect 31245 2441 31279 2452
rect 31279 2441 31288 2452
rect 31236 2418 31245 2429
rect 31245 2418 31279 2429
rect 31279 2418 31288 2429
rect 31236 2380 31288 2418
rect 31236 2377 31245 2380
rect 31245 2377 31279 2380
rect 31279 2377 31288 2380
rect 31236 2346 31245 2365
rect 31245 2346 31279 2365
rect 31279 2346 31288 2365
rect 31236 2313 31288 2346
rect 31236 2274 31245 2301
rect 31245 2274 31279 2301
rect 31279 2274 31288 2301
rect 31236 2249 31288 2274
rect 31236 2236 31288 2237
rect 31236 2202 31245 2236
rect 31245 2202 31279 2236
rect 31279 2202 31288 2236
rect 31236 2185 31288 2202
rect 31236 2164 31288 2173
rect 31236 2130 31245 2164
rect 31245 2130 31279 2164
rect 31279 2130 31288 2164
rect 31236 2121 31288 2130
rect 31236 2092 31288 2109
rect 31236 2058 31245 2092
rect 31245 2058 31279 2092
rect 31279 2058 31288 2092
rect 31236 2057 31288 2058
rect 31236 2020 31288 2045
rect 31236 1993 31245 2020
rect 31245 1993 31279 2020
rect 31279 1993 31288 2020
rect 31236 1948 31288 1981
rect 31236 1929 31245 1948
rect 31245 1929 31279 1948
rect 31279 1929 31288 1948
rect 31236 1914 31245 1917
rect 31245 1914 31279 1917
rect 31279 1914 31288 1917
rect 31236 1876 31288 1914
rect 31236 1865 31245 1876
rect 31245 1865 31279 1876
rect 31279 1865 31288 1876
rect 31236 1842 31245 1853
rect 31245 1842 31279 1853
rect 31279 1842 31288 1853
rect 31236 1804 31288 1842
rect 31236 1801 31245 1804
rect 31245 1801 31279 1804
rect 31279 1801 31288 1804
rect 31236 1770 31245 1789
rect 31245 1770 31279 1789
rect 31279 1770 31288 1789
rect 31236 1737 31288 1770
rect 31236 1698 31245 1725
rect 31245 1698 31279 1725
rect 31279 1698 31288 1725
rect 31236 1673 31288 1698
rect 31236 1660 31288 1661
rect 31236 1626 31245 1660
rect 31245 1626 31279 1660
rect 31279 1626 31288 1660
rect 31236 1609 31288 1626
rect 31236 1588 31288 1597
rect 31236 1554 31245 1588
rect 31245 1554 31279 1588
rect 31279 1554 31288 1588
rect 31236 1545 31288 1554
rect 31236 1516 31288 1533
rect 31236 1482 31245 1516
rect 31245 1482 31279 1516
rect 31279 1482 31288 1516
rect 31236 1481 31288 1482
rect 31236 1444 31288 1469
rect 31236 1417 31245 1444
rect 31245 1417 31279 1444
rect 31279 1417 31288 1444
rect 31236 1372 31288 1405
rect 31236 1353 31245 1372
rect 31245 1353 31279 1372
rect 31279 1353 31288 1372
rect 31236 1338 31245 1341
rect 31245 1338 31279 1341
rect 31279 1338 31288 1341
rect 31236 1300 31288 1338
rect 31236 1289 31245 1300
rect 31245 1289 31279 1300
rect 31279 1289 31288 1300
rect 31236 1266 31245 1277
rect 31245 1266 31279 1277
rect 31279 1266 31288 1277
rect 31236 1228 31288 1266
rect 31236 1225 31245 1228
rect 31245 1225 31279 1228
rect 31279 1225 31288 1228
rect 31236 1194 31245 1213
rect 31245 1194 31279 1213
rect 31279 1194 31288 1213
rect 31236 1161 31288 1194
rect 31332 3100 31384 3133
rect 31332 3081 31341 3100
rect 31341 3081 31375 3100
rect 31375 3081 31384 3100
rect 31332 3066 31341 3069
rect 31341 3066 31375 3069
rect 31375 3066 31384 3069
rect 31332 3028 31384 3066
rect 31332 3017 31341 3028
rect 31341 3017 31375 3028
rect 31375 3017 31384 3028
rect 31332 2994 31341 3005
rect 31341 2994 31375 3005
rect 31375 2994 31384 3005
rect 31332 2956 31384 2994
rect 31332 2953 31341 2956
rect 31341 2953 31375 2956
rect 31375 2953 31384 2956
rect 31332 2922 31341 2941
rect 31341 2922 31375 2941
rect 31375 2922 31384 2941
rect 31332 2889 31384 2922
rect 31332 2850 31341 2877
rect 31341 2850 31375 2877
rect 31375 2850 31384 2877
rect 31332 2825 31384 2850
rect 31332 2812 31384 2813
rect 31332 2778 31341 2812
rect 31341 2778 31375 2812
rect 31375 2778 31384 2812
rect 31332 2761 31384 2778
rect 31332 2740 31384 2749
rect 31332 2706 31341 2740
rect 31341 2706 31375 2740
rect 31375 2706 31384 2740
rect 31332 2697 31384 2706
rect 31332 2668 31384 2685
rect 31332 2634 31341 2668
rect 31341 2634 31375 2668
rect 31375 2634 31384 2668
rect 31332 2633 31384 2634
rect 31332 2596 31384 2621
rect 31332 2569 31341 2596
rect 31341 2569 31375 2596
rect 31375 2569 31384 2596
rect 31332 2524 31384 2557
rect 31332 2505 31341 2524
rect 31341 2505 31375 2524
rect 31375 2505 31384 2524
rect 31332 2490 31341 2493
rect 31341 2490 31375 2493
rect 31375 2490 31384 2493
rect 31332 2452 31384 2490
rect 31332 2441 31341 2452
rect 31341 2441 31375 2452
rect 31375 2441 31384 2452
rect 31332 2418 31341 2429
rect 31341 2418 31375 2429
rect 31375 2418 31384 2429
rect 31332 2380 31384 2418
rect 31332 2377 31341 2380
rect 31341 2377 31375 2380
rect 31375 2377 31384 2380
rect 31332 2346 31341 2365
rect 31341 2346 31375 2365
rect 31375 2346 31384 2365
rect 31332 2313 31384 2346
rect 31332 2274 31341 2301
rect 31341 2274 31375 2301
rect 31375 2274 31384 2301
rect 31332 2249 31384 2274
rect 31332 2236 31384 2237
rect 31332 2202 31341 2236
rect 31341 2202 31375 2236
rect 31375 2202 31384 2236
rect 31332 2185 31384 2202
rect 31332 2164 31384 2173
rect 31332 2130 31341 2164
rect 31341 2130 31375 2164
rect 31375 2130 31384 2164
rect 31332 2121 31384 2130
rect 31332 2092 31384 2109
rect 31332 2058 31341 2092
rect 31341 2058 31375 2092
rect 31375 2058 31384 2092
rect 31332 2057 31384 2058
rect 31332 2020 31384 2045
rect 31332 1993 31341 2020
rect 31341 1993 31375 2020
rect 31375 1993 31384 2020
rect 31332 1948 31384 1981
rect 31332 1929 31341 1948
rect 31341 1929 31375 1948
rect 31375 1929 31384 1948
rect 31332 1914 31341 1917
rect 31341 1914 31375 1917
rect 31375 1914 31384 1917
rect 31332 1876 31384 1914
rect 31332 1865 31341 1876
rect 31341 1865 31375 1876
rect 31375 1865 31384 1876
rect 31332 1842 31341 1853
rect 31341 1842 31375 1853
rect 31375 1842 31384 1853
rect 31332 1804 31384 1842
rect 31332 1801 31341 1804
rect 31341 1801 31375 1804
rect 31375 1801 31384 1804
rect 31332 1770 31341 1789
rect 31341 1770 31375 1789
rect 31375 1770 31384 1789
rect 31332 1737 31384 1770
rect 31332 1698 31341 1725
rect 31341 1698 31375 1725
rect 31375 1698 31384 1725
rect 31332 1673 31384 1698
rect 31332 1660 31384 1661
rect 31332 1626 31341 1660
rect 31341 1626 31375 1660
rect 31375 1626 31384 1660
rect 31332 1609 31384 1626
rect 31332 1588 31384 1597
rect 31332 1554 31341 1588
rect 31341 1554 31375 1588
rect 31375 1554 31384 1588
rect 31332 1545 31384 1554
rect 31332 1516 31384 1533
rect 31332 1482 31341 1516
rect 31341 1482 31375 1516
rect 31375 1482 31384 1516
rect 31332 1481 31384 1482
rect 31332 1444 31384 1469
rect 31332 1417 31341 1444
rect 31341 1417 31375 1444
rect 31375 1417 31384 1444
rect 31332 1372 31384 1405
rect 31332 1353 31341 1372
rect 31341 1353 31375 1372
rect 31375 1353 31384 1372
rect 31332 1338 31341 1341
rect 31341 1338 31375 1341
rect 31375 1338 31384 1341
rect 31332 1300 31384 1338
rect 31332 1289 31341 1300
rect 31341 1289 31375 1300
rect 31375 1289 31384 1300
rect 31332 1266 31341 1277
rect 31341 1266 31375 1277
rect 31375 1266 31384 1277
rect 31332 1228 31384 1266
rect 31332 1225 31341 1228
rect 31341 1225 31375 1228
rect 31375 1225 31384 1228
rect 31332 1194 31341 1213
rect 31341 1194 31375 1213
rect 31375 1194 31384 1213
rect 31332 1161 31384 1194
rect 31428 3100 31480 3133
rect 31428 3081 31437 3100
rect 31437 3081 31471 3100
rect 31471 3081 31480 3100
rect 31428 3066 31437 3069
rect 31437 3066 31471 3069
rect 31471 3066 31480 3069
rect 31428 3028 31480 3066
rect 31428 3017 31437 3028
rect 31437 3017 31471 3028
rect 31471 3017 31480 3028
rect 31428 2994 31437 3005
rect 31437 2994 31471 3005
rect 31471 2994 31480 3005
rect 31428 2956 31480 2994
rect 31428 2953 31437 2956
rect 31437 2953 31471 2956
rect 31471 2953 31480 2956
rect 31428 2922 31437 2941
rect 31437 2922 31471 2941
rect 31471 2922 31480 2941
rect 31428 2889 31480 2922
rect 31428 2850 31437 2877
rect 31437 2850 31471 2877
rect 31471 2850 31480 2877
rect 31428 2825 31480 2850
rect 31428 2812 31480 2813
rect 31428 2778 31437 2812
rect 31437 2778 31471 2812
rect 31471 2778 31480 2812
rect 31428 2761 31480 2778
rect 31428 2740 31480 2749
rect 31428 2706 31437 2740
rect 31437 2706 31471 2740
rect 31471 2706 31480 2740
rect 31428 2697 31480 2706
rect 31428 2668 31480 2685
rect 31428 2634 31437 2668
rect 31437 2634 31471 2668
rect 31471 2634 31480 2668
rect 31428 2633 31480 2634
rect 31428 2596 31480 2621
rect 31428 2569 31437 2596
rect 31437 2569 31471 2596
rect 31471 2569 31480 2596
rect 31428 2524 31480 2557
rect 31428 2505 31437 2524
rect 31437 2505 31471 2524
rect 31471 2505 31480 2524
rect 31428 2490 31437 2493
rect 31437 2490 31471 2493
rect 31471 2490 31480 2493
rect 31428 2452 31480 2490
rect 31428 2441 31437 2452
rect 31437 2441 31471 2452
rect 31471 2441 31480 2452
rect 31428 2418 31437 2429
rect 31437 2418 31471 2429
rect 31471 2418 31480 2429
rect 31428 2380 31480 2418
rect 31428 2377 31437 2380
rect 31437 2377 31471 2380
rect 31471 2377 31480 2380
rect 31428 2346 31437 2365
rect 31437 2346 31471 2365
rect 31471 2346 31480 2365
rect 31428 2313 31480 2346
rect 31428 2274 31437 2301
rect 31437 2274 31471 2301
rect 31471 2274 31480 2301
rect 31428 2249 31480 2274
rect 31428 2236 31480 2237
rect 31428 2202 31437 2236
rect 31437 2202 31471 2236
rect 31471 2202 31480 2236
rect 31428 2185 31480 2202
rect 31428 2164 31480 2173
rect 31428 2130 31437 2164
rect 31437 2130 31471 2164
rect 31471 2130 31480 2164
rect 31428 2121 31480 2130
rect 31428 2092 31480 2109
rect 31428 2058 31437 2092
rect 31437 2058 31471 2092
rect 31471 2058 31480 2092
rect 31428 2057 31480 2058
rect 31428 2020 31480 2045
rect 31428 1993 31437 2020
rect 31437 1993 31471 2020
rect 31471 1993 31480 2020
rect 31428 1948 31480 1981
rect 31428 1929 31437 1948
rect 31437 1929 31471 1948
rect 31471 1929 31480 1948
rect 31428 1914 31437 1917
rect 31437 1914 31471 1917
rect 31471 1914 31480 1917
rect 31428 1876 31480 1914
rect 31428 1865 31437 1876
rect 31437 1865 31471 1876
rect 31471 1865 31480 1876
rect 31428 1842 31437 1853
rect 31437 1842 31471 1853
rect 31471 1842 31480 1853
rect 31428 1804 31480 1842
rect 31428 1801 31437 1804
rect 31437 1801 31471 1804
rect 31471 1801 31480 1804
rect 31428 1770 31437 1789
rect 31437 1770 31471 1789
rect 31471 1770 31480 1789
rect 31428 1737 31480 1770
rect 31428 1698 31437 1725
rect 31437 1698 31471 1725
rect 31471 1698 31480 1725
rect 31428 1673 31480 1698
rect 31428 1660 31480 1661
rect 31428 1626 31437 1660
rect 31437 1626 31471 1660
rect 31471 1626 31480 1660
rect 31428 1609 31480 1626
rect 31428 1588 31480 1597
rect 31428 1554 31437 1588
rect 31437 1554 31471 1588
rect 31471 1554 31480 1588
rect 31428 1545 31480 1554
rect 31428 1516 31480 1533
rect 31428 1482 31437 1516
rect 31437 1482 31471 1516
rect 31471 1482 31480 1516
rect 31428 1481 31480 1482
rect 31428 1444 31480 1469
rect 31428 1417 31437 1444
rect 31437 1417 31471 1444
rect 31471 1417 31480 1444
rect 31428 1372 31480 1405
rect 31428 1353 31437 1372
rect 31437 1353 31471 1372
rect 31471 1353 31480 1372
rect 31428 1338 31437 1341
rect 31437 1338 31471 1341
rect 31471 1338 31480 1341
rect 31428 1300 31480 1338
rect 31428 1289 31437 1300
rect 31437 1289 31471 1300
rect 31471 1289 31480 1300
rect 31428 1266 31437 1277
rect 31437 1266 31471 1277
rect 31471 1266 31480 1277
rect 31428 1228 31480 1266
rect 31428 1225 31437 1228
rect 31437 1225 31471 1228
rect 31471 1225 31480 1228
rect 31428 1194 31437 1213
rect 31437 1194 31471 1213
rect 31471 1194 31480 1213
rect 31428 1161 31480 1194
rect 31524 3100 31576 3133
rect 31524 3081 31533 3100
rect 31533 3081 31567 3100
rect 31567 3081 31576 3100
rect 31524 3066 31533 3069
rect 31533 3066 31567 3069
rect 31567 3066 31576 3069
rect 31524 3028 31576 3066
rect 31524 3017 31533 3028
rect 31533 3017 31567 3028
rect 31567 3017 31576 3028
rect 31524 2994 31533 3005
rect 31533 2994 31567 3005
rect 31567 2994 31576 3005
rect 31524 2956 31576 2994
rect 31524 2953 31533 2956
rect 31533 2953 31567 2956
rect 31567 2953 31576 2956
rect 31524 2922 31533 2941
rect 31533 2922 31567 2941
rect 31567 2922 31576 2941
rect 31524 2889 31576 2922
rect 31524 2850 31533 2877
rect 31533 2850 31567 2877
rect 31567 2850 31576 2877
rect 31524 2825 31576 2850
rect 31524 2812 31576 2813
rect 31524 2778 31533 2812
rect 31533 2778 31567 2812
rect 31567 2778 31576 2812
rect 31524 2761 31576 2778
rect 31524 2740 31576 2749
rect 31524 2706 31533 2740
rect 31533 2706 31567 2740
rect 31567 2706 31576 2740
rect 31524 2697 31576 2706
rect 31524 2668 31576 2685
rect 31524 2634 31533 2668
rect 31533 2634 31567 2668
rect 31567 2634 31576 2668
rect 31524 2633 31576 2634
rect 31524 2596 31576 2621
rect 31524 2569 31533 2596
rect 31533 2569 31567 2596
rect 31567 2569 31576 2596
rect 31524 2524 31576 2557
rect 31524 2505 31533 2524
rect 31533 2505 31567 2524
rect 31567 2505 31576 2524
rect 31524 2490 31533 2493
rect 31533 2490 31567 2493
rect 31567 2490 31576 2493
rect 31524 2452 31576 2490
rect 31524 2441 31533 2452
rect 31533 2441 31567 2452
rect 31567 2441 31576 2452
rect 31524 2418 31533 2429
rect 31533 2418 31567 2429
rect 31567 2418 31576 2429
rect 31524 2380 31576 2418
rect 31524 2377 31533 2380
rect 31533 2377 31567 2380
rect 31567 2377 31576 2380
rect 31524 2346 31533 2365
rect 31533 2346 31567 2365
rect 31567 2346 31576 2365
rect 31524 2313 31576 2346
rect 31524 2274 31533 2301
rect 31533 2274 31567 2301
rect 31567 2274 31576 2301
rect 31524 2249 31576 2274
rect 31524 2236 31576 2237
rect 31524 2202 31533 2236
rect 31533 2202 31567 2236
rect 31567 2202 31576 2236
rect 31524 2185 31576 2202
rect 31524 2164 31576 2173
rect 31524 2130 31533 2164
rect 31533 2130 31567 2164
rect 31567 2130 31576 2164
rect 31524 2121 31576 2130
rect 31524 2092 31576 2109
rect 31524 2058 31533 2092
rect 31533 2058 31567 2092
rect 31567 2058 31576 2092
rect 31524 2057 31576 2058
rect 31524 2020 31576 2045
rect 31524 1993 31533 2020
rect 31533 1993 31567 2020
rect 31567 1993 31576 2020
rect 31524 1948 31576 1981
rect 31524 1929 31533 1948
rect 31533 1929 31567 1948
rect 31567 1929 31576 1948
rect 31524 1914 31533 1917
rect 31533 1914 31567 1917
rect 31567 1914 31576 1917
rect 31524 1876 31576 1914
rect 31524 1865 31533 1876
rect 31533 1865 31567 1876
rect 31567 1865 31576 1876
rect 31524 1842 31533 1853
rect 31533 1842 31567 1853
rect 31567 1842 31576 1853
rect 31524 1804 31576 1842
rect 31524 1801 31533 1804
rect 31533 1801 31567 1804
rect 31567 1801 31576 1804
rect 31524 1770 31533 1789
rect 31533 1770 31567 1789
rect 31567 1770 31576 1789
rect 31524 1737 31576 1770
rect 31524 1698 31533 1725
rect 31533 1698 31567 1725
rect 31567 1698 31576 1725
rect 31524 1673 31576 1698
rect 31524 1660 31576 1661
rect 31524 1626 31533 1660
rect 31533 1626 31567 1660
rect 31567 1626 31576 1660
rect 31524 1609 31576 1626
rect 31524 1588 31576 1597
rect 31524 1554 31533 1588
rect 31533 1554 31567 1588
rect 31567 1554 31576 1588
rect 31524 1545 31576 1554
rect 31524 1516 31576 1533
rect 31524 1482 31533 1516
rect 31533 1482 31567 1516
rect 31567 1482 31576 1516
rect 31524 1481 31576 1482
rect 31524 1444 31576 1469
rect 31524 1417 31533 1444
rect 31533 1417 31567 1444
rect 31567 1417 31576 1444
rect 31524 1372 31576 1405
rect 31524 1353 31533 1372
rect 31533 1353 31567 1372
rect 31567 1353 31576 1372
rect 31524 1338 31533 1341
rect 31533 1338 31567 1341
rect 31567 1338 31576 1341
rect 31524 1300 31576 1338
rect 31524 1289 31533 1300
rect 31533 1289 31567 1300
rect 31567 1289 31576 1300
rect 31524 1266 31533 1277
rect 31533 1266 31567 1277
rect 31567 1266 31576 1277
rect 31524 1228 31576 1266
rect 31524 1225 31533 1228
rect 31533 1225 31567 1228
rect 31567 1225 31576 1228
rect 31524 1194 31533 1213
rect 31533 1194 31567 1213
rect 31567 1194 31576 1213
rect 31524 1161 31576 1194
rect 31620 3100 31672 3133
rect 31620 3081 31629 3100
rect 31629 3081 31663 3100
rect 31663 3081 31672 3100
rect 31620 3066 31629 3069
rect 31629 3066 31663 3069
rect 31663 3066 31672 3069
rect 31620 3028 31672 3066
rect 31620 3017 31629 3028
rect 31629 3017 31663 3028
rect 31663 3017 31672 3028
rect 31620 2994 31629 3005
rect 31629 2994 31663 3005
rect 31663 2994 31672 3005
rect 31620 2956 31672 2994
rect 31620 2953 31629 2956
rect 31629 2953 31663 2956
rect 31663 2953 31672 2956
rect 31620 2922 31629 2941
rect 31629 2922 31663 2941
rect 31663 2922 31672 2941
rect 31620 2889 31672 2922
rect 31620 2850 31629 2877
rect 31629 2850 31663 2877
rect 31663 2850 31672 2877
rect 31620 2825 31672 2850
rect 31620 2812 31672 2813
rect 31620 2778 31629 2812
rect 31629 2778 31663 2812
rect 31663 2778 31672 2812
rect 31620 2761 31672 2778
rect 31620 2740 31672 2749
rect 31620 2706 31629 2740
rect 31629 2706 31663 2740
rect 31663 2706 31672 2740
rect 31620 2697 31672 2706
rect 31620 2668 31672 2685
rect 31620 2634 31629 2668
rect 31629 2634 31663 2668
rect 31663 2634 31672 2668
rect 31620 2633 31672 2634
rect 31620 2596 31672 2621
rect 31620 2569 31629 2596
rect 31629 2569 31663 2596
rect 31663 2569 31672 2596
rect 31620 2524 31672 2557
rect 31620 2505 31629 2524
rect 31629 2505 31663 2524
rect 31663 2505 31672 2524
rect 31620 2490 31629 2493
rect 31629 2490 31663 2493
rect 31663 2490 31672 2493
rect 31620 2452 31672 2490
rect 31620 2441 31629 2452
rect 31629 2441 31663 2452
rect 31663 2441 31672 2452
rect 31620 2418 31629 2429
rect 31629 2418 31663 2429
rect 31663 2418 31672 2429
rect 31620 2380 31672 2418
rect 31620 2377 31629 2380
rect 31629 2377 31663 2380
rect 31663 2377 31672 2380
rect 31620 2346 31629 2365
rect 31629 2346 31663 2365
rect 31663 2346 31672 2365
rect 31620 2313 31672 2346
rect 31620 2274 31629 2301
rect 31629 2274 31663 2301
rect 31663 2274 31672 2301
rect 31620 2249 31672 2274
rect 31620 2236 31672 2237
rect 31620 2202 31629 2236
rect 31629 2202 31663 2236
rect 31663 2202 31672 2236
rect 31620 2185 31672 2202
rect 31620 2164 31672 2173
rect 31620 2130 31629 2164
rect 31629 2130 31663 2164
rect 31663 2130 31672 2164
rect 31620 2121 31672 2130
rect 31620 2092 31672 2109
rect 31620 2058 31629 2092
rect 31629 2058 31663 2092
rect 31663 2058 31672 2092
rect 31620 2057 31672 2058
rect 31620 2020 31672 2045
rect 31620 1993 31629 2020
rect 31629 1993 31663 2020
rect 31663 1993 31672 2020
rect 31620 1948 31672 1981
rect 31620 1929 31629 1948
rect 31629 1929 31663 1948
rect 31663 1929 31672 1948
rect 31620 1914 31629 1917
rect 31629 1914 31663 1917
rect 31663 1914 31672 1917
rect 31620 1876 31672 1914
rect 31620 1865 31629 1876
rect 31629 1865 31663 1876
rect 31663 1865 31672 1876
rect 31620 1842 31629 1853
rect 31629 1842 31663 1853
rect 31663 1842 31672 1853
rect 31620 1804 31672 1842
rect 31620 1801 31629 1804
rect 31629 1801 31663 1804
rect 31663 1801 31672 1804
rect 31620 1770 31629 1789
rect 31629 1770 31663 1789
rect 31663 1770 31672 1789
rect 31620 1737 31672 1770
rect 31620 1698 31629 1725
rect 31629 1698 31663 1725
rect 31663 1698 31672 1725
rect 31620 1673 31672 1698
rect 31620 1660 31672 1661
rect 31620 1626 31629 1660
rect 31629 1626 31663 1660
rect 31663 1626 31672 1660
rect 31620 1609 31672 1626
rect 31620 1588 31672 1597
rect 31620 1554 31629 1588
rect 31629 1554 31663 1588
rect 31663 1554 31672 1588
rect 31620 1545 31672 1554
rect 31620 1516 31672 1533
rect 31620 1482 31629 1516
rect 31629 1482 31663 1516
rect 31663 1482 31672 1516
rect 31620 1481 31672 1482
rect 31620 1444 31672 1469
rect 31620 1417 31629 1444
rect 31629 1417 31663 1444
rect 31663 1417 31672 1444
rect 31620 1372 31672 1405
rect 31620 1353 31629 1372
rect 31629 1353 31663 1372
rect 31663 1353 31672 1372
rect 31620 1338 31629 1341
rect 31629 1338 31663 1341
rect 31663 1338 31672 1341
rect 31620 1300 31672 1338
rect 31620 1289 31629 1300
rect 31629 1289 31663 1300
rect 31663 1289 31672 1300
rect 31620 1266 31629 1277
rect 31629 1266 31663 1277
rect 31663 1266 31672 1277
rect 31620 1228 31672 1266
rect 31620 1225 31629 1228
rect 31629 1225 31663 1228
rect 31663 1225 31672 1228
rect 31620 1194 31629 1213
rect 31629 1194 31663 1213
rect 31663 1194 31672 1213
rect 31620 1161 31672 1194
rect 31716 3100 31768 3133
rect 31716 3081 31725 3100
rect 31725 3081 31759 3100
rect 31759 3081 31768 3100
rect 31716 3066 31725 3069
rect 31725 3066 31759 3069
rect 31759 3066 31768 3069
rect 31716 3028 31768 3066
rect 31716 3017 31725 3028
rect 31725 3017 31759 3028
rect 31759 3017 31768 3028
rect 31716 2994 31725 3005
rect 31725 2994 31759 3005
rect 31759 2994 31768 3005
rect 31716 2956 31768 2994
rect 31716 2953 31725 2956
rect 31725 2953 31759 2956
rect 31759 2953 31768 2956
rect 31716 2922 31725 2941
rect 31725 2922 31759 2941
rect 31759 2922 31768 2941
rect 31716 2889 31768 2922
rect 31716 2850 31725 2877
rect 31725 2850 31759 2877
rect 31759 2850 31768 2877
rect 31716 2825 31768 2850
rect 31716 2812 31768 2813
rect 31716 2778 31725 2812
rect 31725 2778 31759 2812
rect 31759 2778 31768 2812
rect 31716 2761 31768 2778
rect 31716 2740 31768 2749
rect 31716 2706 31725 2740
rect 31725 2706 31759 2740
rect 31759 2706 31768 2740
rect 31716 2697 31768 2706
rect 31716 2668 31768 2685
rect 31716 2634 31725 2668
rect 31725 2634 31759 2668
rect 31759 2634 31768 2668
rect 31716 2633 31768 2634
rect 31716 2596 31768 2621
rect 31716 2569 31725 2596
rect 31725 2569 31759 2596
rect 31759 2569 31768 2596
rect 31716 2524 31768 2557
rect 31716 2505 31725 2524
rect 31725 2505 31759 2524
rect 31759 2505 31768 2524
rect 31716 2490 31725 2493
rect 31725 2490 31759 2493
rect 31759 2490 31768 2493
rect 31716 2452 31768 2490
rect 31716 2441 31725 2452
rect 31725 2441 31759 2452
rect 31759 2441 31768 2452
rect 31716 2418 31725 2429
rect 31725 2418 31759 2429
rect 31759 2418 31768 2429
rect 31716 2380 31768 2418
rect 31716 2377 31725 2380
rect 31725 2377 31759 2380
rect 31759 2377 31768 2380
rect 31716 2346 31725 2365
rect 31725 2346 31759 2365
rect 31759 2346 31768 2365
rect 31716 2313 31768 2346
rect 31716 2274 31725 2301
rect 31725 2274 31759 2301
rect 31759 2274 31768 2301
rect 31716 2249 31768 2274
rect 31716 2236 31768 2237
rect 31716 2202 31725 2236
rect 31725 2202 31759 2236
rect 31759 2202 31768 2236
rect 31716 2185 31768 2202
rect 31716 2164 31768 2173
rect 31716 2130 31725 2164
rect 31725 2130 31759 2164
rect 31759 2130 31768 2164
rect 31716 2121 31768 2130
rect 31716 2092 31768 2109
rect 31716 2058 31725 2092
rect 31725 2058 31759 2092
rect 31759 2058 31768 2092
rect 31716 2057 31768 2058
rect 31716 2020 31768 2045
rect 31716 1993 31725 2020
rect 31725 1993 31759 2020
rect 31759 1993 31768 2020
rect 31716 1948 31768 1981
rect 31716 1929 31725 1948
rect 31725 1929 31759 1948
rect 31759 1929 31768 1948
rect 31716 1914 31725 1917
rect 31725 1914 31759 1917
rect 31759 1914 31768 1917
rect 31716 1876 31768 1914
rect 31716 1865 31725 1876
rect 31725 1865 31759 1876
rect 31759 1865 31768 1876
rect 31716 1842 31725 1853
rect 31725 1842 31759 1853
rect 31759 1842 31768 1853
rect 31716 1804 31768 1842
rect 31716 1801 31725 1804
rect 31725 1801 31759 1804
rect 31759 1801 31768 1804
rect 31716 1770 31725 1789
rect 31725 1770 31759 1789
rect 31759 1770 31768 1789
rect 31716 1737 31768 1770
rect 31716 1698 31725 1725
rect 31725 1698 31759 1725
rect 31759 1698 31768 1725
rect 31716 1673 31768 1698
rect 31716 1660 31768 1661
rect 31716 1626 31725 1660
rect 31725 1626 31759 1660
rect 31759 1626 31768 1660
rect 31716 1609 31768 1626
rect 31716 1588 31768 1597
rect 31716 1554 31725 1588
rect 31725 1554 31759 1588
rect 31759 1554 31768 1588
rect 31716 1545 31768 1554
rect 31716 1516 31768 1533
rect 31716 1482 31725 1516
rect 31725 1482 31759 1516
rect 31759 1482 31768 1516
rect 31716 1481 31768 1482
rect 31716 1444 31768 1469
rect 31716 1417 31725 1444
rect 31725 1417 31759 1444
rect 31759 1417 31768 1444
rect 31716 1372 31768 1405
rect 31716 1353 31725 1372
rect 31725 1353 31759 1372
rect 31759 1353 31768 1372
rect 31716 1338 31725 1341
rect 31725 1338 31759 1341
rect 31759 1338 31768 1341
rect 31716 1300 31768 1338
rect 31716 1289 31725 1300
rect 31725 1289 31759 1300
rect 31759 1289 31768 1300
rect 31716 1266 31725 1277
rect 31725 1266 31759 1277
rect 31759 1266 31768 1277
rect 31716 1228 31768 1266
rect 31716 1225 31725 1228
rect 31725 1225 31759 1228
rect 31759 1225 31768 1228
rect 31716 1194 31725 1213
rect 31725 1194 31759 1213
rect 31759 1194 31768 1213
rect 31716 1161 31768 1194
rect 31812 3100 31864 3133
rect 31812 3081 31821 3100
rect 31821 3081 31855 3100
rect 31855 3081 31864 3100
rect 31812 3066 31821 3069
rect 31821 3066 31855 3069
rect 31855 3066 31864 3069
rect 31812 3028 31864 3066
rect 31812 3017 31821 3028
rect 31821 3017 31855 3028
rect 31855 3017 31864 3028
rect 31812 2994 31821 3005
rect 31821 2994 31855 3005
rect 31855 2994 31864 3005
rect 31812 2956 31864 2994
rect 31812 2953 31821 2956
rect 31821 2953 31855 2956
rect 31855 2953 31864 2956
rect 31812 2922 31821 2941
rect 31821 2922 31855 2941
rect 31855 2922 31864 2941
rect 31812 2889 31864 2922
rect 31812 2850 31821 2877
rect 31821 2850 31855 2877
rect 31855 2850 31864 2877
rect 31812 2825 31864 2850
rect 31812 2812 31864 2813
rect 31812 2778 31821 2812
rect 31821 2778 31855 2812
rect 31855 2778 31864 2812
rect 31812 2761 31864 2778
rect 31812 2740 31864 2749
rect 31812 2706 31821 2740
rect 31821 2706 31855 2740
rect 31855 2706 31864 2740
rect 31812 2697 31864 2706
rect 31812 2668 31864 2685
rect 31812 2634 31821 2668
rect 31821 2634 31855 2668
rect 31855 2634 31864 2668
rect 31812 2633 31864 2634
rect 31812 2596 31864 2621
rect 31812 2569 31821 2596
rect 31821 2569 31855 2596
rect 31855 2569 31864 2596
rect 31812 2524 31864 2557
rect 31812 2505 31821 2524
rect 31821 2505 31855 2524
rect 31855 2505 31864 2524
rect 31812 2490 31821 2493
rect 31821 2490 31855 2493
rect 31855 2490 31864 2493
rect 31812 2452 31864 2490
rect 31812 2441 31821 2452
rect 31821 2441 31855 2452
rect 31855 2441 31864 2452
rect 31812 2418 31821 2429
rect 31821 2418 31855 2429
rect 31855 2418 31864 2429
rect 31812 2380 31864 2418
rect 31812 2377 31821 2380
rect 31821 2377 31855 2380
rect 31855 2377 31864 2380
rect 31812 2346 31821 2365
rect 31821 2346 31855 2365
rect 31855 2346 31864 2365
rect 31812 2313 31864 2346
rect 31812 2274 31821 2301
rect 31821 2274 31855 2301
rect 31855 2274 31864 2301
rect 31812 2249 31864 2274
rect 31812 2236 31864 2237
rect 31812 2202 31821 2236
rect 31821 2202 31855 2236
rect 31855 2202 31864 2236
rect 31812 2185 31864 2202
rect 31812 2164 31864 2173
rect 31812 2130 31821 2164
rect 31821 2130 31855 2164
rect 31855 2130 31864 2164
rect 31812 2121 31864 2130
rect 31812 2092 31864 2109
rect 31812 2058 31821 2092
rect 31821 2058 31855 2092
rect 31855 2058 31864 2092
rect 31812 2057 31864 2058
rect 31812 2020 31864 2045
rect 31812 1993 31821 2020
rect 31821 1993 31855 2020
rect 31855 1993 31864 2020
rect 31812 1948 31864 1981
rect 31812 1929 31821 1948
rect 31821 1929 31855 1948
rect 31855 1929 31864 1948
rect 31812 1914 31821 1917
rect 31821 1914 31855 1917
rect 31855 1914 31864 1917
rect 31812 1876 31864 1914
rect 31812 1865 31821 1876
rect 31821 1865 31855 1876
rect 31855 1865 31864 1876
rect 31812 1842 31821 1853
rect 31821 1842 31855 1853
rect 31855 1842 31864 1853
rect 31812 1804 31864 1842
rect 31812 1801 31821 1804
rect 31821 1801 31855 1804
rect 31855 1801 31864 1804
rect 31812 1770 31821 1789
rect 31821 1770 31855 1789
rect 31855 1770 31864 1789
rect 31812 1737 31864 1770
rect 31812 1698 31821 1725
rect 31821 1698 31855 1725
rect 31855 1698 31864 1725
rect 31812 1673 31864 1698
rect 31812 1660 31864 1661
rect 31812 1626 31821 1660
rect 31821 1626 31855 1660
rect 31855 1626 31864 1660
rect 31812 1609 31864 1626
rect 31812 1588 31864 1597
rect 31812 1554 31821 1588
rect 31821 1554 31855 1588
rect 31855 1554 31864 1588
rect 31812 1545 31864 1554
rect 31812 1516 31864 1533
rect 31812 1482 31821 1516
rect 31821 1482 31855 1516
rect 31855 1482 31864 1516
rect 31812 1481 31864 1482
rect 31812 1444 31864 1469
rect 31812 1417 31821 1444
rect 31821 1417 31855 1444
rect 31855 1417 31864 1444
rect 31812 1372 31864 1405
rect 31812 1353 31821 1372
rect 31821 1353 31855 1372
rect 31855 1353 31864 1372
rect 31812 1338 31821 1341
rect 31821 1338 31855 1341
rect 31855 1338 31864 1341
rect 31812 1300 31864 1338
rect 31812 1289 31821 1300
rect 31821 1289 31855 1300
rect 31855 1289 31864 1300
rect 31812 1266 31821 1277
rect 31821 1266 31855 1277
rect 31855 1266 31864 1277
rect 31812 1228 31864 1266
rect 31812 1225 31821 1228
rect 31821 1225 31855 1228
rect 31855 1225 31864 1228
rect 31812 1194 31821 1213
rect 31821 1194 31855 1213
rect 31855 1194 31864 1213
rect 31812 1161 31864 1194
rect 31908 3100 31960 3133
rect 31908 3081 31917 3100
rect 31917 3081 31951 3100
rect 31951 3081 31960 3100
rect 31908 3066 31917 3069
rect 31917 3066 31951 3069
rect 31951 3066 31960 3069
rect 31908 3028 31960 3066
rect 31908 3017 31917 3028
rect 31917 3017 31951 3028
rect 31951 3017 31960 3028
rect 31908 2994 31917 3005
rect 31917 2994 31951 3005
rect 31951 2994 31960 3005
rect 31908 2956 31960 2994
rect 31908 2953 31917 2956
rect 31917 2953 31951 2956
rect 31951 2953 31960 2956
rect 31908 2922 31917 2941
rect 31917 2922 31951 2941
rect 31951 2922 31960 2941
rect 31908 2889 31960 2922
rect 31908 2850 31917 2877
rect 31917 2850 31951 2877
rect 31951 2850 31960 2877
rect 31908 2825 31960 2850
rect 31908 2812 31960 2813
rect 31908 2778 31917 2812
rect 31917 2778 31951 2812
rect 31951 2778 31960 2812
rect 31908 2761 31960 2778
rect 31908 2740 31960 2749
rect 31908 2706 31917 2740
rect 31917 2706 31951 2740
rect 31951 2706 31960 2740
rect 31908 2697 31960 2706
rect 31908 2668 31960 2685
rect 31908 2634 31917 2668
rect 31917 2634 31951 2668
rect 31951 2634 31960 2668
rect 31908 2633 31960 2634
rect 31908 2596 31960 2621
rect 31908 2569 31917 2596
rect 31917 2569 31951 2596
rect 31951 2569 31960 2596
rect 31908 2524 31960 2557
rect 31908 2505 31917 2524
rect 31917 2505 31951 2524
rect 31951 2505 31960 2524
rect 31908 2490 31917 2493
rect 31917 2490 31951 2493
rect 31951 2490 31960 2493
rect 31908 2452 31960 2490
rect 31908 2441 31917 2452
rect 31917 2441 31951 2452
rect 31951 2441 31960 2452
rect 31908 2418 31917 2429
rect 31917 2418 31951 2429
rect 31951 2418 31960 2429
rect 31908 2380 31960 2418
rect 31908 2377 31917 2380
rect 31917 2377 31951 2380
rect 31951 2377 31960 2380
rect 31908 2346 31917 2365
rect 31917 2346 31951 2365
rect 31951 2346 31960 2365
rect 31908 2313 31960 2346
rect 31908 2274 31917 2301
rect 31917 2274 31951 2301
rect 31951 2274 31960 2301
rect 31908 2249 31960 2274
rect 31908 2236 31960 2237
rect 31908 2202 31917 2236
rect 31917 2202 31951 2236
rect 31951 2202 31960 2236
rect 31908 2185 31960 2202
rect 31908 2164 31960 2173
rect 31908 2130 31917 2164
rect 31917 2130 31951 2164
rect 31951 2130 31960 2164
rect 31908 2121 31960 2130
rect 31908 2092 31960 2109
rect 31908 2058 31917 2092
rect 31917 2058 31951 2092
rect 31951 2058 31960 2092
rect 31908 2057 31960 2058
rect 31908 2020 31960 2045
rect 31908 1993 31917 2020
rect 31917 1993 31951 2020
rect 31951 1993 31960 2020
rect 31908 1948 31960 1981
rect 31908 1929 31917 1948
rect 31917 1929 31951 1948
rect 31951 1929 31960 1948
rect 31908 1914 31917 1917
rect 31917 1914 31951 1917
rect 31951 1914 31960 1917
rect 31908 1876 31960 1914
rect 31908 1865 31917 1876
rect 31917 1865 31951 1876
rect 31951 1865 31960 1876
rect 31908 1842 31917 1853
rect 31917 1842 31951 1853
rect 31951 1842 31960 1853
rect 31908 1804 31960 1842
rect 31908 1801 31917 1804
rect 31917 1801 31951 1804
rect 31951 1801 31960 1804
rect 31908 1770 31917 1789
rect 31917 1770 31951 1789
rect 31951 1770 31960 1789
rect 31908 1737 31960 1770
rect 31908 1698 31917 1725
rect 31917 1698 31951 1725
rect 31951 1698 31960 1725
rect 31908 1673 31960 1698
rect 31908 1660 31960 1661
rect 31908 1626 31917 1660
rect 31917 1626 31951 1660
rect 31951 1626 31960 1660
rect 31908 1609 31960 1626
rect 31908 1588 31960 1597
rect 31908 1554 31917 1588
rect 31917 1554 31951 1588
rect 31951 1554 31960 1588
rect 31908 1545 31960 1554
rect 31908 1516 31960 1533
rect 31908 1482 31917 1516
rect 31917 1482 31951 1516
rect 31951 1482 31960 1516
rect 31908 1481 31960 1482
rect 31908 1444 31960 1469
rect 31908 1417 31917 1444
rect 31917 1417 31951 1444
rect 31951 1417 31960 1444
rect 31908 1372 31960 1405
rect 31908 1353 31917 1372
rect 31917 1353 31951 1372
rect 31951 1353 31960 1372
rect 31908 1338 31917 1341
rect 31917 1338 31951 1341
rect 31951 1338 31960 1341
rect 31908 1300 31960 1338
rect 31908 1289 31917 1300
rect 31917 1289 31951 1300
rect 31951 1289 31960 1300
rect 31908 1266 31917 1277
rect 31917 1266 31951 1277
rect 31951 1266 31960 1277
rect 31908 1228 31960 1266
rect 31908 1225 31917 1228
rect 31917 1225 31951 1228
rect 31951 1225 31960 1228
rect 31908 1194 31917 1213
rect 31917 1194 31951 1213
rect 31951 1194 31960 1213
rect 31908 1161 31960 1194
rect 32004 3100 32056 3133
rect 32004 3081 32013 3100
rect 32013 3081 32047 3100
rect 32047 3081 32056 3100
rect 32004 3066 32013 3069
rect 32013 3066 32047 3069
rect 32047 3066 32056 3069
rect 32004 3028 32056 3066
rect 32004 3017 32013 3028
rect 32013 3017 32047 3028
rect 32047 3017 32056 3028
rect 32004 2994 32013 3005
rect 32013 2994 32047 3005
rect 32047 2994 32056 3005
rect 32004 2956 32056 2994
rect 32004 2953 32013 2956
rect 32013 2953 32047 2956
rect 32047 2953 32056 2956
rect 32004 2922 32013 2941
rect 32013 2922 32047 2941
rect 32047 2922 32056 2941
rect 32004 2889 32056 2922
rect 32004 2850 32013 2877
rect 32013 2850 32047 2877
rect 32047 2850 32056 2877
rect 32004 2825 32056 2850
rect 32004 2812 32056 2813
rect 32004 2778 32013 2812
rect 32013 2778 32047 2812
rect 32047 2778 32056 2812
rect 32004 2761 32056 2778
rect 32004 2740 32056 2749
rect 32004 2706 32013 2740
rect 32013 2706 32047 2740
rect 32047 2706 32056 2740
rect 32004 2697 32056 2706
rect 32004 2668 32056 2685
rect 32004 2634 32013 2668
rect 32013 2634 32047 2668
rect 32047 2634 32056 2668
rect 32004 2633 32056 2634
rect 32004 2596 32056 2621
rect 32004 2569 32013 2596
rect 32013 2569 32047 2596
rect 32047 2569 32056 2596
rect 32004 2524 32056 2557
rect 32004 2505 32013 2524
rect 32013 2505 32047 2524
rect 32047 2505 32056 2524
rect 32004 2490 32013 2493
rect 32013 2490 32047 2493
rect 32047 2490 32056 2493
rect 32004 2452 32056 2490
rect 32004 2441 32013 2452
rect 32013 2441 32047 2452
rect 32047 2441 32056 2452
rect 32004 2418 32013 2429
rect 32013 2418 32047 2429
rect 32047 2418 32056 2429
rect 32004 2380 32056 2418
rect 32004 2377 32013 2380
rect 32013 2377 32047 2380
rect 32047 2377 32056 2380
rect 32004 2346 32013 2365
rect 32013 2346 32047 2365
rect 32047 2346 32056 2365
rect 32004 2313 32056 2346
rect 32004 2274 32013 2301
rect 32013 2274 32047 2301
rect 32047 2274 32056 2301
rect 32004 2249 32056 2274
rect 32004 2236 32056 2237
rect 32004 2202 32013 2236
rect 32013 2202 32047 2236
rect 32047 2202 32056 2236
rect 32004 2185 32056 2202
rect 32004 2164 32056 2173
rect 32004 2130 32013 2164
rect 32013 2130 32047 2164
rect 32047 2130 32056 2164
rect 32004 2121 32056 2130
rect 32004 2092 32056 2109
rect 32004 2058 32013 2092
rect 32013 2058 32047 2092
rect 32047 2058 32056 2092
rect 32004 2057 32056 2058
rect 32004 2020 32056 2045
rect 32004 1993 32013 2020
rect 32013 1993 32047 2020
rect 32047 1993 32056 2020
rect 32004 1948 32056 1981
rect 32004 1929 32013 1948
rect 32013 1929 32047 1948
rect 32047 1929 32056 1948
rect 32004 1914 32013 1917
rect 32013 1914 32047 1917
rect 32047 1914 32056 1917
rect 32004 1876 32056 1914
rect 32004 1865 32013 1876
rect 32013 1865 32047 1876
rect 32047 1865 32056 1876
rect 32004 1842 32013 1853
rect 32013 1842 32047 1853
rect 32047 1842 32056 1853
rect 32004 1804 32056 1842
rect 32004 1801 32013 1804
rect 32013 1801 32047 1804
rect 32047 1801 32056 1804
rect 32004 1770 32013 1789
rect 32013 1770 32047 1789
rect 32047 1770 32056 1789
rect 32004 1737 32056 1770
rect 32004 1698 32013 1725
rect 32013 1698 32047 1725
rect 32047 1698 32056 1725
rect 32004 1673 32056 1698
rect 32004 1660 32056 1661
rect 32004 1626 32013 1660
rect 32013 1626 32047 1660
rect 32047 1626 32056 1660
rect 32004 1609 32056 1626
rect 32004 1588 32056 1597
rect 32004 1554 32013 1588
rect 32013 1554 32047 1588
rect 32047 1554 32056 1588
rect 32004 1545 32056 1554
rect 32004 1516 32056 1533
rect 32004 1482 32013 1516
rect 32013 1482 32047 1516
rect 32047 1482 32056 1516
rect 32004 1481 32056 1482
rect 32004 1444 32056 1469
rect 32004 1417 32013 1444
rect 32013 1417 32047 1444
rect 32047 1417 32056 1444
rect 32004 1372 32056 1405
rect 32004 1353 32013 1372
rect 32013 1353 32047 1372
rect 32047 1353 32056 1372
rect 32004 1338 32013 1341
rect 32013 1338 32047 1341
rect 32047 1338 32056 1341
rect 32004 1300 32056 1338
rect 32004 1289 32013 1300
rect 32013 1289 32047 1300
rect 32047 1289 32056 1300
rect 32004 1266 32013 1277
rect 32013 1266 32047 1277
rect 32047 1266 32056 1277
rect 32004 1228 32056 1266
rect 32004 1225 32013 1228
rect 32013 1225 32047 1228
rect 32047 1225 32056 1228
rect 32004 1194 32013 1213
rect 32013 1194 32047 1213
rect 32047 1194 32056 1213
rect 32004 1161 32056 1194
rect 32100 3100 32152 3133
rect 32100 3081 32109 3100
rect 32109 3081 32143 3100
rect 32143 3081 32152 3100
rect 32100 3066 32109 3069
rect 32109 3066 32143 3069
rect 32143 3066 32152 3069
rect 32100 3028 32152 3066
rect 32100 3017 32109 3028
rect 32109 3017 32143 3028
rect 32143 3017 32152 3028
rect 32100 2994 32109 3005
rect 32109 2994 32143 3005
rect 32143 2994 32152 3005
rect 32100 2956 32152 2994
rect 32100 2953 32109 2956
rect 32109 2953 32143 2956
rect 32143 2953 32152 2956
rect 32100 2922 32109 2941
rect 32109 2922 32143 2941
rect 32143 2922 32152 2941
rect 32100 2889 32152 2922
rect 32100 2850 32109 2877
rect 32109 2850 32143 2877
rect 32143 2850 32152 2877
rect 32100 2825 32152 2850
rect 32100 2812 32152 2813
rect 32100 2778 32109 2812
rect 32109 2778 32143 2812
rect 32143 2778 32152 2812
rect 32100 2761 32152 2778
rect 32100 2740 32152 2749
rect 32100 2706 32109 2740
rect 32109 2706 32143 2740
rect 32143 2706 32152 2740
rect 32100 2697 32152 2706
rect 32100 2668 32152 2685
rect 32100 2634 32109 2668
rect 32109 2634 32143 2668
rect 32143 2634 32152 2668
rect 32100 2633 32152 2634
rect 32100 2596 32152 2621
rect 32100 2569 32109 2596
rect 32109 2569 32143 2596
rect 32143 2569 32152 2596
rect 32100 2524 32152 2557
rect 32100 2505 32109 2524
rect 32109 2505 32143 2524
rect 32143 2505 32152 2524
rect 32100 2490 32109 2493
rect 32109 2490 32143 2493
rect 32143 2490 32152 2493
rect 32100 2452 32152 2490
rect 32100 2441 32109 2452
rect 32109 2441 32143 2452
rect 32143 2441 32152 2452
rect 32100 2418 32109 2429
rect 32109 2418 32143 2429
rect 32143 2418 32152 2429
rect 32100 2380 32152 2418
rect 32100 2377 32109 2380
rect 32109 2377 32143 2380
rect 32143 2377 32152 2380
rect 32100 2346 32109 2365
rect 32109 2346 32143 2365
rect 32143 2346 32152 2365
rect 32100 2313 32152 2346
rect 32100 2274 32109 2301
rect 32109 2274 32143 2301
rect 32143 2274 32152 2301
rect 32100 2249 32152 2274
rect 32100 2236 32152 2237
rect 32100 2202 32109 2236
rect 32109 2202 32143 2236
rect 32143 2202 32152 2236
rect 32100 2185 32152 2202
rect 32100 2164 32152 2173
rect 32100 2130 32109 2164
rect 32109 2130 32143 2164
rect 32143 2130 32152 2164
rect 32100 2121 32152 2130
rect 32100 2092 32152 2109
rect 32100 2058 32109 2092
rect 32109 2058 32143 2092
rect 32143 2058 32152 2092
rect 32100 2057 32152 2058
rect 32100 2020 32152 2045
rect 32100 1993 32109 2020
rect 32109 1993 32143 2020
rect 32143 1993 32152 2020
rect 32100 1948 32152 1981
rect 32100 1929 32109 1948
rect 32109 1929 32143 1948
rect 32143 1929 32152 1948
rect 32100 1914 32109 1917
rect 32109 1914 32143 1917
rect 32143 1914 32152 1917
rect 32100 1876 32152 1914
rect 32100 1865 32109 1876
rect 32109 1865 32143 1876
rect 32143 1865 32152 1876
rect 32100 1842 32109 1853
rect 32109 1842 32143 1853
rect 32143 1842 32152 1853
rect 32100 1804 32152 1842
rect 32100 1801 32109 1804
rect 32109 1801 32143 1804
rect 32143 1801 32152 1804
rect 32100 1770 32109 1789
rect 32109 1770 32143 1789
rect 32143 1770 32152 1789
rect 32100 1737 32152 1770
rect 32100 1698 32109 1725
rect 32109 1698 32143 1725
rect 32143 1698 32152 1725
rect 32100 1673 32152 1698
rect 32100 1660 32152 1661
rect 32100 1626 32109 1660
rect 32109 1626 32143 1660
rect 32143 1626 32152 1660
rect 32100 1609 32152 1626
rect 32100 1588 32152 1597
rect 32100 1554 32109 1588
rect 32109 1554 32143 1588
rect 32143 1554 32152 1588
rect 32100 1545 32152 1554
rect 32100 1516 32152 1533
rect 32100 1482 32109 1516
rect 32109 1482 32143 1516
rect 32143 1482 32152 1516
rect 32100 1481 32152 1482
rect 32100 1444 32152 1469
rect 32100 1417 32109 1444
rect 32109 1417 32143 1444
rect 32143 1417 32152 1444
rect 32100 1372 32152 1405
rect 32100 1353 32109 1372
rect 32109 1353 32143 1372
rect 32143 1353 32152 1372
rect 32100 1338 32109 1341
rect 32109 1338 32143 1341
rect 32143 1338 32152 1341
rect 32100 1300 32152 1338
rect 32100 1289 32109 1300
rect 32109 1289 32143 1300
rect 32143 1289 32152 1300
rect 32100 1266 32109 1277
rect 32109 1266 32143 1277
rect 32143 1266 32152 1277
rect 32100 1228 32152 1266
rect 32100 1225 32109 1228
rect 32109 1225 32143 1228
rect 32143 1225 32152 1228
rect 32100 1194 32109 1213
rect 32109 1194 32143 1213
rect 32143 1194 32152 1213
rect 32100 1161 32152 1194
rect 32196 3100 32248 3133
rect 32196 3081 32205 3100
rect 32205 3081 32239 3100
rect 32239 3081 32248 3100
rect 32196 3066 32205 3069
rect 32205 3066 32239 3069
rect 32239 3066 32248 3069
rect 32196 3028 32248 3066
rect 32196 3017 32205 3028
rect 32205 3017 32239 3028
rect 32239 3017 32248 3028
rect 32196 2994 32205 3005
rect 32205 2994 32239 3005
rect 32239 2994 32248 3005
rect 32196 2956 32248 2994
rect 32196 2953 32205 2956
rect 32205 2953 32239 2956
rect 32239 2953 32248 2956
rect 32196 2922 32205 2941
rect 32205 2922 32239 2941
rect 32239 2922 32248 2941
rect 32196 2889 32248 2922
rect 32196 2850 32205 2877
rect 32205 2850 32239 2877
rect 32239 2850 32248 2877
rect 32196 2825 32248 2850
rect 32196 2812 32248 2813
rect 32196 2778 32205 2812
rect 32205 2778 32239 2812
rect 32239 2778 32248 2812
rect 32196 2761 32248 2778
rect 32196 2740 32248 2749
rect 32196 2706 32205 2740
rect 32205 2706 32239 2740
rect 32239 2706 32248 2740
rect 32196 2697 32248 2706
rect 32196 2668 32248 2685
rect 32196 2634 32205 2668
rect 32205 2634 32239 2668
rect 32239 2634 32248 2668
rect 32196 2633 32248 2634
rect 32196 2596 32248 2621
rect 32196 2569 32205 2596
rect 32205 2569 32239 2596
rect 32239 2569 32248 2596
rect 32196 2524 32248 2557
rect 32196 2505 32205 2524
rect 32205 2505 32239 2524
rect 32239 2505 32248 2524
rect 32196 2490 32205 2493
rect 32205 2490 32239 2493
rect 32239 2490 32248 2493
rect 32196 2452 32248 2490
rect 32196 2441 32205 2452
rect 32205 2441 32239 2452
rect 32239 2441 32248 2452
rect 32196 2418 32205 2429
rect 32205 2418 32239 2429
rect 32239 2418 32248 2429
rect 32196 2380 32248 2418
rect 32196 2377 32205 2380
rect 32205 2377 32239 2380
rect 32239 2377 32248 2380
rect 32196 2346 32205 2365
rect 32205 2346 32239 2365
rect 32239 2346 32248 2365
rect 32196 2313 32248 2346
rect 32196 2274 32205 2301
rect 32205 2274 32239 2301
rect 32239 2274 32248 2301
rect 32196 2249 32248 2274
rect 32196 2236 32248 2237
rect 32196 2202 32205 2236
rect 32205 2202 32239 2236
rect 32239 2202 32248 2236
rect 32196 2185 32248 2202
rect 32196 2164 32248 2173
rect 32196 2130 32205 2164
rect 32205 2130 32239 2164
rect 32239 2130 32248 2164
rect 32196 2121 32248 2130
rect 32196 2092 32248 2109
rect 32196 2058 32205 2092
rect 32205 2058 32239 2092
rect 32239 2058 32248 2092
rect 32196 2057 32248 2058
rect 32196 2020 32248 2045
rect 32196 1993 32205 2020
rect 32205 1993 32239 2020
rect 32239 1993 32248 2020
rect 32196 1948 32248 1981
rect 32196 1929 32205 1948
rect 32205 1929 32239 1948
rect 32239 1929 32248 1948
rect 32196 1914 32205 1917
rect 32205 1914 32239 1917
rect 32239 1914 32248 1917
rect 32196 1876 32248 1914
rect 32196 1865 32205 1876
rect 32205 1865 32239 1876
rect 32239 1865 32248 1876
rect 32196 1842 32205 1853
rect 32205 1842 32239 1853
rect 32239 1842 32248 1853
rect 32196 1804 32248 1842
rect 32196 1801 32205 1804
rect 32205 1801 32239 1804
rect 32239 1801 32248 1804
rect 32196 1770 32205 1789
rect 32205 1770 32239 1789
rect 32239 1770 32248 1789
rect 32196 1737 32248 1770
rect 32196 1698 32205 1725
rect 32205 1698 32239 1725
rect 32239 1698 32248 1725
rect 32196 1673 32248 1698
rect 32196 1660 32248 1661
rect 32196 1626 32205 1660
rect 32205 1626 32239 1660
rect 32239 1626 32248 1660
rect 32196 1609 32248 1626
rect 32196 1588 32248 1597
rect 32196 1554 32205 1588
rect 32205 1554 32239 1588
rect 32239 1554 32248 1588
rect 32196 1545 32248 1554
rect 32196 1516 32248 1533
rect 32196 1482 32205 1516
rect 32205 1482 32239 1516
rect 32239 1482 32248 1516
rect 32196 1481 32248 1482
rect 32196 1444 32248 1469
rect 32196 1417 32205 1444
rect 32205 1417 32239 1444
rect 32239 1417 32248 1444
rect 32196 1372 32248 1405
rect 32196 1353 32205 1372
rect 32205 1353 32239 1372
rect 32239 1353 32248 1372
rect 32196 1338 32205 1341
rect 32205 1338 32239 1341
rect 32239 1338 32248 1341
rect 32196 1300 32248 1338
rect 32196 1289 32205 1300
rect 32205 1289 32239 1300
rect 32239 1289 32248 1300
rect 32196 1266 32205 1277
rect 32205 1266 32239 1277
rect 32239 1266 32248 1277
rect 32196 1228 32248 1266
rect 32196 1225 32205 1228
rect 32205 1225 32239 1228
rect 32239 1225 32248 1228
rect 32196 1194 32205 1213
rect 32205 1194 32239 1213
rect 32239 1194 32248 1213
rect 32196 1161 32248 1194
rect 32292 3100 32344 3133
rect 32292 3081 32301 3100
rect 32301 3081 32335 3100
rect 32335 3081 32344 3100
rect 32292 3066 32301 3069
rect 32301 3066 32335 3069
rect 32335 3066 32344 3069
rect 32292 3028 32344 3066
rect 32292 3017 32301 3028
rect 32301 3017 32335 3028
rect 32335 3017 32344 3028
rect 32292 2994 32301 3005
rect 32301 2994 32335 3005
rect 32335 2994 32344 3005
rect 32292 2956 32344 2994
rect 32292 2953 32301 2956
rect 32301 2953 32335 2956
rect 32335 2953 32344 2956
rect 32292 2922 32301 2941
rect 32301 2922 32335 2941
rect 32335 2922 32344 2941
rect 32292 2889 32344 2922
rect 32292 2850 32301 2877
rect 32301 2850 32335 2877
rect 32335 2850 32344 2877
rect 32292 2825 32344 2850
rect 32292 2812 32344 2813
rect 32292 2778 32301 2812
rect 32301 2778 32335 2812
rect 32335 2778 32344 2812
rect 32292 2761 32344 2778
rect 32292 2740 32344 2749
rect 32292 2706 32301 2740
rect 32301 2706 32335 2740
rect 32335 2706 32344 2740
rect 32292 2697 32344 2706
rect 32292 2668 32344 2685
rect 32292 2634 32301 2668
rect 32301 2634 32335 2668
rect 32335 2634 32344 2668
rect 32292 2633 32344 2634
rect 32292 2596 32344 2621
rect 32292 2569 32301 2596
rect 32301 2569 32335 2596
rect 32335 2569 32344 2596
rect 32292 2524 32344 2557
rect 32292 2505 32301 2524
rect 32301 2505 32335 2524
rect 32335 2505 32344 2524
rect 32292 2490 32301 2493
rect 32301 2490 32335 2493
rect 32335 2490 32344 2493
rect 32292 2452 32344 2490
rect 32292 2441 32301 2452
rect 32301 2441 32335 2452
rect 32335 2441 32344 2452
rect 32292 2418 32301 2429
rect 32301 2418 32335 2429
rect 32335 2418 32344 2429
rect 32292 2380 32344 2418
rect 32292 2377 32301 2380
rect 32301 2377 32335 2380
rect 32335 2377 32344 2380
rect 32292 2346 32301 2365
rect 32301 2346 32335 2365
rect 32335 2346 32344 2365
rect 32292 2313 32344 2346
rect 32292 2274 32301 2301
rect 32301 2274 32335 2301
rect 32335 2274 32344 2301
rect 32292 2249 32344 2274
rect 32292 2236 32344 2237
rect 32292 2202 32301 2236
rect 32301 2202 32335 2236
rect 32335 2202 32344 2236
rect 32292 2185 32344 2202
rect 32292 2164 32344 2173
rect 32292 2130 32301 2164
rect 32301 2130 32335 2164
rect 32335 2130 32344 2164
rect 32292 2121 32344 2130
rect 32292 2092 32344 2109
rect 32292 2058 32301 2092
rect 32301 2058 32335 2092
rect 32335 2058 32344 2092
rect 32292 2057 32344 2058
rect 32292 2020 32344 2045
rect 32292 1993 32301 2020
rect 32301 1993 32335 2020
rect 32335 1993 32344 2020
rect 32292 1948 32344 1981
rect 32292 1929 32301 1948
rect 32301 1929 32335 1948
rect 32335 1929 32344 1948
rect 32292 1914 32301 1917
rect 32301 1914 32335 1917
rect 32335 1914 32344 1917
rect 32292 1876 32344 1914
rect 32292 1865 32301 1876
rect 32301 1865 32335 1876
rect 32335 1865 32344 1876
rect 32292 1842 32301 1853
rect 32301 1842 32335 1853
rect 32335 1842 32344 1853
rect 32292 1804 32344 1842
rect 32292 1801 32301 1804
rect 32301 1801 32335 1804
rect 32335 1801 32344 1804
rect 32292 1770 32301 1789
rect 32301 1770 32335 1789
rect 32335 1770 32344 1789
rect 32292 1737 32344 1770
rect 32292 1698 32301 1725
rect 32301 1698 32335 1725
rect 32335 1698 32344 1725
rect 32292 1673 32344 1698
rect 32292 1660 32344 1661
rect 32292 1626 32301 1660
rect 32301 1626 32335 1660
rect 32335 1626 32344 1660
rect 32292 1609 32344 1626
rect 32292 1588 32344 1597
rect 32292 1554 32301 1588
rect 32301 1554 32335 1588
rect 32335 1554 32344 1588
rect 32292 1545 32344 1554
rect 32292 1516 32344 1533
rect 32292 1482 32301 1516
rect 32301 1482 32335 1516
rect 32335 1482 32344 1516
rect 32292 1481 32344 1482
rect 32292 1444 32344 1469
rect 32292 1417 32301 1444
rect 32301 1417 32335 1444
rect 32335 1417 32344 1444
rect 32292 1372 32344 1405
rect 32292 1353 32301 1372
rect 32301 1353 32335 1372
rect 32335 1353 32344 1372
rect 32292 1338 32301 1341
rect 32301 1338 32335 1341
rect 32335 1338 32344 1341
rect 32292 1300 32344 1338
rect 32292 1289 32301 1300
rect 32301 1289 32335 1300
rect 32335 1289 32344 1300
rect 32292 1266 32301 1277
rect 32301 1266 32335 1277
rect 32335 1266 32344 1277
rect 32292 1228 32344 1266
rect 32292 1225 32301 1228
rect 32301 1225 32335 1228
rect 32335 1225 32344 1228
rect 32292 1194 32301 1213
rect 32301 1194 32335 1213
rect 32335 1194 32344 1213
rect 32292 1161 32344 1194
rect 32388 3100 32440 3133
rect 32388 3081 32397 3100
rect 32397 3081 32431 3100
rect 32431 3081 32440 3100
rect 32388 3066 32397 3069
rect 32397 3066 32431 3069
rect 32431 3066 32440 3069
rect 32388 3028 32440 3066
rect 32388 3017 32397 3028
rect 32397 3017 32431 3028
rect 32431 3017 32440 3028
rect 32388 2994 32397 3005
rect 32397 2994 32431 3005
rect 32431 2994 32440 3005
rect 32388 2956 32440 2994
rect 32388 2953 32397 2956
rect 32397 2953 32431 2956
rect 32431 2953 32440 2956
rect 32388 2922 32397 2941
rect 32397 2922 32431 2941
rect 32431 2922 32440 2941
rect 32388 2889 32440 2922
rect 32388 2850 32397 2877
rect 32397 2850 32431 2877
rect 32431 2850 32440 2877
rect 32388 2825 32440 2850
rect 32388 2812 32440 2813
rect 32388 2778 32397 2812
rect 32397 2778 32431 2812
rect 32431 2778 32440 2812
rect 32388 2761 32440 2778
rect 32388 2740 32440 2749
rect 32388 2706 32397 2740
rect 32397 2706 32431 2740
rect 32431 2706 32440 2740
rect 32388 2697 32440 2706
rect 32388 2668 32440 2685
rect 32388 2634 32397 2668
rect 32397 2634 32431 2668
rect 32431 2634 32440 2668
rect 32388 2633 32440 2634
rect 32388 2596 32440 2621
rect 32388 2569 32397 2596
rect 32397 2569 32431 2596
rect 32431 2569 32440 2596
rect 32388 2524 32440 2557
rect 32388 2505 32397 2524
rect 32397 2505 32431 2524
rect 32431 2505 32440 2524
rect 32388 2490 32397 2493
rect 32397 2490 32431 2493
rect 32431 2490 32440 2493
rect 32388 2452 32440 2490
rect 32388 2441 32397 2452
rect 32397 2441 32431 2452
rect 32431 2441 32440 2452
rect 32388 2418 32397 2429
rect 32397 2418 32431 2429
rect 32431 2418 32440 2429
rect 32388 2380 32440 2418
rect 32388 2377 32397 2380
rect 32397 2377 32431 2380
rect 32431 2377 32440 2380
rect 32388 2346 32397 2365
rect 32397 2346 32431 2365
rect 32431 2346 32440 2365
rect 32388 2313 32440 2346
rect 32388 2274 32397 2301
rect 32397 2274 32431 2301
rect 32431 2274 32440 2301
rect 32388 2249 32440 2274
rect 32388 2236 32440 2237
rect 32388 2202 32397 2236
rect 32397 2202 32431 2236
rect 32431 2202 32440 2236
rect 32388 2185 32440 2202
rect 32388 2164 32440 2173
rect 32388 2130 32397 2164
rect 32397 2130 32431 2164
rect 32431 2130 32440 2164
rect 32388 2121 32440 2130
rect 32388 2092 32440 2109
rect 32388 2058 32397 2092
rect 32397 2058 32431 2092
rect 32431 2058 32440 2092
rect 32388 2057 32440 2058
rect 32388 2020 32440 2045
rect 32388 1993 32397 2020
rect 32397 1993 32431 2020
rect 32431 1993 32440 2020
rect 32388 1948 32440 1981
rect 32388 1929 32397 1948
rect 32397 1929 32431 1948
rect 32431 1929 32440 1948
rect 32388 1914 32397 1917
rect 32397 1914 32431 1917
rect 32431 1914 32440 1917
rect 32388 1876 32440 1914
rect 32388 1865 32397 1876
rect 32397 1865 32431 1876
rect 32431 1865 32440 1876
rect 32388 1842 32397 1853
rect 32397 1842 32431 1853
rect 32431 1842 32440 1853
rect 32388 1804 32440 1842
rect 32388 1801 32397 1804
rect 32397 1801 32431 1804
rect 32431 1801 32440 1804
rect 32388 1770 32397 1789
rect 32397 1770 32431 1789
rect 32431 1770 32440 1789
rect 32388 1737 32440 1770
rect 32388 1698 32397 1725
rect 32397 1698 32431 1725
rect 32431 1698 32440 1725
rect 32388 1673 32440 1698
rect 32388 1660 32440 1661
rect 32388 1626 32397 1660
rect 32397 1626 32431 1660
rect 32431 1626 32440 1660
rect 32388 1609 32440 1626
rect 32388 1588 32440 1597
rect 32388 1554 32397 1588
rect 32397 1554 32431 1588
rect 32431 1554 32440 1588
rect 32388 1545 32440 1554
rect 32388 1516 32440 1533
rect 32388 1482 32397 1516
rect 32397 1482 32431 1516
rect 32431 1482 32440 1516
rect 32388 1481 32440 1482
rect 32388 1444 32440 1469
rect 32388 1417 32397 1444
rect 32397 1417 32431 1444
rect 32431 1417 32440 1444
rect 32388 1372 32440 1405
rect 32388 1353 32397 1372
rect 32397 1353 32431 1372
rect 32431 1353 32440 1372
rect 32388 1338 32397 1341
rect 32397 1338 32431 1341
rect 32431 1338 32440 1341
rect 32388 1300 32440 1338
rect 32388 1289 32397 1300
rect 32397 1289 32431 1300
rect 32431 1289 32440 1300
rect 32388 1266 32397 1277
rect 32397 1266 32431 1277
rect 32431 1266 32440 1277
rect 32388 1228 32440 1266
rect 32388 1225 32397 1228
rect 32397 1225 32431 1228
rect 32431 1225 32440 1228
rect 32388 1194 32397 1213
rect 32397 1194 32431 1213
rect 32431 1194 32440 1213
rect 32388 1161 32440 1194
rect 32484 3100 32536 3133
rect 32484 3081 32493 3100
rect 32493 3081 32527 3100
rect 32527 3081 32536 3100
rect 32484 3066 32493 3069
rect 32493 3066 32527 3069
rect 32527 3066 32536 3069
rect 32484 3028 32536 3066
rect 32484 3017 32493 3028
rect 32493 3017 32527 3028
rect 32527 3017 32536 3028
rect 32484 2994 32493 3005
rect 32493 2994 32527 3005
rect 32527 2994 32536 3005
rect 32484 2956 32536 2994
rect 32484 2953 32493 2956
rect 32493 2953 32527 2956
rect 32527 2953 32536 2956
rect 32484 2922 32493 2941
rect 32493 2922 32527 2941
rect 32527 2922 32536 2941
rect 32484 2889 32536 2922
rect 32484 2850 32493 2877
rect 32493 2850 32527 2877
rect 32527 2850 32536 2877
rect 32484 2825 32536 2850
rect 32484 2812 32536 2813
rect 32484 2778 32493 2812
rect 32493 2778 32527 2812
rect 32527 2778 32536 2812
rect 32484 2761 32536 2778
rect 32484 2740 32536 2749
rect 32484 2706 32493 2740
rect 32493 2706 32527 2740
rect 32527 2706 32536 2740
rect 32484 2697 32536 2706
rect 32484 2668 32536 2685
rect 32484 2634 32493 2668
rect 32493 2634 32527 2668
rect 32527 2634 32536 2668
rect 32484 2633 32536 2634
rect 32484 2596 32536 2621
rect 32484 2569 32493 2596
rect 32493 2569 32527 2596
rect 32527 2569 32536 2596
rect 32484 2524 32536 2557
rect 32484 2505 32493 2524
rect 32493 2505 32527 2524
rect 32527 2505 32536 2524
rect 32484 2490 32493 2493
rect 32493 2490 32527 2493
rect 32527 2490 32536 2493
rect 32484 2452 32536 2490
rect 32484 2441 32493 2452
rect 32493 2441 32527 2452
rect 32527 2441 32536 2452
rect 32484 2418 32493 2429
rect 32493 2418 32527 2429
rect 32527 2418 32536 2429
rect 32484 2380 32536 2418
rect 32484 2377 32493 2380
rect 32493 2377 32527 2380
rect 32527 2377 32536 2380
rect 32484 2346 32493 2365
rect 32493 2346 32527 2365
rect 32527 2346 32536 2365
rect 32484 2313 32536 2346
rect 32484 2274 32493 2301
rect 32493 2274 32527 2301
rect 32527 2274 32536 2301
rect 32484 2249 32536 2274
rect 32484 2236 32536 2237
rect 32484 2202 32493 2236
rect 32493 2202 32527 2236
rect 32527 2202 32536 2236
rect 32484 2185 32536 2202
rect 32484 2164 32536 2173
rect 32484 2130 32493 2164
rect 32493 2130 32527 2164
rect 32527 2130 32536 2164
rect 32484 2121 32536 2130
rect 32484 2092 32536 2109
rect 32484 2058 32493 2092
rect 32493 2058 32527 2092
rect 32527 2058 32536 2092
rect 32484 2057 32536 2058
rect 32484 2020 32536 2045
rect 32484 1993 32493 2020
rect 32493 1993 32527 2020
rect 32527 1993 32536 2020
rect 32484 1948 32536 1981
rect 32484 1929 32493 1948
rect 32493 1929 32527 1948
rect 32527 1929 32536 1948
rect 32484 1914 32493 1917
rect 32493 1914 32527 1917
rect 32527 1914 32536 1917
rect 32484 1876 32536 1914
rect 32484 1865 32493 1876
rect 32493 1865 32527 1876
rect 32527 1865 32536 1876
rect 32484 1842 32493 1853
rect 32493 1842 32527 1853
rect 32527 1842 32536 1853
rect 32484 1804 32536 1842
rect 32484 1801 32493 1804
rect 32493 1801 32527 1804
rect 32527 1801 32536 1804
rect 32484 1770 32493 1789
rect 32493 1770 32527 1789
rect 32527 1770 32536 1789
rect 32484 1737 32536 1770
rect 32484 1698 32493 1725
rect 32493 1698 32527 1725
rect 32527 1698 32536 1725
rect 32484 1673 32536 1698
rect 32484 1660 32536 1661
rect 32484 1626 32493 1660
rect 32493 1626 32527 1660
rect 32527 1626 32536 1660
rect 32484 1609 32536 1626
rect 32484 1588 32536 1597
rect 32484 1554 32493 1588
rect 32493 1554 32527 1588
rect 32527 1554 32536 1588
rect 32484 1545 32536 1554
rect 32484 1516 32536 1533
rect 32484 1482 32493 1516
rect 32493 1482 32527 1516
rect 32527 1482 32536 1516
rect 32484 1481 32536 1482
rect 32484 1444 32536 1469
rect 32484 1417 32493 1444
rect 32493 1417 32527 1444
rect 32527 1417 32536 1444
rect 32484 1372 32536 1405
rect 32484 1353 32493 1372
rect 32493 1353 32527 1372
rect 32527 1353 32536 1372
rect 32484 1338 32493 1341
rect 32493 1338 32527 1341
rect 32527 1338 32536 1341
rect 32484 1300 32536 1338
rect 32484 1289 32493 1300
rect 32493 1289 32527 1300
rect 32527 1289 32536 1300
rect 32484 1266 32493 1277
rect 32493 1266 32527 1277
rect 32527 1266 32536 1277
rect 32484 1228 32536 1266
rect 32484 1225 32493 1228
rect 32493 1225 32527 1228
rect 32527 1225 32536 1228
rect 32484 1194 32493 1213
rect 32493 1194 32527 1213
rect 32527 1194 32536 1213
rect 32484 1161 32536 1194
rect 32580 3100 32632 3133
rect 32580 3081 32589 3100
rect 32589 3081 32623 3100
rect 32623 3081 32632 3100
rect 32580 3066 32589 3069
rect 32589 3066 32623 3069
rect 32623 3066 32632 3069
rect 32580 3028 32632 3066
rect 32580 3017 32589 3028
rect 32589 3017 32623 3028
rect 32623 3017 32632 3028
rect 32580 2994 32589 3005
rect 32589 2994 32623 3005
rect 32623 2994 32632 3005
rect 32580 2956 32632 2994
rect 32580 2953 32589 2956
rect 32589 2953 32623 2956
rect 32623 2953 32632 2956
rect 32580 2922 32589 2941
rect 32589 2922 32623 2941
rect 32623 2922 32632 2941
rect 32580 2889 32632 2922
rect 32580 2850 32589 2877
rect 32589 2850 32623 2877
rect 32623 2850 32632 2877
rect 32580 2825 32632 2850
rect 32580 2812 32632 2813
rect 32580 2778 32589 2812
rect 32589 2778 32623 2812
rect 32623 2778 32632 2812
rect 32580 2761 32632 2778
rect 32580 2740 32632 2749
rect 32580 2706 32589 2740
rect 32589 2706 32623 2740
rect 32623 2706 32632 2740
rect 32580 2697 32632 2706
rect 32580 2668 32632 2685
rect 32580 2634 32589 2668
rect 32589 2634 32623 2668
rect 32623 2634 32632 2668
rect 32580 2633 32632 2634
rect 32580 2596 32632 2621
rect 32580 2569 32589 2596
rect 32589 2569 32623 2596
rect 32623 2569 32632 2596
rect 32580 2524 32632 2557
rect 32580 2505 32589 2524
rect 32589 2505 32623 2524
rect 32623 2505 32632 2524
rect 32580 2490 32589 2493
rect 32589 2490 32623 2493
rect 32623 2490 32632 2493
rect 32580 2452 32632 2490
rect 32580 2441 32589 2452
rect 32589 2441 32623 2452
rect 32623 2441 32632 2452
rect 32580 2418 32589 2429
rect 32589 2418 32623 2429
rect 32623 2418 32632 2429
rect 32580 2380 32632 2418
rect 32580 2377 32589 2380
rect 32589 2377 32623 2380
rect 32623 2377 32632 2380
rect 32580 2346 32589 2365
rect 32589 2346 32623 2365
rect 32623 2346 32632 2365
rect 32580 2313 32632 2346
rect 32580 2274 32589 2301
rect 32589 2274 32623 2301
rect 32623 2274 32632 2301
rect 32580 2249 32632 2274
rect 32580 2236 32632 2237
rect 32580 2202 32589 2236
rect 32589 2202 32623 2236
rect 32623 2202 32632 2236
rect 32580 2185 32632 2202
rect 32580 2164 32632 2173
rect 32580 2130 32589 2164
rect 32589 2130 32623 2164
rect 32623 2130 32632 2164
rect 32580 2121 32632 2130
rect 32580 2092 32632 2109
rect 32580 2058 32589 2092
rect 32589 2058 32623 2092
rect 32623 2058 32632 2092
rect 32580 2057 32632 2058
rect 32580 2020 32632 2045
rect 32580 1993 32589 2020
rect 32589 1993 32623 2020
rect 32623 1993 32632 2020
rect 32580 1948 32632 1981
rect 32580 1929 32589 1948
rect 32589 1929 32623 1948
rect 32623 1929 32632 1948
rect 32580 1914 32589 1917
rect 32589 1914 32623 1917
rect 32623 1914 32632 1917
rect 32580 1876 32632 1914
rect 32580 1865 32589 1876
rect 32589 1865 32623 1876
rect 32623 1865 32632 1876
rect 32580 1842 32589 1853
rect 32589 1842 32623 1853
rect 32623 1842 32632 1853
rect 32580 1804 32632 1842
rect 32580 1801 32589 1804
rect 32589 1801 32623 1804
rect 32623 1801 32632 1804
rect 32580 1770 32589 1789
rect 32589 1770 32623 1789
rect 32623 1770 32632 1789
rect 32580 1737 32632 1770
rect 32580 1698 32589 1725
rect 32589 1698 32623 1725
rect 32623 1698 32632 1725
rect 32580 1673 32632 1698
rect 32580 1660 32632 1661
rect 32580 1626 32589 1660
rect 32589 1626 32623 1660
rect 32623 1626 32632 1660
rect 32580 1609 32632 1626
rect 32580 1588 32632 1597
rect 32580 1554 32589 1588
rect 32589 1554 32623 1588
rect 32623 1554 32632 1588
rect 32580 1545 32632 1554
rect 32580 1516 32632 1533
rect 32580 1482 32589 1516
rect 32589 1482 32623 1516
rect 32623 1482 32632 1516
rect 32580 1481 32632 1482
rect 32580 1444 32632 1469
rect 32580 1417 32589 1444
rect 32589 1417 32623 1444
rect 32623 1417 32632 1444
rect 32580 1372 32632 1405
rect 32580 1353 32589 1372
rect 32589 1353 32623 1372
rect 32623 1353 32632 1372
rect 32580 1338 32589 1341
rect 32589 1338 32623 1341
rect 32623 1338 32632 1341
rect 32580 1300 32632 1338
rect 32580 1289 32589 1300
rect 32589 1289 32623 1300
rect 32623 1289 32632 1300
rect 32580 1266 32589 1277
rect 32589 1266 32623 1277
rect 32623 1266 32632 1277
rect 32580 1228 32632 1266
rect 32580 1225 32589 1228
rect 32589 1225 32623 1228
rect 32623 1225 32632 1228
rect 32580 1194 32589 1213
rect 32589 1194 32623 1213
rect 32623 1194 32632 1213
rect 32580 1161 32632 1194
rect 32676 3100 32728 3133
rect 32676 3081 32685 3100
rect 32685 3081 32719 3100
rect 32719 3081 32728 3100
rect 32676 3066 32685 3069
rect 32685 3066 32719 3069
rect 32719 3066 32728 3069
rect 32676 3028 32728 3066
rect 32676 3017 32685 3028
rect 32685 3017 32719 3028
rect 32719 3017 32728 3028
rect 32676 2994 32685 3005
rect 32685 2994 32719 3005
rect 32719 2994 32728 3005
rect 32676 2956 32728 2994
rect 32676 2953 32685 2956
rect 32685 2953 32719 2956
rect 32719 2953 32728 2956
rect 32676 2922 32685 2941
rect 32685 2922 32719 2941
rect 32719 2922 32728 2941
rect 32676 2889 32728 2922
rect 32676 2850 32685 2877
rect 32685 2850 32719 2877
rect 32719 2850 32728 2877
rect 32676 2825 32728 2850
rect 32676 2812 32728 2813
rect 32676 2778 32685 2812
rect 32685 2778 32719 2812
rect 32719 2778 32728 2812
rect 32676 2761 32728 2778
rect 32676 2740 32728 2749
rect 32676 2706 32685 2740
rect 32685 2706 32719 2740
rect 32719 2706 32728 2740
rect 32676 2697 32728 2706
rect 32676 2668 32728 2685
rect 32676 2634 32685 2668
rect 32685 2634 32719 2668
rect 32719 2634 32728 2668
rect 32676 2633 32728 2634
rect 32676 2596 32728 2621
rect 32676 2569 32685 2596
rect 32685 2569 32719 2596
rect 32719 2569 32728 2596
rect 32676 2524 32728 2557
rect 32676 2505 32685 2524
rect 32685 2505 32719 2524
rect 32719 2505 32728 2524
rect 32676 2490 32685 2493
rect 32685 2490 32719 2493
rect 32719 2490 32728 2493
rect 32676 2452 32728 2490
rect 32676 2441 32685 2452
rect 32685 2441 32719 2452
rect 32719 2441 32728 2452
rect 32676 2418 32685 2429
rect 32685 2418 32719 2429
rect 32719 2418 32728 2429
rect 32676 2380 32728 2418
rect 32676 2377 32685 2380
rect 32685 2377 32719 2380
rect 32719 2377 32728 2380
rect 32676 2346 32685 2365
rect 32685 2346 32719 2365
rect 32719 2346 32728 2365
rect 32676 2313 32728 2346
rect 32676 2274 32685 2301
rect 32685 2274 32719 2301
rect 32719 2274 32728 2301
rect 32676 2249 32728 2274
rect 32676 2236 32728 2237
rect 32676 2202 32685 2236
rect 32685 2202 32719 2236
rect 32719 2202 32728 2236
rect 32676 2185 32728 2202
rect 32676 2164 32728 2173
rect 32676 2130 32685 2164
rect 32685 2130 32719 2164
rect 32719 2130 32728 2164
rect 32676 2121 32728 2130
rect 32676 2092 32728 2109
rect 32676 2058 32685 2092
rect 32685 2058 32719 2092
rect 32719 2058 32728 2092
rect 32676 2057 32728 2058
rect 32676 2020 32728 2045
rect 32676 1993 32685 2020
rect 32685 1993 32719 2020
rect 32719 1993 32728 2020
rect 32676 1948 32728 1981
rect 32676 1929 32685 1948
rect 32685 1929 32719 1948
rect 32719 1929 32728 1948
rect 32676 1914 32685 1917
rect 32685 1914 32719 1917
rect 32719 1914 32728 1917
rect 32676 1876 32728 1914
rect 32676 1865 32685 1876
rect 32685 1865 32719 1876
rect 32719 1865 32728 1876
rect 32676 1842 32685 1853
rect 32685 1842 32719 1853
rect 32719 1842 32728 1853
rect 32676 1804 32728 1842
rect 32676 1801 32685 1804
rect 32685 1801 32719 1804
rect 32719 1801 32728 1804
rect 32676 1770 32685 1789
rect 32685 1770 32719 1789
rect 32719 1770 32728 1789
rect 32676 1737 32728 1770
rect 32676 1698 32685 1725
rect 32685 1698 32719 1725
rect 32719 1698 32728 1725
rect 32676 1673 32728 1698
rect 32676 1660 32728 1661
rect 32676 1626 32685 1660
rect 32685 1626 32719 1660
rect 32719 1626 32728 1660
rect 32676 1609 32728 1626
rect 32676 1588 32728 1597
rect 32676 1554 32685 1588
rect 32685 1554 32719 1588
rect 32719 1554 32728 1588
rect 32676 1545 32728 1554
rect 32676 1516 32728 1533
rect 32676 1482 32685 1516
rect 32685 1482 32719 1516
rect 32719 1482 32728 1516
rect 32676 1481 32728 1482
rect 32676 1444 32728 1469
rect 32676 1417 32685 1444
rect 32685 1417 32719 1444
rect 32719 1417 32728 1444
rect 32676 1372 32728 1405
rect 32676 1353 32685 1372
rect 32685 1353 32719 1372
rect 32719 1353 32728 1372
rect 32676 1338 32685 1341
rect 32685 1338 32719 1341
rect 32719 1338 32728 1341
rect 32676 1300 32728 1338
rect 32676 1289 32685 1300
rect 32685 1289 32719 1300
rect 32719 1289 32728 1300
rect 32676 1266 32685 1277
rect 32685 1266 32719 1277
rect 32719 1266 32728 1277
rect 32676 1228 32728 1266
rect 32676 1225 32685 1228
rect 32685 1225 32719 1228
rect 32719 1225 32728 1228
rect 32676 1194 32685 1213
rect 32685 1194 32719 1213
rect 32719 1194 32728 1213
rect 32676 1161 32728 1194
rect 32772 3100 32824 3133
rect 32772 3081 32781 3100
rect 32781 3081 32815 3100
rect 32815 3081 32824 3100
rect 32772 3066 32781 3069
rect 32781 3066 32815 3069
rect 32815 3066 32824 3069
rect 32772 3028 32824 3066
rect 32772 3017 32781 3028
rect 32781 3017 32815 3028
rect 32815 3017 32824 3028
rect 32772 2994 32781 3005
rect 32781 2994 32815 3005
rect 32815 2994 32824 3005
rect 32772 2956 32824 2994
rect 32772 2953 32781 2956
rect 32781 2953 32815 2956
rect 32815 2953 32824 2956
rect 32772 2922 32781 2941
rect 32781 2922 32815 2941
rect 32815 2922 32824 2941
rect 32772 2889 32824 2922
rect 32772 2850 32781 2877
rect 32781 2850 32815 2877
rect 32815 2850 32824 2877
rect 32772 2825 32824 2850
rect 32772 2812 32824 2813
rect 32772 2778 32781 2812
rect 32781 2778 32815 2812
rect 32815 2778 32824 2812
rect 32772 2761 32824 2778
rect 32772 2740 32824 2749
rect 32772 2706 32781 2740
rect 32781 2706 32815 2740
rect 32815 2706 32824 2740
rect 32772 2697 32824 2706
rect 32772 2668 32824 2685
rect 32772 2634 32781 2668
rect 32781 2634 32815 2668
rect 32815 2634 32824 2668
rect 32772 2633 32824 2634
rect 32772 2596 32824 2621
rect 32772 2569 32781 2596
rect 32781 2569 32815 2596
rect 32815 2569 32824 2596
rect 32772 2524 32824 2557
rect 32772 2505 32781 2524
rect 32781 2505 32815 2524
rect 32815 2505 32824 2524
rect 32772 2490 32781 2493
rect 32781 2490 32815 2493
rect 32815 2490 32824 2493
rect 32772 2452 32824 2490
rect 32772 2441 32781 2452
rect 32781 2441 32815 2452
rect 32815 2441 32824 2452
rect 32772 2418 32781 2429
rect 32781 2418 32815 2429
rect 32815 2418 32824 2429
rect 32772 2380 32824 2418
rect 32772 2377 32781 2380
rect 32781 2377 32815 2380
rect 32815 2377 32824 2380
rect 32772 2346 32781 2365
rect 32781 2346 32815 2365
rect 32815 2346 32824 2365
rect 32772 2313 32824 2346
rect 32772 2274 32781 2301
rect 32781 2274 32815 2301
rect 32815 2274 32824 2301
rect 32772 2249 32824 2274
rect 32772 2236 32824 2237
rect 32772 2202 32781 2236
rect 32781 2202 32815 2236
rect 32815 2202 32824 2236
rect 32772 2185 32824 2202
rect 32772 2164 32824 2173
rect 32772 2130 32781 2164
rect 32781 2130 32815 2164
rect 32815 2130 32824 2164
rect 32772 2121 32824 2130
rect 32772 2092 32824 2109
rect 32772 2058 32781 2092
rect 32781 2058 32815 2092
rect 32815 2058 32824 2092
rect 32772 2057 32824 2058
rect 32772 2020 32824 2045
rect 32772 1993 32781 2020
rect 32781 1993 32815 2020
rect 32815 1993 32824 2020
rect 32772 1948 32824 1981
rect 32772 1929 32781 1948
rect 32781 1929 32815 1948
rect 32815 1929 32824 1948
rect 32772 1914 32781 1917
rect 32781 1914 32815 1917
rect 32815 1914 32824 1917
rect 32772 1876 32824 1914
rect 32772 1865 32781 1876
rect 32781 1865 32815 1876
rect 32815 1865 32824 1876
rect 32772 1842 32781 1853
rect 32781 1842 32815 1853
rect 32815 1842 32824 1853
rect 32772 1804 32824 1842
rect 32772 1801 32781 1804
rect 32781 1801 32815 1804
rect 32815 1801 32824 1804
rect 32772 1770 32781 1789
rect 32781 1770 32815 1789
rect 32815 1770 32824 1789
rect 32772 1737 32824 1770
rect 32772 1698 32781 1725
rect 32781 1698 32815 1725
rect 32815 1698 32824 1725
rect 32772 1673 32824 1698
rect 32772 1660 32824 1661
rect 32772 1626 32781 1660
rect 32781 1626 32815 1660
rect 32815 1626 32824 1660
rect 32772 1609 32824 1626
rect 32772 1588 32824 1597
rect 32772 1554 32781 1588
rect 32781 1554 32815 1588
rect 32815 1554 32824 1588
rect 32772 1545 32824 1554
rect 32772 1516 32824 1533
rect 32772 1482 32781 1516
rect 32781 1482 32815 1516
rect 32815 1482 32824 1516
rect 32772 1481 32824 1482
rect 32772 1444 32824 1469
rect 32772 1417 32781 1444
rect 32781 1417 32815 1444
rect 32815 1417 32824 1444
rect 32772 1372 32824 1405
rect 32772 1353 32781 1372
rect 32781 1353 32815 1372
rect 32815 1353 32824 1372
rect 32772 1338 32781 1341
rect 32781 1338 32815 1341
rect 32815 1338 32824 1341
rect 32772 1300 32824 1338
rect 32772 1289 32781 1300
rect 32781 1289 32815 1300
rect 32815 1289 32824 1300
rect 32772 1266 32781 1277
rect 32781 1266 32815 1277
rect 32815 1266 32824 1277
rect 32772 1228 32824 1266
rect 32772 1225 32781 1228
rect 32781 1225 32815 1228
rect 32815 1225 32824 1228
rect 32772 1194 32781 1213
rect 32781 1194 32815 1213
rect 32815 1194 32824 1213
rect 32772 1161 32824 1194
rect 32868 3100 32920 3133
rect 32868 3081 32877 3100
rect 32877 3081 32911 3100
rect 32911 3081 32920 3100
rect 32868 3066 32877 3069
rect 32877 3066 32911 3069
rect 32911 3066 32920 3069
rect 32868 3028 32920 3066
rect 32868 3017 32877 3028
rect 32877 3017 32911 3028
rect 32911 3017 32920 3028
rect 32868 2994 32877 3005
rect 32877 2994 32911 3005
rect 32911 2994 32920 3005
rect 32868 2956 32920 2994
rect 32868 2953 32877 2956
rect 32877 2953 32911 2956
rect 32911 2953 32920 2956
rect 32868 2922 32877 2941
rect 32877 2922 32911 2941
rect 32911 2922 32920 2941
rect 32868 2889 32920 2922
rect 32868 2850 32877 2877
rect 32877 2850 32911 2877
rect 32911 2850 32920 2877
rect 32868 2825 32920 2850
rect 32868 2812 32920 2813
rect 32868 2778 32877 2812
rect 32877 2778 32911 2812
rect 32911 2778 32920 2812
rect 32868 2761 32920 2778
rect 32868 2740 32920 2749
rect 32868 2706 32877 2740
rect 32877 2706 32911 2740
rect 32911 2706 32920 2740
rect 32868 2697 32920 2706
rect 32868 2668 32920 2685
rect 32868 2634 32877 2668
rect 32877 2634 32911 2668
rect 32911 2634 32920 2668
rect 32868 2633 32920 2634
rect 32868 2596 32920 2621
rect 32868 2569 32877 2596
rect 32877 2569 32911 2596
rect 32911 2569 32920 2596
rect 32868 2524 32920 2557
rect 32868 2505 32877 2524
rect 32877 2505 32911 2524
rect 32911 2505 32920 2524
rect 32868 2490 32877 2493
rect 32877 2490 32911 2493
rect 32911 2490 32920 2493
rect 32868 2452 32920 2490
rect 32868 2441 32877 2452
rect 32877 2441 32911 2452
rect 32911 2441 32920 2452
rect 32868 2418 32877 2429
rect 32877 2418 32911 2429
rect 32911 2418 32920 2429
rect 32868 2380 32920 2418
rect 32868 2377 32877 2380
rect 32877 2377 32911 2380
rect 32911 2377 32920 2380
rect 32868 2346 32877 2365
rect 32877 2346 32911 2365
rect 32911 2346 32920 2365
rect 32868 2313 32920 2346
rect 32868 2274 32877 2301
rect 32877 2274 32911 2301
rect 32911 2274 32920 2301
rect 32868 2249 32920 2274
rect 32868 2236 32920 2237
rect 32868 2202 32877 2236
rect 32877 2202 32911 2236
rect 32911 2202 32920 2236
rect 32868 2185 32920 2202
rect 32868 2164 32920 2173
rect 32868 2130 32877 2164
rect 32877 2130 32911 2164
rect 32911 2130 32920 2164
rect 32868 2121 32920 2130
rect 32868 2092 32920 2109
rect 32868 2058 32877 2092
rect 32877 2058 32911 2092
rect 32911 2058 32920 2092
rect 32868 2057 32920 2058
rect 32868 2020 32920 2045
rect 32868 1993 32877 2020
rect 32877 1993 32911 2020
rect 32911 1993 32920 2020
rect 32868 1948 32920 1981
rect 32868 1929 32877 1948
rect 32877 1929 32911 1948
rect 32911 1929 32920 1948
rect 32868 1914 32877 1917
rect 32877 1914 32911 1917
rect 32911 1914 32920 1917
rect 32868 1876 32920 1914
rect 32868 1865 32877 1876
rect 32877 1865 32911 1876
rect 32911 1865 32920 1876
rect 32868 1842 32877 1853
rect 32877 1842 32911 1853
rect 32911 1842 32920 1853
rect 32868 1804 32920 1842
rect 32868 1801 32877 1804
rect 32877 1801 32911 1804
rect 32911 1801 32920 1804
rect 32868 1770 32877 1789
rect 32877 1770 32911 1789
rect 32911 1770 32920 1789
rect 32868 1737 32920 1770
rect 32868 1698 32877 1725
rect 32877 1698 32911 1725
rect 32911 1698 32920 1725
rect 32868 1673 32920 1698
rect 32868 1660 32920 1661
rect 32868 1626 32877 1660
rect 32877 1626 32911 1660
rect 32911 1626 32920 1660
rect 32868 1609 32920 1626
rect 32868 1588 32920 1597
rect 32868 1554 32877 1588
rect 32877 1554 32911 1588
rect 32911 1554 32920 1588
rect 32868 1545 32920 1554
rect 32868 1516 32920 1533
rect 32868 1482 32877 1516
rect 32877 1482 32911 1516
rect 32911 1482 32920 1516
rect 32868 1481 32920 1482
rect 32868 1444 32920 1469
rect 32868 1417 32877 1444
rect 32877 1417 32911 1444
rect 32911 1417 32920 1444
rect 32868 1372 32920 1405
rect 32868 1353 32877 1372
rect 32877 1353 32911 1372
rect 32911 1353 32920 1372
rect 32868 1338 32877 1341
rect 32877 1338 32911 1341
rect 32911 1338 32920 1341
rect 32868 1300 32920 1338
rect 32868 1289 32877 1300
rect 32877 1289 32911 1300
rect 32911 1289 32920 1300
rect 32868 1266 32877 1277
rect 32877 1266 32911 1277
rect 32911 1266 32920 1277
rect 32868 1228 32920 1266
rect 32868 1225 32877 1228
rect 32877 1225 32911 1228
rect 32911 1225 32920 1228
rect 32868 1194 32877 1213
rect 32877 1194 32911 1213
rect 32911 1194 32920 1213
rect 32868 1161 32920 1194
rect 32964 3100 33016 3133
rect 32964 3081 32973 3100
rect 32973 3081 33007 3100
rect 33007 3081 33016 3100
rect 32964 3066 32973 3069
rect 32973 3066 33007 3069
rect 33007 3066 33016 3069
rect 32964 3028 33016 3066
rect 32964 3017 32973 3028
rect 32973 3017 33007 3028
rect 33007 3017 33016 3028
rect 32964 2994 32973 3005
rect 32973 2994 33007 3005
rect 33007 2994 33016 3005
rect 32964 2956 33016 2994
rect 32964 2953 32973 2956
rect 32973 2953 33007 2956
rect 33007 2953 33016 2956
rect 32964 2922 32973 2941
rect 32973 2922 33007 2941
rect 33007 2922 33016 2941
rect 32964 2889 33016 2922
rect 32964 2850 32973 2877
rect 32973 2850 33007 2877
rect 33007 2850 33016 2877
rect 32964 2825 33016 2850
rect 32964 2812 33016 2813
rect 32964 2778 32973 2812
rect 32973 2778 33007 2812
rect 33007 2778 33016 2812
rect 32964 2761 33016 2778
rect 32964 2740 33016 2749
rect 32964 2706 32973 2740
rect 32973 2706 33007 2740
rect 33007 2706 33016 2740
rect 32964 2697 33016 2706
rect 32964 2668 33016 2685
rect 32964 2634 32973 2668
rect 32973 2634 33007 2668
rect 33007 2634 33016 2668
rect 32964 2633 33016 2634
rect 32964 2596 33016 2621
rect 32964 2569 32973 2596
rect 32973 2569 33007 2596
rect 33007 2569 33016 2596
rect 32964 2524 33016 2557
rect 32964 2505 32973 2524
rect 32973 2505 33007 2524
rect 33007 2505 33016 2524
rect 32964 2490 32973 2493
rect 32973 2490 33007 2493
rect 33007 2490 33016 2493
rect 32964 2452 33016 2490
rect 32964 2441 32973 2452
rect 32973 2441 33007 2452
rect 33007 2441 33016 2452
rect 32964 2418 32973 2429
rect 32973 2418 33007 2429
rect 33007 2418 33016 2429
rect 32964 2380 33016 2418
rect 32964 2377 32973 2380
rect 32973 2377 33007 2380
rect 33007 2377 33016 2380
rect 32964 2346 32973 2365
rect 32973 2346 33007 2365
rect 33007 2346 33016 2365
rect 32964 2313 33016 2346
rect 32964 2274 32973 2301
rect 32973 2274 33007 2301
rect 33007 2274 33016 2301
rect 32964 2249 33016 2274
rect 32964 2236 33016 2237
rect 32964 2202 32973 2236
rect 32973 2202 33007 2236
rect 33007 2202 33016 2236
rect 32964 2185 33016 2202
rect 32964 2164 33016 2173
rect 32964 2130 32973 2164
rect 32973 2130 33007 2164
rect 33007 2130 33016 2164
rect 32964 2121 33016 2130
rect 32964 2092 33016 2109
rect 32964 2058 32973 2092
rect 32973 2058 33007 2092
rect 33007 2058 33016 2092
rect 32964 2057 33016 2058
rect 32964 2020 33016 2045
rect 32964 1993 32973 2020
rect 32973 1993 33007 2020
rect 33007 1993 33016 2020
rect 32964 1948 33016 1981
rect 32964 1929 32973 1948
rect 32973 1929 33007 1948
rect 33007 1929 33016 1948
rect 32964 1914 32973 1917
rect 32973 1914 33007 1917
rect 33007 1914 33016 1917
rect 32964 1876 33016 1914
rect 32964 1865 32973 1876
rect 32973 1865 33007 1876
rect 33007 1865 33016 1876
rect 32964 1842 32973 1853
rect 32973 1842 33007 1853
rect 33007 1842 33016 1853
rect 32964 1804 33016 1842
rect 32964 1801 32973 1804
rect 32973 1801 33007 1804
rect 33007 1801 33016 1804
rect 32964 1770 32973 1789
rect 32973 1770 33007 1789
rect 33007 1770 33016 1789
rect 32964 1737 33016 1770
rect 32964 1698 32973 1725
rect 32973 1698 33007 1725
rect 33007 1698 33016 1725
rect 32964 1673 33016 1698
rect 32964 1660 33016 1661
rect 32964 1626 32973 1660
rect 32973 1626 33007 1660
rect 33007 1626 33016 1660
rect 32964 1609 33016 1626
rect 32964 1588 33016 1597
rect 32964 1554 32973 1588
rect 32973 1554 33007 1588
rect 33007 1554 33016 1588
rect 32964 1545 33016 1554
rect 32964 1516 33016 1533
rect 32964 1482 32973 1516
rect 32973 1482 33007 1516
rect 33007 1482 33016 1516
rect 32964 1481 33016 1482
rect 32964 1444 33016 1469
rect 32964 1417 32973 1444
rect 32973 1417 33007 1444
rect 33007 1417 33016 1444
rect 32964 1372 33016 1405
rect 32964 1353 32973 1372
rect 32973 1353 33007 1372
rect 33007 1353 33016 1372
rect 32964 1338 32973 1341
rect 32973 1338 33007 1341
rect 33007 1338 33016 1341
rect 32964 1300 33016 1338
rect 32964 1289 32973 1300
rect 32973 1289 33007 1300
rect 33007 1289 33016 1300
rect 32964 1266 32973 1277
rect 32973 1266 33007 1277
rect 33007 1266 33016 1277
rect 32964 1228 33016 1266
rect 32964 1225 32973 1228
rect 32973 1225 33007 1228
rect 33007 1225 33016 1228
rect 32964 1194 32973 1213
rect 32973 1194 33007 1213
rect 33007 1194 33016 1213
rect 32964 1161 33016 1194
rect 33060 3100 33112 3133
rect 33060 3081 33069 3100
rect 33069 3081 33103 3100
rect 33103 3081 33112 3100
rect 33060 3066 33069 3069
rect 33069 3066 33103 3069
rect 33103 3066 33112 3069
rect 33060 3028 33112 3066
rect 33060 3017 33069 3028
rect 33069 3017 33103 3028
rect 33103 3017 33112 3028
rect 33060 2994 33069 3005
rect 33069 2994 33103 3005
rect 33103 2994 33112 3005
rect 33060 2956 33112 2994
rect 33060 2953 33069 2956
rect 33069 2953 33103 2956
rect 33103 2953 33112 2956
rect 33060 2922 33069 2941
rect 33069 2922 33103 2941
rect 33103 2922 33112 2941
rect 33060 2889 33112 2922
rect 33060 2850 33069 2877
rect 33069 2850 33103 2877
rect 33103 2850 33112 2877
rect 33060 2825 33112 2850
rect 33060 2812 33112 2813
rect 33060 2778 33069 2812
rect 33069 2778 33103 2812
rect 33103 2778 33112 2812
rect 33060 2761 33112 2778
rect 33060 2740 33112 2749
rect 33060 2706 33069 2740
rect 33069 2706 33103 2740
rect 33103 2706 33112 2740
rect 33060 2697 33112 2706
rect 33060 2668 33112 2685
rect 33060 2634 33069 2668
rect 33069 2634 33103 2668
rect 33103 2634 33112 2668
rect 33060 2633 33112 2634
rect 33060 2596 33112 2621
rect 33060 2569 33069 2596
rect 33069 2569 33103 2596
rect 33103 2569 33112 2596
rect 33060 2524 33112 2557
rect 33060 2505 33069 2524
rect 33069 2505 33103 2524
rect 33103 2505 33112 2524
rect 33060 2490 33069 2493
rect 33069 2490 33103 2493
rect 33103 2490 33112 2493
rect 33060 2452 33112 2490
rect 33060 2441 33069 2452
rect 33069 2441 33103 2452
rect 33103 2441 33112 2452
rect 33060 2418 33069 2429
rect 33069 2418 33103 2429
rect 33103 2418 33112 2429
rect 33060 2380 33112 2418
rect 33060 2377 33069 2380
rect 33069 2377 33103 2380
rect 33103 2377 33112 2380
rect 33060 2346 33069 2365
rect 33069 2346 33103 2365
rect 33103 2346 33112 2365
rect 33060 2313 33112 2346
rect 33060 2274 33069 2301
rect 33069 2274 33103 2301
rect 33103 2274 33112 2301
rect 33060 2249 33112 2274
rect 33060 2236 33112 2237
rect 33060 2202 33069 2236
rect 33069 2202 33103 2236
rect 33103 2202 33112 2236
rect 33060 2185 33112 2202
rect 33060 2164 33112 2173
rect 33060 2130 33069 2164
rect 33069 2130 33103 2164
rect 33103 2130 33112 2164
rect 33060 2121 33112 2130
rect 33060 2092 33112 2109
rect 33060 2058 33069 2092
rect 33069 2058 33103 2092
rect 33103 2058 33112 2092
rect 33060 2057 33112 2058
rect 33060 2020 33112 2045
rect 33060 1993 33069 2020
rect 33069 1993 33103 2020
rect 33103 1993 33112 2020
rect 33060 1948 33112 1981
rect 33060 1929 33069 1948
rect 33069 1929 33103 1948
rect 33103 1929 33112 1948
rect 33060 1914 33069 1917
rect 33069 1914 33103 1917
rect 33103 1914 33112 1917
rect 33060 1876 33112 1914
rect 33060 1865 33069 1876
rect 33069 1865 33103 1876
rect 33103 1865 33112 1876
rect 33060 1842 33069 1853
rect 33069 1842 33103 1853
rect 33103 1842 33112 1853
rect 33060 1804 33112 1842
rect 33060 1801 33069 1804
rect 33069 1801 33103 1804
rect 33103 1801 33112 1804
rect 33060 1770 33069 1789
rect 33069 1770 33103 1789
rect 33103 1770 33112 1789
rect 33060 1737 33112 1770
rect 33060 1698 33069 1725
rect 33069 1698 33103 1725
rect 33103 1698 33112 1725
rect 33060 1673 33112 1698
rect 33060 1660 33112 1661
rect 33060 1626 33069 1660
rect 33069 1626 33103 1660
rect 33103 1626 33112 1660
rect 33060 1609 33112 1626
rect 33060 1588 33112 1597
rect 33060 1554 33069 1588
rect 33069 1554 33103 1588
rect 33103 1554 33112 1588
rect 33060 1545 33112 1554
rect 33060 1516 33112 1533
rect 33060 1482 33069 1516
rect 33069 1482 33103 1516
rect 33103 1482 33112 1516
rect 33060 1481 33112 1482
rect 33060 1444 33112 1469
rect 33060 1417 33069 1444
rect 33069 1417 33103 1444
rect 33103 1417 33112 1444
rect 33060 1372 33112 1405
rect 33060 1353 33069 1372
rect 33069 1353 33103 1372
rect 33103 1353 33112 1372
rect 33060 1338 33069 1341
rect 33069 1338 33103 1341
rect 33103 1338 33112 1341
rect 33060 1300 33112 1338
rect 33060 1289 33069 1300
rect 33069 1289 33103 1300
rect 33103 1289 33112 1300
rect 33060 1266 33069 1277
rect 33069 1266 33103 1277
rect 33103 1266 33112 1277
rect 33060 1228 33112 1266
rect 33060 1225 33069 1228
rect 33069 1225 33103 1228
rect 33103 1225 33112 1228
rect 33060 1194 33069 1213
rect 33069 1194 33103 1213
rect 33103 1194 33112 1213
rect 33060 1161 33112 1194
rect 33156 3100 33208 3133
rect 33156 3081 33165 3100
rect 33165 3081 33199 3100
rect 33199 3081 33208 3100
rect 33156 3066 33165 3069
rect 33165 3066 33199 3069
rect 33199 3066 33208 3069
rect 33156 3028 33208 3066
rect 33156 3017 33165 3028
rect 33165 3017 33199 3028
rect 33199 3017 33208 3028
rect 33156 2994 33165 3005
rect 33165 2994 33199 3005
rect 33199 2994 33208 3005
rect 33156 2956 33208 2994
rect 33156 2953 33165 2956
rect 33165 2953 33199 2956
rect 33199 2953 33208 2956
rect 33156 2922 33165 2941
rect 33165 2922 33199 2941
rect 33199 2922 33208 2941
rect 33156 2889 33208 2922
rect 33156 2850 33165 2877
rect 33165 2850 33199 2877
rect 33199 2850 33208 2877
rect 33156 2825 33208 2850
rect 33156 2812 33208 2813
rect 33156 2778 33165 2812
rect 33165 2778 33199 2812
rect 33199 2778 33208 2812
rect 33156 2761 33208 2778
rect 33156 2740 33208 2749
rect 33156 2706 33165 2740
rect 33165 2706 33199 2740
rect 33199 2706 33208 2740
rect 33156 2697 33208 2706
rect 33156 2668 33208 2685
rect 33156 2634 33165 2668
rect 33165 2634 33199 2668
rect 33199 2634 33208 2668
rect 33156 2633 33208 2634
rect 33156 2596 33208 2621
rect 33156 2569 33165 2596
rect 33165 2569 33199 2596
rect 33199 2569 33208 2596
rect 33156 2524 33208 2557
rect 33156 2505 33165 2524
rect 33165 2505 33199 2524
rect 33199 2505 33208 2524
rect 33156 2490 33165 2493
rect 33165 2490 33199 2493
rect 33199 2490 33208 2493
rect 33156 2452 33208 2490
rect 33156 2441 33165 2452
rect 33165 2441 33199 2452
rect 33199 2441 33208 2452
rect 33156 2418 33165 2429
rect 33165 2418 33199 2429
rect 33199 2418 33208 2429
rect 33156 2380 33208 2418
rect 33156 2377 33165 2380
rect 33165 2377 33199 2380
rect 33199 2377 33208 2380
rect 33156 2346 33165 2365
rect 33165 2346 33199 2365
rect 33199 2346 33208 2365
rect 33156 2313 33208 2346
rect 33156 2274 33165 2301
rect 33165 2274 33199 2301
rect 33199 2274 33208 2301
rect 33156 2249 33208 2274
rect 33156 2236 33208 2237
rect 33156 2202 33165 2236
rect 33165 2202 33199 2236
rect 33199 2202 33208 2236
rect 33156 2185 33208 2202
rect 33156 2164 33208 2173
rect 33156 2130 33165 2164
rect 33165 2130 33199 2164
rect 33199 2130 33208 2164
rect 33156 2121 33208 2130
rect 33156 2092 33208 2109
rect 33156 2058 33165 2092
rect 33165 2058 33199 2092
rect 33199 2058 33208 2092
rect 33156 2057 33208 2058
rect 33156 2020 33208 2045
rect 33156 1993 33165 2020
rect 33165 1993 33199 2020
rect 33199 1993 33208 2020
rect 33156 1948 33208 1981
rect 33156 1929 33165 1948
rect 33165 1929 33199 1948
rect 33199 1929 33208 1948
rect 33156 1914 33165 1917
rect 33165 1914 33199 1917
rect 33199 1914 33208 1917
rect 33156 1876 33208 1914
rect 33156 1865 33165 1876
rect 33165 1865 33199 1876
rect 33199 1865 33208 1876
rect 33156 1842 33165 1853
rect 33165 1842 33199 1853
rect 33199 1842 33208 1853
rect 33156 1804 33208 1842
rect 33156 1801 33165 1804
rect 33165 1801 33199 1804
rect 33199 1801 33208 1804
rect 33156 1770 33165 1789
rect 33165 1770 33199 1789
rect 33199 1770 33208 1789
rect 33156 1737 33208 1770
rect 33156 1698 33165 1725
rect 33165 1698 33199 1725
rect 33199 1698 33208 1725
rect 33156 1673 33208 1698
rect 33156 1660 33208 1661
rect 33156 1626 33165 1660
rect 33165 1626 33199 1660
rect 33199 1626 33208 1660
rect 33156 1609 33208 1626
rect 33156 1588 33208 1597
rect 33156 1554 33165 1588
rect 33165 1554 33199 1588
rect 33199 1554 33208 1588
rect 33156 1545 33208 1554
rect 33156 1516 33208 1533
rect 33156 1482 33165 1516
rect 33165 1482 33199 1516
rect 33199 1482 33208 1516
rect 33156 1481 33208 1482
rect 33156 1444 33208 1469
rect 33156 1417 33165 1444
rect 33165 1417 33199 1444
rect 33199 1417 33208 1444
rect 33156 1372 33208 1405
rect 33156 1353 33165 1372
rect 33165 1353 33199 1372
rect 33199 1353 33208 1372
rect 33156 1338 33165 1341
rect 33165 1338 33199 1341
rect 33199 1338 33208 1341
rect 33156 1300 33208 1338
rect 33156 1289 33165 1300
rect 33165 1289 33199 1300
rect 33199 1289 33208 1300
rect 33156 1266 33165 1277
rect 33165 1266 33199 1277
rect 33199 1266 33208 1277
rect 33156 1228 33208 1266
rect 33156 1225 33165 1228
rect 33165 1225 33199 1228
rect 33199 1225 33208 1228
rect 33156 1194 33165 1213
rect 33165 1194 33199 1213
rect 33199 1194 33208 1213
rect 33156 1161 33208 1194
rect 33252 3100 33304 3133
rect 33252 3081 33261 3100
rect 33261 3081 33295 3100
rect 33295 3081 33304 3100
rect 33252 3066 33261 3069
rect 33261 3066 33295 3069
rect 33295 3066 33304 3069
rect 33252 3028 33304 3066
rect 33252 3017 33261 3028
rect 33261 3017 33295 3028
rect 33295 3017 33304 3028
rect 33252 2994 33261 3005
rect 33261 2994 33295 3005
rect 33295 2994 33304 3005
rect 33252 2956 33304 2994
rect 33252 2953 33261 2956
rect 33261 2953 33295 2956
rect 33295 2953 33304 2956
rect 33252 2922 33261 2941
rect 33261 2922 33295 2941
rect 33295 2922 33304 2941
rect 33252 2889 33304 2922
rect 33252 2850 33261 2877
rect 33261 2850 33295 2877
rect 33295 2850 33304 2877
rect 33252 2825 33304 2850
rect 33252 2812 33304 2813
rect 33252 2778 33261 2812
rect 33261 2778 33295 2812
rect 33295 2778 33304 2812
rect 33252 2761 33304 2778
rect 33252 2740 33304 2749
rect 33252 2706 33261 2740
rect 33261 2706 33295 2740
rect 33295 2706 33304 2740
rect 33252 2697 33304 2706
rect 33252 2668 33304 2685
rect 33252 2634 33261 2668
rect 33261 2634 33295 2668
rect 33295 2634 33304 2668
rect 33252 2633 33304 2634
rect 33252 2596 33304 2621
rect 33252 2569 33261 2596
rect 33261 2569 33295 2596
rect 33295 2569 33304 2596
rect 33252 2524 33304 2557
rect 33252 2505 33261 2524
rect 33261 2505 33295 2524
rect 33295 2505 33304 2524
rect 33252 2490 33261 2493
rect 33261 2490 33295 2493
rect 33295 2490 33304 2493
rect 33252 2452 33304 2490
rect 33252 2441 33261 2452
rect 33261 2441 33295 2452
rect 33295 2441 33304 2452
rect 33252 2418 33261 2429
rect 33261 2418 33295 2429
rect 33295 2418 33304 2429
rect 33252 2380 33304 2418
rect 33252 2377 33261 2380
rect 33261 2377 33295 2380
rect 33295 2377 33304 2380
rect 33252 2346 33261 2365
rect 33261 2346 33295 2365
rect 33295 2346 33304 2365
rect 33252 2313 33304 2346
rect 33252 2274 33261 2301
rect 33261 2274 33295 2301
rect 33295 2274 33304 2301
rect 33252 2249 33304 2274
rect 33252 2236 33304 2237
rect 33252 2202 33261 2236
rect 33261 2202 33295 2236
rect 33295 2202 33304 2236
rect 33252 2185 33304 2202
rect 33252 2164 33304 2173
rect 33252 2130 33261 2164
rect 33261 2130 33295 2164
rect 33295 2130 33304 2164
rect 33252 2121 33304 2130
rect 33252 2092 33304 2109
rect 33252 2058 33261 2092
rect 33261 2058 33295 2092
rect 33295 2058 33304 2092
rect 33252 2057 33304 2058
rect 33252 2020 33304 2045
rect 33252 1993 33261 2020
rect 33261 1993 33295 2020
rect 33295 1993 33304 2020
rect 33252 1948 33304 1981
rect 33252 1929 33261 1948
rect 33261 1929 33295 1948
rect 33295 1929 33304 1948
rect 33252 1914 33261 1917
rect 33261 1914 33295 1917
rect 33295 1914 33304 1917
rect 33252 1876 33304 1914
rect 33252 1865 33261 1876
rect 33261 1865 33295 1876
rect 33295 1865 33304 1876
rect 33252 1842 33261 1853
rect 33261 1842 33295 1853
rect 33295 1842 33304 1853
rect 33252 1804 33304 1842
rect 33252 1801 33261 1804
rect 33261 1801 33295 1804
rect 33295 1801 33304 1804
rect 33252 1770 33261 1789
rect 33261 1770 33295 1789
rect 33295 1770 33304 1789
rect 33252 1737 33304 1770
rect 33252 1698 33261 1725
rect 33261 1698 33295 1725
rect 33295 1698 33304 1725
rect 33252 1673 33304 1698
rect 33252 1660 33304 1661
rect 33252 1626 33261 1660
rect 33261 1626 33295 1660
rect 33295 1626 33304 1660
rect 33252 1609 33304 1626
rect 33252 1588 33304 1597
rect 33252 1554 33261 1588
rect 33261 1554 33295 1588
rect 33295 1554 33304 1588
rect 33252 1545 33304 1554
rect 33252 1516 33304 1533
rect 33252 1482 33261 1516
rect 33261 1482 33295 1516
rect 33295 1482 33304 1516
rect 33252 1481 33304 1482
rect 33252 1444 33304 1469
rect 33252 1417 33261 1444
rect 33261 1417 33295 1444
rect 33295 1417 33304 1444
rect 33252 1372 33304 1405
rect 33252 1353 33261 1372
rect 33261 1353 33295 1372
rect 33295 1353 33304 1372
rect 33252 1338 33261 1341
rect 33261 1338 33295 1341
rect 33295 1338 33304 1341
rect 33252 1300 33304 1338
rect 33252 1289 33261 1300
rect 33261 1289 33295 1300
rect 33295 1289 33304 1300
rect 33252 1266 33261 1277
rect 33261 1266 33295 1277
rect 33295 1266 33304 1277
rect 33252 1228 33304 1266
rect 33252 1225 33261 1228
rect 33261 1225 33295 1228
rect 33295 1225 33304 1228
rect 33252 1194 33261 1213
rect 33261 1194 33295 1213
rect 33295 1194 33304 1213
rect 33252 1161 33304 1194
rect 33348 3100 33400 3133
rect 33348 3081 33357 3100
rect 33357 3081 33391 3100
rect 33391 3081 33400 3100
rect 33348 3066 33357 3069
rect 33357 3066 33391 3069
rect 33391 3066 33400 3069
rect 33348 3028 33400 3066
rect 33348 3017 33357 3028
rect 33357 3017 33391 3028
rect 33391 3017 33400 3028
rect 33348 2994 33357 3005
rect 33357 2994 33391 3005
rect 33391 2994 33400 3005
rect 33348 2956 33400 2994
rect 33348 2953 33357 2956
rect 33357 2953 33391 2956
rect 33391 2953 33400 2956
rect 33348 2922 33357 2941
rect 33357 2922 33391 2941
rect 33391 2922 33400 2941
rect 33348 2889 33400 2922
rect 33348 2850 33357 2877
rect 33357 2850 33391 2877
rect 33391 2850 33400 2877
rect 33348 2825 33400 2850
rect 33348 2812 33400 2813
rect 33348 2778 33357 2812
rect 33357 2778 33391 2812
rect 33391 2778 33400 2812
rect 33348 2761 33400 2778
rect 33348 2740 33400 2749
rect 33348 2706 33357 2740
rect 33357 2706 33391 2740
rect 33391 2706 33400 2740
rect 33348 2697 33400 2706
rect 33348 2668 33400 2685
rect 33348 2634 33357 2668
rect 33357 2634 33391 2668
rect 33391 2634 33400 2668
rect 33348 2633 33400 2634
rect 33348 2596 33400 2621
rect 33348 2569 33357 2596
rect 33357 2569 33391 2596
rect 33391 2569 33400 2596
rect 33348 2524 33400 2557
rect 33348 2505 33357 2524
rect 33357 2505 33391 2524
rect 33391 2505 33400 2524
rect 33348 2490 33357 2493
rect 33357 2490 33391 2493
rect 33391 2490 33400 2493
rect 33348 2452 33400 2490
rect 33348 2441 33357 2452
rect 33357 2441 33391 2452
rect 33391 2441 33400 2452
rect 33348 2418 33357 2429
rect 33357 2418 33391 2429
rect 33391 2418 33400 2429
rect 33348 2380 33400 2418
rect 33348 2377 33357 2380
rect 33357 2377 33391 2380
rect 33391 2377 33400 2380
rect 33348 2346 33357 2365
rect 33357 2346 33391 2365
rect 33391 2346 33400 2365
rect 33348 2313 33400 2346
rect 33348 2274 33357 2301
rect 33357 2274 33391 2301
rect 33391 2274 33400 2301
rect 33348 2249 33400 2274
rect 33348 2236 33400 2237
rect 33348 2202 33357 2236
rect 33357 2202 33391 2236
rect 33391 2202 33400 2236
rect 33348 2185 33400 2202
rect 33348 2164 33400 2173
rect 33348 2130 33357 2164
rect 33357 2130 33391 2164
rect 33391 2130 33400 2164
rect 33348 2121 33400 2130
rect 33348 2092 33400 2109
rect 33348 2058 33357 2092
rect 33357 2058 33391 2092
rect 33391 2058 33400 2092
rect 33348 2057 33400 2058
rect 33348 2020 33400 2045
rect 33348 1993 33357 2020
rect 33357 1993 33391 2020
rect 33391 1993 33400 2020
rect 33348 1948 33400 1981
rect 33348 1929 33357 1948
rect 33357 1929 33391 1948
rect 33391 1929 33400 1948
rect 33348 1914 33357 1917
rect 33357 1914 33391 1917
rect 33391 1914 33400 1917
rect 33348 1876 33400 1914
rect 33348 1865 33357 1876
rect 33357 1865 33391 1876
rect 33391 1865 33400 1876
rect 33348 1842 33357 1853
rect 33357 1842 33391 1853
rect 33391 1842 33400 1853
rect 33348 1804 33400 1842
rect 33348 1801 33357 1804
rect 33357 1801 33391 1804
rect 33391 1801 33400 1804
rect 33348 1770 33357 1789
rect 33357 1770 33391 1789
rect 33391 1770 33400 1789
rect 33348 1737 33400 1770
rect 33348 1698 33357 1725
rect 33357 1698 33391 1725
rect 33391 1698 33400 1725
rect 33348 1673 33400 1698
rect 33348 1660 33400 1661
rect 33348 1626 33357 1660
rect 33357 1626 33391 1660
rect 33391 1626 33400 1660
rect 33348 1609 33400 1626
rect 33348 1588 33400 1597
rect 33348 1554 33357 1588
rect 33357 1554 33391 1588
rect 33391 1554 33400 1588
rect 33348 1545 33400 1554
rect 33348 1516 33400 1533
rect 33348 1482 33357 1516
rect 33357 1482 33391 1516
rect 33391 1482 33400 1516
rect 33348 1481 33400 1482
rect 33348 1444 33400 1469
rect 33348 1417 33357 1444
rect 33357 1417 33391 1444
rect 33391 1417 33400 1444
rect 33348 1372 33400 1405
rect 33348 1353 33357 1372
rect 33357 1353 33391 1372
rect 33391 1353 33400 1372
rect 33348 1338 33357 1341
rect 33357 1338 33391 1341
rect 33391 1338 33400 1341
rect 33348 1300 33400 1338
rect 33348 1289 33357 1300
rect 33357 1289 33391 1300
rect 33391 1289 33400 1300
rect 33348 1266 33357 1277
rect 33357 1266 33391 1277
rect 33391 1266 33400 1277
rect 33348 1228 33400 1266
rect 33348 1225 33357 1228
rect 33357 1225 33391 1228
rect 33391 1225 33400 1228
rect 33348 1194 33357 1213
rect 33357 1194 33391 1213
rect 33391 1194 33400 1213
rect 33348 1161 33400 1194
rect 33444 3100 33496 3133
rect 33444 3081 33453 3100
rect 33453 3081 33487 3100
rect 33487 3081 33496 3100
rect 33444 3066 33453 3069
rect 33453 3066 33487 3069
rect 33487 3066 33496 3069
rect 33444 3028 33496 3066
rect 33444 3017 33453 3028
rect 33453 3017 33487 3028
rect 33487 3017 33496 3028
rect 33444 2994 33453 3005
rect 33453 2994 33487 3005
rect 33487 2994 33496 3005
rect 33444 2956 33496 2994
rect 33444 2953 33453 2956
rect 33453 2953 33487 2956
rect 33487 2953 33496 2956
rect 33444 2922 33453 2941
rect 33453 2922 33487 2941
rect 33487 2922 33496 2941
rect 33444 2889 33496 2922
rect 33444 2850 33453 2877
rect 33453 2850 33487 2877
rect 33487 2850 33496 2877
rect 33444 2825 33496 2850
rect 33444 2812 33496 2813
rect 33444 2778 33453 2812
rect 33453 2778 33487 2812
rect 33487 2778 33496 2812
rect 33444 2761 33496 2778
rect 33444 2740 33496 2749
rect 33444 2706 33453 2740
rect 33453 2706 33487 2740
rect 33487 2706 33496 2740
rect 33444 2697 33496 2706
rect 33444 2668 33496 2685
rect 33444 2634 33453 2668
rect 33453 2634 33487 2668
rect 33487 2634 33496 2668
rect 33444 2633 33496 2634
rect 33444 2596 33496 2621
rect 33444 2569 33453 2596
rect 33453 2569 33487 2596
rect 33487 2569 33496 2596
rect 33444 2524 33496 2557
rect 33444 2505 33453 2524
rect 33453 2505 33487 2524
rect 33487 2505 33496 2524
rect 33444 2490 33453 2493
rect 33453 2490 33487 2493
rect 33487 2490 33496 2493
rect 33444 2452 33496 2490
rect 33444 2441 33453 2452
rect 33453 2441 33487 2452
rect 33487 2441 33496 2452
rect 33444 2418 33453 2429
rect 33453 2418 33487 2429
rect 33487 2418 33496 2429
rect 33444 2380 33496 2418
rect 33444 2377 33453 2380
rect 33453 2377 33487 2380
rect 33487 2377 33496 2380
rect 33444 2346 33453 2365
rect 33453 2346 33487 2365
rect 33487 2346 33496 2365
rect 33444 2313 33496 2346
rect 33444 2274 33453 2301
rect 33453 2274 33487 2301
rect 33487 2274 33496 2301
rect 33444 2249 33496 2274
rect 33444 2236 33496 2237
rect 33444 2202 33453 2236
rect 33453 2202 33487 2236
rect 33487 2202 33496 2236
rect 33444 2185 33496 2202
rect 33444 2164 33496 2173
rect 33444 2130 33453 2164
rect 33453 2130 33487 2164
rect 33487 2130 33496 2164
rect 33444 2121 33496 2130
rect 33444 2092 33496 2109
rect 33444 2058 33453 2092
rect 33453 2058 33487 2092
rect 33487 2058 33496 2092
rect 33444 2057 33496 2058
rect 33444 2020 33496 2045
rect 33444 1993 33453 2020
rect 33453 1993 33487 2020
rect 33487 1993 33496 2020
rect 33444 1948 33496 1981
rect 33444 1929 33453 1948
rect 33453 1929 33487 1948
rect 33487 1929 33496 1948
rect 33444 1914 33453 1917
rect 33453 1914 33487 1917
rect 33487 1914 33496 1917
rect 33444 1876 33496 1914
rect 33444 1865 33453 1876
rect 33453 1865 33487 1876
rect 33487 1865 33496 1876
rect 33444 1842 33453 1853
rect 33453 1842 33487 1853
rect 33487 1842 33496 1853
rect 33444 1804 33496 1842
rect 33444 1801 33453 1804
rect 33453 1801 33487 1804
rect 33487 1801 33496 1804
rect 33444 1770 33453 1789
rect 33453 1770 33487 1789
rect 33487 1770 33496 1789
rect 33444 1737 33496 1770
rect 33444 1698 33453 1725
rect 33453 1698 33487 1725
rect 33487 1698 33496 1725
rect 33444 1673 33496 1698
rect 33444 1660 33496 1661
rect 33444 1626 33453 1660
rect 33453 1626 33487 1660
rect 33487 1626 33496 1660
rect 33444 1609 33496 1626
rect 33444 1588 33496 1597
rect 33444 1554 33453 1588
rect 33453 1554 33487 1588
rect 33487 1554 33496 1588
rect 33444 1545 33496 1554
rect 33444 1516 33496 1533
rect 33444 1482 33453 1516
rect 33453 1482 33487 1516
rect 33487 1482 33496 1516
rect 33444 1481 33496 1482
rect 33444 1444 33496 1469
rect 33444 1417 33453 1444
rect 33453 1417 33487 1444
rect 33487 1417 33496 1444
rect 33444 1372 33496 1405
rect 33444 1353 33453 1372
rect 33453 1353 33487 1372
rect 33487 1353 33496 1372
rect 33444 1338 33453 1341
rect 33453 1338 33487 1341
rect 33487 1338 33496 1341
rect 33444 1300 33496 1338
rect 33444 1289 33453 1300
rect 33453 1289 33487 1300
rect 33487 1289 33496 1300
rect 33444 1266 33453 1277
rect 33453 1266 33487 1277
rect 33487 1266 33496 1277
rect 33444 1228 33496 1266
rect 33444 1225 33453 1228
rect 33453 1225 33487 1228
rect 33487 1225 33496 1228
rect 33444 1194 33453 1213
rect 33453 1194 33487 1213
rect 33487 1194 33496 1213
rect 33444 1161 33496 1194
rect 33540 3100 33592 3133
rect 33540 3081 33549 3100
rect 33549 3081 33583 3100
rect 33583 3081 33592 3100
rect 33540 3066 33549 3069
rect 33549 3066 33583 3069
rect 33583 3066 33592 3069
rect 33540 3028 33592 3066
rect 33540 3017 33549 3028
rect 33549 3017 33583 3028
rect 33583 3017 33592 3028
rect 33540 2994 33549 3005
rect 33549 2994 33583 3005
rect 33583 2994 33592 3005
rect 33540 2956 33592 2994
rect 33540 2953 33549 2956
rect 33549 2953 33583 2956
rect 33583 2953 33592 2956
rect 33540 2922 33549 2941
rect 33549 2922 33583 2941
rect 33583 2922 33592 2941
rect 33540 2889 33592 2922
rect 33540 2850 33549 2877
rect 33549 2850 33583 2877
rect 33583 2850 33592 2877
rect 33540 2825 33592 2850
rect 33540 2812 33592 2813
rect 33540 2778 33549 2812
rect 33549 2778 33583 2812
rect 33583 2778 33592 2812
rect 33540 2761 33592 2778
rect 33540 2740 33592 2749
rect 33540 2706 33549 2740
rect 33549 2706 33583 2740
rect 33583 2706 33592 2740
rect 33540 2697 33592 2706
rect 33540 2668 33592 2685
rect 33540 2634 33549 2668
rect 33549 2634 33583 2668
rect 33583 2634 33592 2668
rect 33540 2633 33592 2634
rect 33540 2596 33592 2621
rect 33540 2569 33549 2596
rect 33549 2569 33583 2596
rect 33583 2569 33592 2596
rect 33540 2524 33592 2557
rect 33540 2505 33549 2524
rect 33549 2505 33583 2524
rect 33583 2505 33592 2524
rect 33540 2490 33549 2493
rect 33549 2490 33583 2493
rect 33583 2490 33592 2493
rect 33540 2452 33592 2490
rect 33540 2441 33549 2452
rect 33549 2441 33583 2452
rect 33583 2441 33592 2452
rect 33540 2418 33549 2429
rect 33549 2418 33583 2429
rect 33583 2418 33592 2429
rect 33540 2380 33592 2418
rect 33540 2377 33549 2380
rect 33549 2377 33583 2380
rect 33583 2377 33592 2380
rect 33540 2346 33549 2365
rect 33549 2346 33583 2365
rect 33583 2346 33592 2365
rect 33540 2313 33592 2346
rect 33540 2274 33549 2301
rect 33549 2274 33583 2301
rect 33583 2274 33592 2301
rect 33540 2249 33592 2274
rect 33540 2236 33592 2237
rect 33540 2202 33549 2236
rect 33549 2202 33583 2236
rect 33583 2202 33592 2236
rect 33540 2185 33592 2202
rect 33540 2164 33592 2173
rect 33540 2130 33549 2164
rect 33549 2130 33583 2164
rect 33583 2130 33592 2164
rect 33540 2121 33592 2130
rect 33540 2092 33592 2109
rect 33540 2058 33549 2092
rect 33549 2058 33583 2092
rect 33583 2058 33592 2092
rect 33540 2057 33592 2058
rect 33540 2020 33592 2045
rect 33540 1993 33549 2020
rect 33549 1993 33583 2020
rect 33583 1993 33592 2020
rect 33540 1948 33592 1981
rect 33540 1929 33549 1948
rect 33549 1929 33583 1948
rect 33583 1929 33592 1948
rect 33540 1914 33549 1917
rect 33549 1914 33583 1917
rect 33583 1914 33592 1917
rect 33540 1876 33592 1914
rect 33540 1865 33549 1876
rect 33549 1865 33583 1876
rect 33583 1865 33592 1876
rect 33540 1842 33549 1853
rect 33549 1842 33583 1853
rect 33583 1842 33592 1853
rect 33540 1804 33592 1842
rect 33540 1801 33549 1804
rect 33549 1801 33583 1804
rect 33583 1801 33592 1804
rect 33540 1770 33549 1789
rect 33549 1770 33583 1789
rect 33583 1770 33592 1789
rect 33540 1737 33592 1770
rect 33540 1698 33549 1725
rect 33549 1698 33583 1725
rect 33583 1698 33592 1725
rect 33540 1673 33592 1698
rect 33540 1660 33592 1661
rect 33540 1626 33549 1660
rect 33549 1626 33583 1660
rect 33583 1626 33592 1660
rect 33540 1609 33592 1626
rect 33540 1588 33592 1597
rect 33540 1554 33549 1588
rect 33549 1554 33583 1588
rect 33583 1554 33592 1588
rect 33540 1545 33592 1554
rect 33540 1516 33592 1533
rect 33540 1482 33549 1516
rect 33549 1482 33583 1516
rect 33583 1482 33592 1516
rect 33540 1481 33592 1482
rect 33540 1444 33592 1469
rect 33540 1417 33549 1444
rect 33549 1417 33583 1444
rect 33583 1417 33592 1444
rect 33540 1372 33592 1405
rect 33540 1353 33549 1372
rect 33549 1353 33583 1372
rect 33583 1353 33592 1372
rect 33540 1338 33549 1341
rect 33549 1338 33583 1341
rect 33583 1338 33592 1341
rect 33540 1300 33592 1338
rect 33540 1289 33549 1300
rect 33549 1289 33583 1300
rect 33583 1289 33592 1300
rect 33540 1266 33549 1277
rect 33549 1266 33583 1277
rect 33583 1266 33592 1277
rect 33540 1228 33592 1266
rect 33540 1225 33549 1228
rect 33549 1225 33583 1228
rect 33583 1225 33592 1228
rect 33540 1194 33549 1213
rect 33549 1194 33583 1213
rect 33583 1194 33592 1213
rect 33540 1161 33592 1194
rect 33636 3100 33688 3133
rect 33636 3081 33645 3100
rect 33645 3081 33679 3100
rect 33679 3081 33688 3100
rect 33636 3066 33645 3069
rect 33645 3066 33679 3069
rect 33679 3066 33688 3069
rect 33636 3028 33688 3066
rect 33636 3017 33645 3028
rect 33645 3017 33679 3028
rect 33679 3017 33688 3028
rect 33636 2994 33645 3005
rect 33645 2994 33679 3005
rect 33679 2994 33688 3005
rect 33636 2956 33688 2994
rect 33636 2953 33645 2956
rect 33645 2953 33679 2956
rect 33679 2953 33688 2956
rect 33636 2922 33645 2941
rect 33645 2922 33679 2941
rect 33679 2922 33688 2941
rect 33636 2889 33688 2922
rect 33636 2850 33645 2877
rect 33645 2850 33679 2877
rect 33679 2850 33688 2877
rect 33636 2825 33688 2850
rect 33636 2812 33688 2813
rect 33636 2778 33645 2812
rect 33645 2778 33679 2812
rect 33679 2778 33688 2812
rect 33636 2761 33688 2778
rect 33636 2740 33688 2749
rect 33636 2706 33645 2740
rect 33645 2706 33679 2740
rect 33679 2706 33688 2740
rect 33636 2697 33688 2706
rect 33636 2668 33688 2685
rect 33636 2634 33645 2668
rect 33645 2634 33679 2668
rect 33679 2634 33688 2668
rect 33636 2633 33688 2634
rect 33636 2596 33688 2621
rect 33636 2569 33645 2596
rect 33645 2569 33679 2596
rect 33679 2569 33688 2596
rect 33636 2524 33688 2557
rect 33636 2505 33645 2524
rect 33645 2505 33679 2524
rect 33679 2505 33688 2524
rect 33636 2490 33645 2493
rect 33645 2490 33679 2493
rect 33679 2490 33688 2493
rect 33636 2452 33688 2490
rect 33636 2441 33645 2452
rect 33645 2441 33679 2452
rect 33679 2441 33688 2452
rect 33636 2418 33645 2429
rect 33645 2418 33679 2429
rect 33679 2418 33688 2429
rect 33636 2380 33688 2418
rect 33636 2377 33645 2380
rect 33645 2377 33679 2380
rect 33679 2377 33688 2380
rect 33636 2346 33645 2365
rect 33645 2346 33679 2365
rect 33679 2346 33688 2365
rect 33636 2313 33688 2346
rect 33636 2274 33645 2301
rect 33645 2274 33679 2301
rect 33679 2274 33688 2301
rect 33636 2249 33688 2274
rect 33636 2236 33688 2237
rect 33636 2202 33645 2236
rect 33645 2202 33679 2236
rect 33679 2202 33688 2236
rect 33636 2185 33688 2202
rect 33636 2164 33688 2173
rect 33636 2130 33645 2164
rect 33645 2130 33679 2164
rect 33679 2130 33688 2164
rect 33636 2121 33688 2130
rect 33636 2092 33688 2109
rect 33636 2058 33645 2092
rect 33645 2058 33679 2092
rect 33679 2058 33688 2092
rect 33636 2057 33688 2058
rect 33636 2020 33688 2045
rect 33636 1993 33645 2020
rect 33645 1993 33679 2020
rect 33679 1993 33688 2020
rect 33636 1948 33688 1981
rect 33636 1929 33645 1948
rect 33645 1929 33679 1948
rect 33679 1929 33688 1948
rect 33636 1914 33645 1917
rect 33645 1914 33679 1917
rect 33679 1914 33688 1917
rect 33636 1876 33688 1914
rect 33636 1865 33645 1876
rect 33645 1865 33679 1876
rect 33679 1865 33688 1876
rect 33636 1842 33645 1853
rect 33645 1842 33679 1853
rect 33679 1842 33688 1853
rect 33636 1804 33688 1842
rect 33636 1801 33645 1804
rect 33645 1801 33679 1804
rect 33679 1801 33688 1804
rect 33636 1770 33645 1789
rect 33645 1770 33679 1789
rect 33679 1770 33688 1789
rect 33636 1737 33688 1770
rect 33636 1698 33645 1725
rect 33645 1698 33679 1725
rect 33679 1698 33688 1725
rect 33636 1673 33688 1698
rect 33636 1660 33688 1661
rect 33636 1626 33645 1660
rect 33645 1626 33679 1660
rect 33679 1626 33688 1660
rect 33636 1609 33688 1626
rect 33636 1588 33688 1597
rect 33636 1554 33645 1588
rect 33645 1554 33679 1588
rect 33679 1554 33688 1588
rect 33636 1545 33688 1554
rect 33636 1516 33688 1533
rect 33636 1482 33645 1516
rect 33645 1482 33679 1516
rect 33679 1482 33688 1516
rect 33636 1481 33688 1482
rect 33636 1444 33688 1469
rect 33636 1417 33645 1444
rect 33645 1417 33679 1444
rect 33679 1417 33688 1444
rect 33636 1372 33688 1405
rect 33636 1353 33645 1372
rect 33645 1353 33679 1372
rect 33679 1353 33688 1372
rect 33636 1338 33645 1341
rect 33645 1338 33679 1341
rect 33679 1338 33688 1341
rect 33636 1300 33688 1338
rect 33636 1289 33645 1300
rect 33645 1289 33679 1300
rect 33679 1289 33688 1300
rect 33636 1266 33645 1277
rect 33645 1266 33679 1277
rect 33679 1266 33688 1277
rect 33636 1228 33688 1266
rect 33636 1225 33645 1228
rect 33645 1225 33679 1228
rect 33679 1225 33688 1228
rect 33636 1194 33645 1213
rect 33645 1194 33679 1213
rect 33679 1194 33688 1213
rect 33636 1161 33688 1194
rect 33732 3100 33784 3133
rect 33732 3081 33741 3100
rect 33741 3081 33775 3100
rect 33775 3081 33784 3100
rect 33732 3066 33741 3069
rect 33741 3066 33775 3069
rect 33775 3066 33784 3069
rect 33732 3028 33784 3066
rect 33732 3017 33741 3028
rect 33741 3017 33775 3028
rect 33775 3017 33784 3028
rect 33732 2994 33741 3005
rect 33741 2994 33775 3005
rect 33775 2994 33784 3005
rect 33732 2956 33784 2994
rect 33732 2953 33741 2956
rect 33741 2953 33775 2956
rect 33775 2953 33784 2956
rect 33732 2922 33741 2941
rect 33741 2922 33775 2941
rect 33775 2922 33784 2941
rect 33732 2889 33784 2922
rect 33732 2850 33741 2877
rect 33741 2850 33775 2877
rect 33775 2850 33784 2877
rect 33732 2825 33784 2850
rect 33732 2812 33784 2813
rect 33732 2778 33741 2812
rect 33741 2778 33775 2812
rect 33775 2778 33784 2812
rect 33732 2761 33784 2778
rect 33732 2740 33784 2749
rect 33732 2706 33741 2740
rect 33741 2706 33775 2740
rect 33775 2706 33784 2740
rect 33732 2697 33784 2706
rect 33732 2668 33784 2685
rect 33732 2634 33741 2668
rect 33741 2634 33775 2668
rect 33775 2634 33784 2668
rect 33732 2633 33784 2634
rect 33732 2596 33784 2621
rect 33732 2569 33741 2596
rect 33741 2569 33775 2596
rect 33775 2569 33784 2596
rect 33732 2524 33784 2557
rect 33732 2505 33741 2524
rect 33741 2505 33775 2524
rect 33775 2505 33784 2524
rect 33732 2490 33741 2493
rect 33741 2490 33775 2493
rect 33775 2490 33784 2493
rect 33732 2452 33784 2490
rect 33732 2441 33741 2452
rect 33741 2441 33775 2452
rect 33775 2441 33784 2452
rect 33732 2418 33741 2429
rect 33741 2418 33775 2429
rect 33775 2418 33784 2429
rect 33732 2380 33784 2418
rect 33732 2377 33741 2380
rect 33741 2377 33775 2380
rect 33775 2377 33784 2380
rect 33732 2346 33741 2365
rect 33741 2346 33775 2365
rect 33775 2346 33784 2365
rect 33732 2313 33784 2346
rect 33732 2274 33741 2301
rect 33741 2274 33775 2301
rect 33775 2274 33784 2301
rect 33732 2249 33784 2274
rect 33732 2236 33784 2237
rect 33732 2202 33741 2236
rect 33741 2202 33775 2236
rect 33775 2202 33784 2236
rect 33732 2185 33784 2202
rect 33732 2164 33784 2173
rect 33732 2130 33741 2164
rect 33741 2130 33775 2164
rect 33775 2130 33784 2164
rect 33732 2121 33784 2130
rect 33732 2092 33784 2109
rect 33732 2058 33741 2092
rect 33741 2058 33775 2092
rect 33775 2058 33784 2092
rect 33732 2057 33784 2058
rect 33732 2020 33784 2045
rect 33732 1993 33741 2020
rect 33741 1993 33775 2020
rect 33775 1993 33784 2020
rect 33732 1948 33784 1981
rect 33732 1929 33741 1948
rect 33741 1929 33775 1948
rect 33775 1929 33784 1948
rect 33732 1914 33741 1917
rect 33741 1914 33775 1917
rect 33775 1914 33784 1917
rect 33732 1876 33784 1914
rect 33732 1865 33741 1876
rect 33741 1865 33775 1876
rect 33775 1865 33784 1876
rect 33732 1842 33741 1853
rect 33741 1842 33775 1853
rect 33775 1842 33784 1853
rect 33732 1804 33784 1842
rect 33732 1801 33741 1804
rect 33741 1801 33775 1804
rect 33775 1801 33784 1804
rect 33732 1770 33741 1789
rect 33741 1770 33775 1789
rect 33775 1770 33784 1789
rect 33732 1737 33784 1770
rect 33732 1698 33741 1725
rect 33741 1698 33775 1725
rect 33775 1698 33784 1725
rect 33732 1673 33784 1698
rect 33732 1660 33784 1661
rect 33732 1626 33741 1660
rect 33741 1626 33775 1660
rect 33775 1626 33784 1660
rect 33732 1609 33784 1626
rect 33732 1588 33784 1597
rect 33732 1554 33741 1588
rect 33741 1554 33775 1588
rect 33775 1554 33784 1588
rect 33732 1545 33784 1554
rect 33732 1516 33784 1533
rect 33732 1482 33741 1516
rect 33741 1482 33775 1516
rect 33775 1482 33784 1516
rect 33732 1481 33784 1482
rect 33732 1444 33784 1469
rect 33732 1417 33741 1444
rect 33741 1417 33775 1444
rect 33775 1417 33784 1444
rect 33732 1372 33784 1405
rect 33732 1353 33741 1372
rect 33741 1353 33775 1372
rect 33775 1353 33784 1372
rect 33732 1338 33741 1341
rect 33741 1338 33775 1341
rect 33775 1338 33784 1341
rect 33732 1300 33784 1338
rect 33732 1289 33741 1300
rect 33741 1289 33775 1300
rect 33775 1289 33784 1300
rect 33732 1266 33741 1277
rect 33741 1266 33775 1277
rect 33775 1266 33784 1277
rect 33732 1228 33784 1266
rect 33732 1225 33741 1228
rect 33741 1225 33775 1228
rect 33775 1225 33784 1228
rect 33732 1194 33741 1213
rect 33741 1194 33775 1213
rect 33775 1194 33784 1213
rect 33732 1161 33784 1194
rect 33828 3100 33880 3133
rect 33828 3081 33837 3100
rect 33837 3081 33871 3100
rect 33871 3081 33880 3100
rect 33828 3066 33837 3069
rect 33837 3066 33871 3069
rect 33871 3066 33880 3069
rect 33828 3028 33880 3066
rect 33828 3017 33837 3028
rect 33837 3017 33871 3028
rect 33871 3017 33880 3028
rect 33828 2994 33837 3005
rect 33837 2994 33871 3005
rect 33871 2994 33880 3005
rect 33828 2956 33880 2994
rect 33828 2953 33837 2956
rect 33837 2953 33871 2956
rect 33871 2953 33880 2956
rect 33828 2922 33837 2941
rect 33837 2922 33871 2941
rect 33871 2922 33880 2941
rect 33828 2889 33880 2922
rect 33828 2850 33837 2877
rect 33837 2850 33871 2877
rect 33871 2850 33880 2877
rect 33828 2825 33880 2850
rect 33828 2812 33880 2813
rect 33828 2778 33837 2812
rect 33837 2778 33871 2812
rect 33871 2778 33880 2812
rect 33828 2761 33880 2778
rect 33828 2740 33880 2749
rect 33828 2706 33837 2740
rect 33837 2706 33871 2740
rect 33871 2706 33880 2740
rect 33828 2697 33880 2706
rect 33828 2668 33880 2685
rect 33828 2634 33837 2668
rect 33837 2634 33871 2668
rect 33871 2634 33880 2668
rect 33828 2633 33880 2634
rect 33828 2596 33880 2621
rect 33828 2569 33837 2596
rect 33837 2569 33871 2596
rect 33871 2569 33880 2596
rect 33828 2524 33880 2557
rect 33828 2505 33837 2524
rect 33837 2505 33871 2524
rect 33871 2505 33880 2524
rect 33828 2490 33837 2493
rect 33837 2490 33871 2493
rect 33871 2490 33880 2493
rect 33828 2452 33880 2490
rect 33828 2441 33837 2452
rect 33837 2441 33871 2452
rect 33871 2441 33880 2452
rect 33828 2418 33837 2429
rect 33837 2418 33871 2429
rect 33871 2418 33880 2429
rect 33828 2380 33880 2418
rect 33828 2377 33837 2380
rect 33837 2377 33871 2380
rect 33871 2377 33880 2380
rect 33828 2346 33837 2365
rect 33837 2346 33871 2365
rect 33871 2346 33880 2365
rect 33828 2313 33880 2346
rect 33828 2274 33837 2301
rect 33837 2274 33871 2301
rect 33871 2274 33880 2301
rect 33828 2249 33880 2274
rect 33828 2236 33880 2237
rect 33828 2202 33837 2236
rect 33837 2202 33871 2236
rect 33871 2202 33880 2236
rect 33828 2185 33880 2202
rect 33828 2164 33880 2173
rect 33828 2130 33837 2164
rect 33837 2130 33871 2164
rect 33871 2130 33880 2164
rect 33828 2121 33880 2130
rect 33828 2092 33880 2109
rect 33828 2058 33837 2092
rect 33837 2058 33871 2092
rect 33871 2058 33880 2092
rect 33828 2057 33880 2058
rect 33828 2020 33880 2045
rect 33828 1993 33837 2020
rect 33837 1993 33871 2020
rect 33871 1993 33880 2020
rect 33828 1948 33880 1981
rect 33828 1929 33837 1948
rect 33837 1929 33871 1948
rect 33871 1929 33880 1948
rect 33828 1914 33837 1917
rect 33837 1914 33871 1917
rect 33871 1914 33880 1917
rect 33828 1876 33880 1914
rect 33828 1865 33837 1876
rect 33837 1865 33871 1876
rect 33871 1865 33880 1876
rect 33828 1842 33837 1853
rect 33837 1842 33871 1853
rect 33871 1842 33880 1853
rect 33828 1804 33880 1842
rect 33828 1801 33837 1804
rect 33837 1801 33871 1804
rect 33871 1801 33880 1804
rect 33828 1770 33837 1789
rect 33837 1770 33871 1789
rect 33871 1770 33880 1789
rect 33828 1737 33880 1770
rect 33828 1698 33837 1725
rect 33837 1698 33871 1725
rect 33871 1698 33880 1725
rect 33828 1673 33880 1698
rect 33828 1660 33880 1661
rect 33828 1626 33837 1660
rect 33837 1626 33871 1660
rect 33871 1626 33880 1660
rect 33828 1609 33880 1626
rect 33828 1588 33880 1597
rect 33828 1554 33837 1588
rect 33837 1554 33871 1588
rect 33871 1554 33880 1588
rect 33828 1545 33880 1554
rect 33828 1516 33880 1533
rect 33828 1482 33837 1516
rect 33837 1482 33871 1516
rect 33871 1482 33880 1516
rect 33828 1481 33880 1482
rect 33828 1444 33880 1469
rect 33828 1417 33837 1444
rect 33837 1417 33871 1444
rect 33871 1417 33880 1444
rect 33828 1372 33880 1405
rect 33828 1353 33837 1372
rect 33837 1353 33871 1372
rect 33871 1353 33880 1372
rect 33828 1338 33837 1341
rect 33837 1338 33871 1341
rect 33871 1338 33880 1341
rect 33828 1300 33880 1338
rect 33828 1289 33837 1300
rect 33837 1289 33871 1300
rect 33871 1289 33880 1300
rect 33828 1266 33837 1277
rect 33837 1266 33871 1277
rect 33871 1266 33880 1277
rect 33828 1228 33880 1266
rect 33828 1225 33837 1228
rect 33837 1225 33871 1228
rect 33871 1225 33880 1228
rect 33828 1194 33837 1213
rect 33837 1194 33871 1213
rect 33871 1194 33880 1213
rect 33828 1161 33880 1194
rect 33924 3100 33976 3133
rect 33924 3081 33933 3100
rect 33933 3081 33967 3100
rect 33967 3081 33976 3100
rect 33924 3066 33933 3069
rect 33933 3066 33967 3069
rect 33967 3066 33976 3069
rect 33924 3028 33976 3066
rect 33924 3017 33933 3028
rect 33933 3017 33967 3028
rect 33967 3017 33976 3028
rect 33924 2994 33933 3005
rect 33933 2994 33967 3005
rect 33967 2994 33976 3005
rect 33924 2956 33976 2994
rect 33924 2953 33933 2956
rect 33933 2953 33967 2956
rect 33967 2953 33976 2956
rect 33924 2922 33933 2941
rect 33933 2922 33967 2941
rect 33967 2922 33976 2941
rect 33924 2889 33976 2922
rect 33924 2850 33933 2877
rect 33933 2850 33967 2877
rect 33967 2850 33976 2877
rect 33924 2825 33976 2850
rect 33924 2812 33976 2813
rect 33924 2778 33933 2812
rect 33933 2778 33967 2812
rect 33967 2778 33976 2812
rect 33924 2761 33976 2778
rect 33924 2740 33976 2749
rect 33924 2706 33933 2740
rect 33933 2706 33967 2740
rect 33967 2706 33976 2740
rect 33924 2697 33976 2706
rect 33924 2668 33976 2685
rect 33924 2634 33933 2668
rect 33933 2634 33967 2668
rect 33967 2634 33976 2668
rect 33924 2633 33976 2634
rect 33924 2596 33976 2621
rect 33924 2569 33933 2596
rect 33933 2569 33967 2596
rect 33967 2569 33976 2596
rect 33924 2524 33976 2557
rect 33924 2505 33933 2524
rect 33933 2505 33967 2524
rect 33967 2505 33976 2524
rect 33924 2490 33933 2493
rect 33933 2490 33967 2493
rect 33967 2490 33976 2493
rect 33924 2452 33976 2490
rect 33924 2441 33933 2452
rect 33933 2441 33967 2452
rect 33967 2441 33976 2452
rect 33924 2418 33933 2429
rect 33933 2418 33967 2429
rect 33967 2418 33976 2429
rect 33924 2380 33976 2418
rect 33924 2377 33933 2380
rect 33933 2377 33967 2380
rect 33967 2377 33976 2380
rect 33924 2346 33933 2365
rect 33933 2346 33967 2365
rect 33967 2346 33976 2365
rect 33924 2313 33976 2346
rect 33924 2274 33933 2301
rect 33933 2274 33967 2301
rect 33967 2274 33976 2301
rect 33924 2249 33976 2274
rect 33924 2236 33976 2237
rect 33924 2202 33933 2236
rect 33933 2202 33967 2236
rect 33967 2202 33976 2236
rect 33924 2185 33976 2202
rect 33924 2164 33976 2173
rect 33924 2130 33933 2164
rect 33933 2130 33967 2164
rect 33967 2130 33976 2164
rect 33924 2121 33976 2130
rect 33924 2092 33976 2109
rect 33924 2058 33933 2092
rect 33933 2058 33967 2092
rect 33967 2058 33976 2092
rect 33924 2057 33976 2058
rect 33924 2020 33976 2045
rect 33924 1993 33933 2020
rect 33933 1993 33967 2020
rect 33967 1993 33976 2020
rect 33924 1948 33976 1981
rect 33924 1929 33933 1948
rect 33933 1929 33967 1948
rect 33967 1929 33976 1948
rect 33924 1914 33933 1917
rect 33933 1914 33967 1917
rect 33967 1914 33976 1917
rect 33924 1876 33976 1914
rect 33924 1865 33933 1876
rect 33933 1865 33967 1876
rect 33967 1865 33976 1876
rect 33924 1842 33933 1853
rect 33933 1842 33967 1853
rect 33967 1842 33976 1853
rect 33924 1804 33976 1842
rect 33924 1801 33933 1804
rect 33933 1801 33967 1804
rect 33967 1801 33976 1804
rect 33924 1770 33933 1789
rect 33933 1770 33967 1789
rect 33967 1770 33976 1789
rect 33924 1737 33976 1770
rect 33924 1698 33933 1725
rect 33933 1698 33967 1725
rect 33967 1698 33976 1725
rect 33924 1673 33976 1698
rect 33924 1660 33976 1661
rect 33924 1626 33933 1660
rect 33933 1626 33967 1660
rect 33967 1626 33976 1660
rect 33924 1609 33976 1626
rect 33924 1588 33976 1597
rect 33924 1554 33933 1588
rect 33933 1554 33967 1588
rect 33967 1554 33976 1588
rect 33924 1545 33976 1554
rect 33924 1516 33976 1533
rect 33924 1482 33933 1516
rect 33933 1482 33967 1516
rect 33967 1482 33976 1516
rect 33924 1481 33976 1482
rect 33924 1444 33976 1469
rect 33924 1417 33933 1444
rect 33933 1417 33967 1444
rect 33967 1417 33976 1444
rect 33924 1372 33976 1405
rect 33924 1353 33933 1372
rect 33933 1353 33967 1372
rect 33967 1353 33976 1372
rect 33924 1338 33933 1341
rect 33933 1338 33967 1341
rect 33967 1338 33976 1341
rect 33924 1300 33976 1338
rect 33924 1289 33933 1300
rect 33933 1289 33967 1300
rect 33967 1289 33976 1300
rect 33924 1266 33933 1277
rect 33933 1266 33967 1277
rect 33967 1266 33976 1277
rect 33924 1228 33976 1266
rect 33924 1225 33933 1228
rect 33933 1225 33967 1228
rect 33967 1225 33976 1228
rect 33924 1194 33933 1213
rect 33933 1194 33967 1213
rect 33967 1194 33976 1213
rect 33924 1161 33976 1194
rect 34020 3100 34072 3133
rect 34020 3081 34029 3100
rect 34029 3081 34063 3100
rect 34063 3081 34072 3100
rect 34020 3066 34029 3069
rect 34029 3066 34063 3069
rect 34063 3066 34072 3069
rect 34020 3028 34072 3066
rect 34020 3017 34029 3028
rect 34029 3017 34063 3028
rect 34063 3017 34072 3028
rect 34020 2994 34029 3005
rect 34029 2994 34063 3005
rect 34063 2994 34072 3005
rect 34020 2956 34072 2994
rect 34020 2953 34029 2956
rect 34029 2953 34063 2956
rect 34063 2953 34072 2956
rect 34020 2922 34029 2941
rect 34029 2922 34063 2941
rect 34063 2922 34072 2941
rect 34020 2889 34072 2922
rect 34020 2850 34029 2877
rect 34029 2850 34063 2877
rect 34063 2850 34072 2877
rect 34020 2825 34072 2850
rect 34020 2812 34072 2813
rect 34020 2778 34029 2812
rect 34029 2778 34063 2812
rect 34063 2778 34072 2812
rect 34020 2761 34072 2778
rect 34020 2740 34072 2749
rect 34020 2706 34029 2740
rect 34029 2706 34063 2740
rect 34063 2706 34072 2740
rect 34020 2697 34072 2706
rect 34020 2668 34072 2685
rect 34020 2634 34029 2668
rect 34029 2634 34063 2668
rect 34063 2634 34072 2668
rect 34020 2633 34072 2634
rect 34020 2596 34072 2621
rect 34020 2569 34029 2596
rect 34029 2569 34063 2596
rect 34063 2569 34072 2596
rect 34020 2524 34072 2557
rect 34020 2505 34029 2524
rect 34029 2505 34063 2524
rect 34063 2505 34072 2524
rect 34020 2490 34029 2493
rect 34029 2490 34063 2493
rect 34063 2490 34072 2493
rect 34020 2452 34072 2490
rect 34020 2441 34029 2452
rect 34029 2441 34063 2452
rect 34063 2441 34072 2452
rect 34020 2418 34029 2429
rect 34029 2418 34063 2429
rect 34063 2418 34072 2429
rect 34020 2380 34072 2418
rect 34020 2377 34029 2380
rect 34029 2377 34063 2380
rect 34063 2377 34072 2380
rect 34020 2346 34029 2365
rect 34029 2346 34063 2365
rect 34063 2346 34072 2365
rect 34020 2313 34072 2346
rect 34020 2274 34029 2301
rect 34029 2274 34063 2301
rect 34063 2274 34072 2301
rect 34020 2249 34072 2274
rect 34020 2236 34072 2237
rect 34020 2202 34029 2236
rect 34029 2202 34063 2236
rect 34063 2202 34072 2236
rect 34020 2185 34072 2202
rect 34020 2164 34072 2173
rect 34020 2130 34029 2164
rect 34029 2130 34063 2164
rect 34063 2130 34072 2164
rect 34020 2121 34072 2130
rect 34020 2092 34072 2109
rect 34020 2058 34029 2092
rect 34029 2058 34063 2092
rect 34063 2058 34072 2092
rect 34020 2057 34072 2058
rect 34020 2020 34072 2045
rect 34020 1993 34029 2020
rect 34029 1993 34063 2020
rect 34063 1993 34072 2020
rect 34020 1948 34072 1981
rect 34020 1929 34029 1948
rect 34029 1929 34063 1948
rect 34063 1929 34072 1948
rect 34020 1914 34029 1917
rect 34029 1914 34063 1917
rect 34063 1914 34072 1917
rect 34020 1876 34072 1914
rect 34020 1865 34029 1876
rect 34029 1865 34063 1876
rect 34063 1865 34072 1876
rect 34020 1842 34029 1853
rect 34029 1842 34063 1853
rect 34063 1842 34072 1853
rect 34020 1804 34072 1842
rect 34020 1801 34029 1804
rect 34029 1801 34063 1804
rect 34063 1801 34072 1804
rect 34020 1770 34029 1789
rect 34029 1770 34063 1789
rect 34063 1770 34072 1789
rect 34020 1737 34072 1770
rect 34020 1698 34029 1725
rect 34029 1698 34063 1725
rect 34063 1698 34072 1725
rect 34020 1673 34072 1698
rect 34020 1660 34072 1661
rect 34020 1626 34029 1660
rect 34029 1626 34063 1660
rect 34063 1626 34072 1660
rect 34020 1609 34072 1626
rect 34020 1588 34072 1597
rect 34020 1554 34029 1588
rect 34029 1554 34063 1588
rect 34063 1554 34072 1588
rect 34020 1545 34072 1554
rect 34020 1516 34072 1533
rect 34020 1482 34029 1516
rect 34029 1482 34063 1516
rect 34063 1482 34072 1516
rect 34020 1481 34072 1482
rect 34020 1444 34072 1469
rect 34020 1417 34029 1444
rect 34029 1417 34063 1444
rect 34063 1417 34072 1444
rect 34020 1372 34072 1405
rect 34020 1353 34029 1372
rect 34029 1353 34063 1372
rect 34063 1353 34072 1372
rect 34020 1338 34029 1341
rect 34029 1338 34063 1341
rect 34063 1338 34072 1341
rect 34020 1300 34072 1338
rect 34020 1289 34029 1300
rect 34029 1289 34063 1300
rect 34063 1289 34072 1300
rect 34020 1266 34029 1277
rect 34029 1266 34063 1277
rect 34063 1266 34072 1277
rect 34020 1228 34072 1266
rect 34020 1225 34029 1228
rect 34029 1225 34063 1228
rect 34063 1225 34072 1228
rect 34020 1194 34029 1213
rect 34029 1194 34063 1213
rect 34063 1194 34072 1213
rect 34020 1161 34072 1194
rect 34116 3100 34168 3133
rect 34116 3081 34125 3100
rect 34125 3081 34159 3100
rect 34159 3081 34168 3100
rect 34116 3066 34125 3069
rect 34125 3066 34159 3069
rect 34159 3066 34168 3069
rect 34116 3028 34168 3066
rect 34116 3017 34125 3028
rect 34125 3017 34159 3028
rect 34159 3017 34168 3028
rect 34116 2994 34125 3005
rect 34125 2994 34159 3005
rect 34159 2994 34168 3005
rect 34116 2956 34168 2994
rect 34116 2953 34125 2956
rect 34125 2953 34159 2956
rect 34159 2953 34168 2956
rect 34116 2922 34125 2941
rect 34125 2922 34159 2941
rect 34159 2922 34168 2941
rect 34116 2889 34168 2922
rect 34116 2850 34125 2877
rect 34125 2850 34159 2877
rect 34159 2850 34168 2877
rect 34116 2825 34168 2850
rect 34116 2812 34168 2813
rect 34116 2778 34125 2812
rect 34125 2778 34159 2812
rect 34159 2778 34168 2812
rect 34116 2761 34168 2778
rect 34116 2740 34168 2749
rect 34116 2706 34125 2740
rect 34125 2706 34159 2740
rect 34159 2706 34168 2740
rect 34116 2697 34168 2706
rect 34116 2668 34168 2685
rect 34116 2634 34125 2668
rect 34125 2634 34159 2668
rect 34159 2634 34168 2668
rect 34116 2633 34168 2634
rect 34116 2596 34168 2621
rect 34116 2569 34125 2596
rect 34125 2569 34159 2596
rect 34159 2569 34168 2596
rect 34116 2524 34168 2557
rect 34116 2505 34125 2524
rect 34125 2505 34159 2524
rect 34159 2505 34168 2524
rect 34116 2490 34125 2493
rect 34125 2490 34159 2493
rect 34159 2490 34168 2493
rect 34116 2452 34168 2490
rect 34116 2441 34125 2452
rect 34125 2441 34159 2452
rect 34159 2441 34168 2452
rect 34116 2418 34125 2429
rect 34125 2418 34159 2429
rect 34159 2418 34168 2429
rect 34116 2380 34168 2418
rect 34116 2377 34125 2380
rect 34125 2377 34159 2380
rect 34159 2377 34168 2380
rect 34116 2346 34125 2365
rect 34125 2346 34159 2365
rect 34159 2346 34168 2365
rect 34116 2313 34168 2346
rect 34116 2274 34125 2301
rect 34125 2274 34159 2301
rect 34159 2274 34168 2301
rect 34116 2249 34168 2274
rect 34116 2236 34168 2237
rect 34116 2202 34125 2236
rect 34125 2202 34159 2236
rect 34159 2202 34168 2236
rect 34116 2185 34168 2202
rect 34116 2164 34168 2173
rect 34116 2130 34125 2164
rect 34125 2130 34159 2164
rect 34159 2130 34168 2164
rect 34116 2121 34168 2130
rect 34116 2092 34168 2109
rect 34116 2058 34125 2092
rect 34125 2058 34159 2092
rect 34159 2058 34168 2092
rect 34116 2057 34168 2058
rect 34116 2020 34168 2045
rect 34116 1993 34125 2020
rect 34125 1993 34159 2020
rect 34159 1993 34168 2020
rect 34116 1948 34168 1981
rect 34116 1929 34125 1948
rect 34125 1929 34159 1948
rect 34159 1929 34168 1948
rect 34116 1914 34125 1917
rect 34125 1914 34159 1917
rect 34159 1914 34168 1917
rect 34116 1876 34168 1914
rect 34116 1865 34125 1876
rect 34125 1865 34159 1876
rect 34159 1865 34168 1876
rect 34116 1842 34125 1853
rect 34125 1842 34159 1853
rect 34159 1842 34168 1853
rect 34116 1804 34168 1842
rect 34116 1801 34125 1804
rect 34125 1801 34159 1804
rect 34159 1801 34168 1804
rect 34116 1770 34125 1789
rect 34125 1770 34159 1789
rect 34159 1770 34168 1789
rect 34116 1737 34168 1770
rect 34116 1698 34125 1725
rect 34125 1698 34159 1725
rect 34159 1698 34168 1725
rect 34116 1673 34168 1698
rect 34116 1660 34168 1661
rect 34116 1626 34125 1660
rect 34125 1626 34159 1660
rect 34159 1626 34168 1660
rect 34116 1609 34168 1626
rect 34116 1588 34168 1597
rect 34116 1554 34125 1588
rect 34125 1554 34159 1588
rect 34159 1554 34168 1588
rect 34116 1545 34168 1554
rect 34116 1516 34168 1533
rect 34116 1482 34125 1516
rect 34125 1482 34159 1516
rect 34159 1482 34168 1516
rect 34116 1481 34168 1482
rect 34116 1444 34168 1469
rect 34116 1417 34125 1444
rect 34125 1417 34159 1444
rect 34159 1417 34168 1444
rect 34116 1372 34168 1405
rect 34116 1353 34125 1372
rect 34125 1353 34159 1372
rect 34159 1353 34168 1372
rect 34116 1338 34125 1341
rect 34125 1338 34159 1341
rect 34159 1338 34168 1341
rect 34116 1300 34168 1338
rect 34116 1289 34125 1300
rect 34125 1289 34159 1300
rect 34159 1289 34168 1300
rect 34116 1266 34125 1277
rect 34125 1266 34159 1277
rect 34159 1266 34168 1277
rect 34116 1228 34168 1266
rect 34116 1225 34125 1228
rect 34125 1225 34159 1228
rect 34159 1225 34168 1228
rect 34116 1194 34125 1213
rect 34125 1194 34159 1213
rect 34159 1194 34168 1213
rect 34116 1161 34168 1194
rect 34212 3100 34264 3133
rect 34212 3081 34221 3100
rect 34221 3081 34255 3100
rect 34255 3081 34264 3100
rect 34212 3066 34221 3069
rect 34221 3066 34255 3069
rect 34255 3066 34264 3069
rect 34212 3028 34264 3066
rect 34212 3017 34221 3028
rect 34221 3017 34255 3028
rect 34255 3017 34264 3028
rect 34212 2994 34221 3005
rect 34221 2994 34255 3005
rect 34255 2994 34264 3005
rect 34212 2956 34264 2994
rect 34212 2953 34221 2956
rect 34221 2953 34255 2956
rect 34255 2953 34264 2956
rect 34212 2922 34221 2941
rect 34221 2922 34255 2941
rect 34255 2922 34264 2941
rect 34212 2889 34264 2922
rect 34212 2850 34221 2877
rect 34221 2850 34255 2877
rect 34255 2850 34264 2877
rect 34212 2825 34264 2850
rect 34212 2812 34264 2813
rect 34212 2778 34221 2812
rect 34221 2778 34255 2812
rect 34255 2778 34264 2812
rect 34212 2761 34264 2778
rect 34212 2740 34264 2749
rect 34212 2706 34221 2740
rect 34221 2706 34255 2740
rect 34255 2706 34264 2740
rect 34212 2697 34264 2706
rect 34212 2668 34264 2685
rect 34212 2634 34221 2668
rect 34221 2634 34255 2668
rect 34255 2634 34264 2668
rect 34212 2633 34264 2634
rect 34212 2596 34264 2621
rect 34212 2569 34221 2596
rect 34221 2569 34255 2596
rect 34255 2569 34264 2596
rect 34212 2524 34264 2557
rect 34212 2505 34221 2524
rect 34221 2505 34255 2524
rect 34255 2505 34264 2524
rect 34212 2490 34221 2493
rect 34221 2490 34255 2493
rect 34255 2490 34264 2493
rect 34212 2452 34264 2490
rect 34212 2441 34221 2452
rect 34221 2441 34255 2452
rect 34255 2441 34264 2452
rect 34212 2418 34221 2429
rect 34221 2418 34255 2429
rect 34255 2418 34264 2429
rect 34212 2380 34264 2418
rect 34212 2377 34221 2380
rect 34221 2377 34255 2380
rect 34255 2377 34264 2380
rect 34212 2346 34221 2365
rect 34221 2346 34255 2365
rect 34255 2346 34264 2365
rect 34212 2313 34264 2346
rect 34212 2274 34221 2301
rect 34221 2274 34255 2301
rect 34255 2274 34264 2301
rect 34212 2249 34264 2274
rect 34212 2236 34264 2237
rect 34212 2202 34221 2236
rect 34221 2202 34255 2236
rect 34255 2202 34264 2236
rect 34212 2185 34264 2202
rect 34212 2164 34264 2173
rect 34212 2130 34221 2164
rect 34221 2130 34255 2164
rect 34255 2130 34264 2164
rect 34212 2121 34264 2130
rect 34212 2092 34264 2109
rect 34212 2058 34221 2092
rect 34221 2058 34255 2092
rect 34255 2058 34264 2092
rect 34212 2057 34264 2058
rect 34212 2020 34264 2045
rect 34212 1993 34221 2020
rect 34221 1993 34255 2020
rect 34255 1993 34264 2020
rect 34212 1948 34264 1981
rect 34212 1929 34221 1948
rect 34221 1929 34255 1948
rect 34255 1929 34264 1948
rect 34212 1914 34221 1917
rect 34221 1914 34255 1917
rect 34255 1914 34264 1917
rect 34212 1876 34264 1914
rect 34212 1865 34221 1876
rect 34221 1865 34255 1876
rect 34255 1865 34264 1876
rect 34212 1842 34221 1853
rect 34221 1842 34255 1853
rect 34255 1842 34264 1853
rect 34212 1804 34264 1842
rect 34212 1801 34221 1804
rect 34221 1801 34255 1804
rect 34255 1801 34264 1804
rect 34212 1770 34221 1789
rect 34221 1770 34255 1789
rect 34255 1770 34264 1789
rect 34212 1737 34264 1770
rect 34212 1698 34221 1725
rect 34221 1698 34255 1725
rect 34255 1698 34264 1725
rect 34212 1673 34264 1698
rect 34212 1660 34264 1661
rect 34212 1626 34221 1660
rect 34221 1626 34255 1660
rect 34255 1626 34264 1660
rect 34212 1609 34264 1626
rect 34212 1588 34264 1597
rect 34212 1554 34221 1588
rect 34221 1554 34255 1588
rect 34255 1554 34264 1588
rect 34212 1545 34264 1554
rect 34212 1516 34264 1533
rect 34212 1482 34221 1516
rect 34221 1482 34255 1516
rect 34255 1482 34264 1516
rect 34212 1481 34264 1482
rect 34212 1444 34264 1469
rect 34212 1417 34221 1444
rect 34221 1417 34255 1444
rect 34255 1417 34264 1444
rect 34212 1372 34264 1405
rect 34212 1353 34221 1372
rect 34221 1353 34255 1372
rect 34255 1353 34264 1372
rect 34212 1338 34221 1341
rect 34221 1338 34255 1341
rect 34255 1338 34264 1341
rect 34212 1300 34264 1338
rect 34212 1289 34221 1300
rect 34221 1289 34255 1300
rect 34255 1289 34264 1300
rect 34212 1266 34221 1277
rect 34221 1266 34255 1277
rect 34255 1266 34264 1277
rect 34212 1228 34264 1266
rect 34212 1225 34221 1228
rect 34221 1225 34255 1228
rect 34255 1225 34264 1228
rect 34212 1194 34221 1213
rect 34221 1194 34255 1213
rect 34255 1194 34264 1213
rect 34212 1161 34264 1194
rect 34308 3100 34360 3133
rect 34308 3081 34317 3100
rect 34317 3081 34351 3100
rect 34351 3081 34360 3100
rect 34308 3066 34317 3069
rect 34317 3066 34351 3069
rect 34351 3066 34360 3069
rect 34308 3028 34360 3066
rect 34308 3017 34317 3028
rect 34317 3017 34351 3028
rect 34351 3017 34360 3028
rect 34308 2994 34317 3005
rect 34317 2994 34351 3005
rect 34351 2994 34360 3005
rect 34308 2956 34360 2994
rect 34308 2953 34317 2956
rect 34317 2953 34351 2956
rect 34351 2953 34360 2956
rect 34308 2922 34317 2941
rect 34317 2922 34351 2941
rect 34351 2922 34360 2941
rect 34308 2889 34360 2922
rect 34308 2850 34317 2877
rect 34317 2850 34351 2877
rect 34351 2850 34360 2877
rect 34308 2825 34360 2850
rect 34308 2812 34360 2813
rect 34308 2778 34317 2812
rect 34317 2778 34351 2812
rect 34351 2778 34360 2812
rect 34308 2761 34360 2778
rect 34308 2740 34360 2749
rect 34308 2706 34317 2740
rect 34317 2706 34351 2740
rect 34351 2706 34360 2740
rect 34308 2697 34360 2706
rect 34308 2668 34360 2685
rect 34308 2634 34317 2668
rect 34317 2634 34351 2668
rect 34351 2634 34360 2668
rect 34308 2633 34360 2634
rect 34308 2596 34360 2621
rect 34308 2569 34317 2596
rect 34317 2569 34351 2596
rect 34351 2569 34360 2596
rect 34308 2524 34360 2557
rect 34308 2505 34317 2524
rect 34317 2505 34351 2524
rect 34351 2505 34360 2524
rect 34308 2490 34317 2493
rect 34317 2490 34351 2493
rect 34351 2490 34360 2493
rect 34308 2452 34360 2490
rect 34308 2441 34317 2452
rect 34317 2441 34351 2452
rect 34351 2441 34360 2452
rect 34308 2418 34317 2429
rect 34317 2418 34351 2429
rect 34351 2418 34360 2429
rect 34308 2380 34360 2418
rect 34308 2377 34317 2380
rect 34317 2377 34351 2380
rect 34351 2377 34360 2380
rect 34308 2346 34317 2365
rect 34317 2346 34351 2365
rect 34351 2346 34360 2365
rect 34308 2313 34360 2346
rect 34308 2274 34317 2301
rect 34317 2274 34351 2301
rect 34351 2274 34360 2301
rect 34308 2249 34360 2274
rect 34308 2236 34360 2237
rect 34308 2202 34317 2236
rect 34317 2202 34351 2236
rect 34351 2202 34360 2236
rect 34308 2185 34360 2202
rect 34308 2164 34360 2173
rect 34308 2130 34317 2164
rect 34317 2130 34351 2164
rect 34351 2130 34360 2164
rect 34308 2121 34360 2130
rect 34308 2092 34360 2109
rect 34308 2058 34317 2092
rect 34317 2058 34351 2092
rect 34351 2058 34360 2092
rect 34308 2057 34360 2058
rect 34308 2020 34360 2045
rect 34308 1993 34317 2020
rect 34317 1993 34351 2020
rect 34351 1993 34360 2020
rect 34308 1948 34360 1981
rect 34308 1929 34317 1948
rect 34317 1929 34351 1948
rect 34351 1929 34360 1948
rect 34308 1914 34317 1917
rect 34317 1914 34351 1917
rect 34351 1914 34360 1917
rect 34308 1876 34360 1914
rect 34308 1865 34317 1876
rect 34317 1865 34351 1876
rect 34351 1865 34360 1876
rect 34308 1842 34317 1853
rect 34317 1842 34351 1853
rect 34351 1842 34360 1853
rect 34308 1804 34360 1842
rect 34308 1801 34317 1804
rect 34317 1801 34351 1804
rect 34351 1801 34360 1804
rect 34308 1770 34317 1789
rect 34317 1770 34351 1789
rect 34351 1770 34360 1789
rect 34308 1737 34360 1770
rect 34308 1698 34317 1725
rect 34317 1698 34351 1725
rect 34351 1698 34360 1725
rect 34308 1673 34360 1698
rect 34308 1660 34360 1661
rect 34308 1626 34317 1660
rect 34317 1626 34351 1660
rect 34351 1626 34360 1660
rect 34308 1609 34360 1626
rect 34308 1588 34360 1597
rect 34308 1554 34317 1588
rect 34317 1554 34351 1588
rect 34351 1554 34360 1588
rect 34308 1545 34360 1554
rect 34308 1516 34360 1533
rect 34308 1482 34317 1516
rect 34317 1482 34351 1516
rect 34351 1482 34360 1516
rect 34308 1481 34360 1482
rect 34308 1444 34360 1469
rect 34308 1417 34317 1444
rect 34317 1417 34351 1444
rect 34351 1417 34360 1444
rect 34308 1372 34360 1405
rect 34308 1353 34317 1372
rect 34317 1353 34351 1372
rect 34351 1353 34360 1372
rect 34308 1338 34317 1341
rect 34317 1338 34351 1341
rect 34351 1338 34360 1341
rect 34308 1300 34360 1338
rect 34308 1289 34317 1300
rect 34317 1289 34351 1300
rect 34351 1289 34360 1300
rect 34308 1266 34317 1277
rect 34317 1266 34351 1277
rect 34351 1266 34360 1277
rect 34308 1228 34360 1266
rect 34308 1225 34317 1228
rect 34317 1225 34351 1228
rect 34351 1225 34360 1228
rect 34308 1194 34317 1213
rect 34317 1194 34351 1213
rect 34351 1194 34360 1213
rect 34308 1161 34360 1194
rect 34404 3100 34456 3133
rect 34404 3081 34413 3100
rect 34413 3081 34447 3100
rect 34447 3081 34456 3100
rect 34404 3066 34413 3069
rect 34413 3066 34447 3069
rect 34447 3066 34456 3069
rect 34404 3028 34456 3066
rect 34404 3017 34413 3028
rect 34413 3017 34447 3028
rect 34447 3017 34456 3028
rect 34404 2994 34413 3005
rect 34413 2994 34447 3005
rect 34447 2994 34456 3005
rect 34404 2956 34456 2994
rect 34404 2953 34413 2956
rect 34413 2953 34447 2956
rect 34447 2953 34456 2956
rect 34404 2922 34413 2941
rect 34413 2922 34447 2941
rect 34447 2922 34456 2941
rect 34404 2889 34456 2922
rect 34404 2850 34413 2877
rect 34413 2850 34447 2877
rect 34447 2850 34456 2877
rect 34404 2825 34456 2850
rect 34404 2812 34456 2813
rect 34404 2778 34413 2812
rect 34413 2778 34447 2812
rect 34447 2778 34456 2812
rect 34404 2761 34456 2778
rect 34404 2740 34456 2749
rect 34404 2706 34413 2740
rect 34413 2706 34447 2740
rect 34447 2706 34456 2740
rect 34404 2697 34456 2706
rect 34404 2668 34456 2685
rect 34404 2634 34413 2668
rect 34413 2634 34447 2668
rect 34447 2634 34456 2668
rect 34404 2633 34456 2634
rect 34404 2596 34456 2621
rect 34404 2569 34413 2596
rect 34413 2569 34447 2596
rect 34447 2569 34456 2596
rect 34404 2524 34456 2557
rect 34404 2505 34413 2524
rect 34413 2505 34447 2524
rect 34447 2505 34456 2524
rect 34404 2490 34413 2493
rect 34413 2490 34447 2493
rect 34447 2490 34456 2493
rect 34404 2452 34456 2490
rect 34404 2441 34413 2452
rect 34413 2441 34447 2452
rect 34447 2441 34456 2452
rect 34404 2418 34413 2429
rect 34413 2418 34447 2429
rect 34447 2418 34456 2429
rect 34404 2380 34456 2418
rect 34404 2377 34413 2380
rect 34413 2377 34447 2380
rect 34447 2377 34456 2380
rect 34404 2346 34413 2365
rect 34413 2346 34447 2365
rect 34447 2346 34456 2365
rect 34404 2313 34456 2346
rect 34404 2274 34413 2301
rect 34413 2274 34447 2301
rect 34447 2274 34456 2301
rect 34404 2249 34456 2274
rect 34404 2236 34456 2237
rect 34404 2202 34413 2236
rect 34413 2202 34447 2236
rect 34447 2202 34456 2236
rect 34404 2185 34456 2202
rect 34404 2164 34456 2173
rect 34404 2130 34413 2164
rect 34413 2130 34447 2164
rect 34447 2130 34456 2164
rect 34404 2121 34456 2130
rect 34404 2092 34456 2109
rect 34404 2058 34413 2092
rect 34413 2058 34447 2092
rect 34447 2058 34456 2092
rect 34404 2057 34456 2058
rect 34404 2020 34456 2045
rect 34404 1993 34413 2020
rect 34413 1993 34447 2020
rect 34447 1993 34456 2020
rect 34404 1948 34456 1981
rect 34404 1929 34413 1948
rect 34413 1929 34447 1948
rect 34447 1929 34456 1948
rect 34404 1914 34413 1917
rect 34413 1914 34447 1917
rect 34447 1914 34456 1917
rect 34404 1876 34456 1914
rect 34404 1865 34413 1876
rect 34413 1865 34447 1876
rect 34447 1865 34456 1876
rect 34404 1842 34413 1853
rect 34413 1842 34447 1853
rect 34447 1842 34456 1853
rect 34404 1804 34456 1842
rect 34404 1801 34413 1804
rect 34413 1801 34447 1804
rect 34447 1801 34456 1804
rect 34404 1770 34413 1789
rect 34413 1770 34447 1789
rect 34447 1770 34456 1789
rect 34404 1737 34456 1770
rect 34404 1698 34413 1725
rect 34413 1698 34447 1725
rect 34447 1698 34456 1725
rect 34404 1673 34456 1698
rect 34404 1660 34456 1661
rect 34404 1626 34413 1660
rect 34413 1626 34447 1660
rect 34447 1626 34456 1660
rect 34404 1609 34456 1626
rect 34404 1588 34456 1597
rect 34404 1554 34413 1588
rect 34413 1554 34447 1588
rect 34447 1554 34456 1588
rect 34404 1545 34456 1554
rect 34404 1516 34456 1533
rect 34404 1482 34413 1516
rect 34413 1482 34447 1516
rect 34447 1482 34456 1516
rect 34404 1481 34456 1482
rect 34404 1444 34456 1469
rect 34404 1417 34413 1444
rect 34413 1417 34447 1444
rect 34447 1417 34456 1444
rect 34404 1372 34456 1405
rect 34404 1353 34413 1372
rect 34413 1353 34447 1372
rect 34447 1353 34456 1372
rect 34404 1338 34413 1341
rect 34413 1338 34447 1341
rect 34447 1338 34456 1341
rect 34404 1300 34456 1338
rect 34404 1289 34413 1300
rect 34413 1289 34447 1300
rect 34447 1289 34456 1300
rect 34404 1266 34413 1277
rect 34413 1266 34447 1277
rect 34447 1266 34456 1277
rect 34404 1228 34456 1266
rect 34404 1225 34413 1228
rect 34413 1225 34447 1228
rect 34447 1225 34456 1228
rect 34404 1194 34413 1213
rect 34413 1194 34447 1213
rect 34447 1194 34456 1213
rect 34404 1161 34456 1194
rect 34500 3100 34552 3133
rect 34500 3081 34509 3100
rect 34509 3081 34543 3100
rect 34543 3081 34552 3100
rect 34500 3066 34509 3069
rect 34509 3066 34543 3069
rect 34543 3066 34552 3069
rect 34500 3028 34552 3066
rect 34500 3017 34509 3028
rect 34509 3017 34543 3028
rect 34543 3017 34552 3028
rect 34500 2994 34509 3005
rect 34509 2994 34543 3005
rect 34543 2994 34552 3005
rect 34500 2956 34552 2994
rect 34500 2953 34509 2956
rect 34509 2953 34543 2956
rect 34543 2953 34552 2956
rect 34500 2922 34509 2941
rect 34509 2922 34543 2941
rect 34543 2922 34552 2941
rect 34500 2889 34552 2922
rect 34500 2850 34509 2877
rect 34509 2850 34543 2877
rect 34543 2850 34552 2877
rect 34500 2825 34552 2850
rect 34500 2812 34552 2813
rect 34500 2778 34509 2812
rect 34509 2778 34543 2812
rect 34543 2778 34552 2812
rect 34500 2761 34552 2778
rect 34500 2740 34552 2749
rect 34500 2706 34509 2740
rect 34509 2706 34543 2740
rect 34543 2706 34552 2740
rect 34500 2697 34552 2706
rect 34500 2668 34552 2685
rect 34500 2634 34509 2668
rect 34509 2634 34543 2668
rect 34543 2634 34552 2668
rect 34500 2633 34552 2634
rect 34500 2596 34552 2621
rect 34500 2569 34509 2596
rect 34509 2569 34543 2596
rect 34543 2569 34552 2596
rect 34500 2524 34552 2557
rect 34500 2505 34509 2524
rect 34509 2505 34543 2524
rect 34543 2505 34552 2524
rect 34500 2490 34509 2493
rect 34509 2490 34543 2493
rect 34543 2490 34552 2493
rect 34500 2452 34552 2490
rect 34500 2441 34509 2452
rect 34509 2441 34543 2452
rect 34543 2441 34552 2452
rect 34500 2418 34509 2429
rect 34509 2418 34543 2429
rect 34543 2418 34552 2429
rect 34500 2380 34552 2418
rect 34500 2377 34509 2380
rect 34509 2377 34543 2380
rect 34543 2377 34552 2380
rect 34500 2346 34509 2365
rect 34509 2346 34543 2365
rect 34543 2346 34552 2365
rect 34500 2313 34552 2346
rect 34500 2274 34509 2301
rect 34509 2274 34543 2301
rect 34543 2274 34552 2301
rect 34500 2249 34552 2274
rect 34500 2236 34552 2237
rect 34500 2202 34509 2236
rect 34509 2202 34543 2236
rect 34543 2202 34552 2236
rect 34500 2185 34552 2202
rect 34500 2164 34552 2173
rect 34500 2130 34509 2164
rect 34509 2130 34543 2164
rect 34543 2130 34552 2164
rect 34500 2121 34552 2130
rect 34500 2092 34552 2109
rect 34500 2058 34509 2092
rect 34509 2058 34543 2092
rect 34543 2058 34552 2092
rect 34500 2057 34552 2058
rect 34500 2020 34552 2045
rect 34500 1993 34509 2020
rect 34509 1993 34543 2020
rect 34543 1993 34552 2020
rect 34500 1948 34552 1981
rect 34500 1929 34509 1948
rect 34509 1929 34543 1948
rect 34543 1929 34552 1948
rect 34500 1914 34509 1917
rect 34509 1914 34543 1917
rect 34543 1914 34552 1917
rect 34500 1876 34552 1914
rect 34500 1865 34509 1876
rect 34509 1865 34543 1876
rect 34543 1865 34552 1876
rect 34500 1842 34509 1853
rect 34509 1842 34543 1853
rect 34543 1842 34552 1853
rect 34500 1804 34552 1842
rect 34500 1801 34509 1804
rect 34509 1801 34543 1804
rect 34543 1801 34552 1804
rect 34500 1770 34509 1789
rect 34509 1770 34543 1789
rect 34543 1770 34552 1789
rect 34500 1737 34552 1770
rect 34500 1698 34509 1725
rect 34509 1698 34543 1725
rect 34543 1698 34552 1725
rect 34500 1673 34552 1698
rect 34500 1660 34552 1661
rect 34500 1626 34509 1660
rect 34509 1626 34543 1660
rect 34543 1626 34552 1660
rect 34500 1609 34552 1626
rect 34500 1588 34552 1597
rect 34500 1554 34509 1588
rect 34509 1554 34543 1588
rect 34543 1554 34552 1588
rect 34500 1545 34552 1554
rect 34500 1516 34552 1533
rect 34500 1482 34509 1516
rect 34509 1482 34543 1516
rect 34543 1482 34552 1516
rect 34500 1481 34552 1482
rect 34500 1444 34552 1469
rect 34500 1417 34509 1444
rect 34509 1417 34543 1444
rect 34543 1417 34552 1444
rect 34500 1372 34552 1405
rect 34500 1353 34509 1372
rect 34509 1353 34543 1372
rect 34543 1353 34552 1372
rect 34500 1338 34509 1341
rect 34509 1338 34543 1341
rect 34543 1338 34552 1341
rect 34500 1300 34552 1338
rect 34500 1289 34509 1300
rect 34509 1289 34543 1300
rect 34543 1289 34552 1300
rect 34500 1266 34509 1277
rect 34509 1266 34543 1277
rect 34543 1266 34552 1277
rect 34500 1228 34552 1266
rect 34500 1225 34509 1228
rect 34509 1225 34543 1228
rect 34543 1225 34552 1228
rect 34500 1194 34509 1213
rect 34509 1194 34543 1213
rect 34543 1194 34552 1213
rect 34500 1161 34552 1194
rect 34596 3100 34648 3133
rect 34596 3081 34605 3100
rect 34605 3081 34639 3100
rect 34639 3081 34648 3100
rect 34596 3066 34605 3069
rect 34605 3066 34639 3069
rect 34639 3066 34648 3069
rect 34596 3028 34648 3066
rect 34596 3017 34605 3028
rect 34605 3017 34639 3028
rect 34639 3017 34648 3028
rect 34596 2994 34605 3005
rect 34605 2994 34639 3005
rect 34639 2994 34648 3005
rect 34596 2956 34648 2994
rect 34596 2953 34605 2956
rect 34605 2953 34639 2956
rect 34639 2953 34648 2956
rect 34596 2922 34605 2941
rect 34605 2922 34639 2941
rect 34639 2922 34648 2941
rect 34596 2889 34648 2922
rect 34596 2850 34605 2877
rect 34605 2850 34639 2877
rect 34639 2850 34648 2877
rect 34596 2825 34648 2850
rect 34596 2812 34648 2813
rect 34596 2778 34605 2812
rect 34605 2778 34639 2812
rect 34639 2778 34648 2812
rect 34596 2761 34648 2778
rect 34596 2740 34648 2749
rect 34596 2706 34605 2740
rect 34605 2706 34639 2740
rect 34639 2706 34648 2740
rect 34596 2697 34648 2706
rect 34596 2668 34648 2685
rect 34596 2634 34605 2668
rect 34605 2634 34639 2668
rect 34639 2634 34648 2668
rect 34596 2633 34648 2634
rect 34596 2596 34648 2621
rect 34596 2569 34605 2596
rect 34605 2569 34639 2596
rect 34639 2569 34648 2596
rect 34596 2524 34648 2557
rect 34596 2505 34605 2524
rect 34605 2505 34639 2524
rect 34639 2505 34648 2524
rect 34596 2490 34605 2493
rect 34605 2490 34639 2493
rect 34639 2490 34648 2493
rect 34596 2452 34648 2490
rect 34596 2441 34605 2452
rect 34605 2441 34639 2452
rect 34639 2441 34648 2452
rect 34596 2418 34605 2429
rect 34605 2418 34639 2429
rect 34639 2418 34648 2429
rect 34596 2380 34648 2418
rect 34596 2377 34605 2380
rect 34605 2377 34639 2380
rect 34639 2377 34648 2380
rect 34596 2346 34605 2365
rect 34605 2346 34639 2365
rect 34639 2346 34648 2365
rect 34596 2313 34648 2346
rect 34596 2274 34605 2301
rect 34605 2274 34639 2301
rect 34639 2274 34648 2301
rect 34596 2249 34648 2274
rect 34596 2236 34648 2237
rect 34596 2202 34605 2236
rect 34605 2202 34639 2236
rect 34639 2202 34648 2236
rect 34596 2185 34648 2202
rect 34596 2164 34648 2173
rect 34596 2130 34605 2164
rect 34605 2130 34639 2164
rect 34639 2130 34648 2164
rect 34596 2121 34648 2130
rect 34596 2092 34648 2109
rect 34596 2058 34605 2092
rect 34605 2058 34639 2092
rect 34639 2058 34648 2092
rect 34596 2057 34648 2058
rect 34596 2020 34648 2045
rect 34596 1993 34605 2020
rect 34605 1993 34639 2020
rect 34639 1993 34648 2020
rect 34596 1948 34648 1981
rect 34596 1929 34605 1948
rect 34605 1929 34639 1948
rect 34639 1929 34648 1948
rect 34596 1914 34605 1917
rect 34605 1914 34639 1917
rect 34639 1914 34648 1917
rect 34596 1876 34648 1914
rect 34596 1865 34605 1876
rect 34605 1865 34639 1876
rect 34639 1865 34648 1876
rect 34596 1842 34605 1853
rect 34605 1842 34639 1853
rect 34639 1842 34648 1853
rect 34596 1804 34648 1842
rect 34596 1801 34605 1804
rect 34605 1801 34639 1804
rect 34639 1801 34648 1804
rect 34596 1770 34605 1789
rect 34605 1770 34639 1789
rect 34639 1770 34648 1789
rect 34596 1737 34648 1770
rect 34596 1698 34605 1725
rect 34605 1698 34639 1725
rect 34639 1698 34648 1725
rect 34596 1673 34648 1698
rect 34596 1660 34648 1661
rect 34596 1626 34605 1660
rect 34605 1626 34639 1660
rect 34639 1626 34648 1660
rect 34596 1609 34648 1626
rect 34596 1588 34648 1597
rect 34596 1554 34605 1588
rect 34605 1554 34639 1588
rect 34639 1554 34648 1588
rect 34596 1545 34648 1554
rect 34596 1516 34648 1533
rect 34596 1482 34605 1516
rect 34605 1482 34639 1516
rect 34639 1482 34648 1516
rect 34596 1481 34648 1482
rect 34596 1444 34648 1469
rect 34596 1417 34605 1444
rect 34605 1417 34639 1444
rect 34639 1417 34648 1444
rect 34596 1372 34648 1405
rect 34596 1353 34605 1372
rect 34605 1353 34639 1372
rect 34639 1353 34648 1372
rect 34596 1338 34605 1341
rect 34605 1338 34639 1341
rect 34639 1338 34648 1341
rect 34596 1300 34648 1338
rect 34596 1289 34605 1300
rect 34605 1289 34639 1300
rect 34639 1289 34648 1300
rect 34596 1266 34605 1277
rect 34605 1266 34639 1277
rect 34639 1266 34648 1277
rect 34596 1228 34648 1266
rect 34596 1225 34605 1228
rect 34605 1225 34639 1228
rect 34639 1225 34648 1228
rect 34596 1194 34605 1213
rect 34605 1194 34639 1213
rect 34639 1194 34648 1213
rect 34596 1161 34648 1194
rect 34692 3100 34744 3133
rect 34692 3081 34701 3100
rect 34701 3081 34735 3100
rect 34735 3081 34744 3100
rect 34692 3066 34701 3069
rect 34701 3066 34735 3069
rect 34735 3066 34744 3069
rect 34692 3028 34744 3066
rect 34692 3017 34701 3028
rect 34701 3017 34735 3028
rect 34735 3017 34744 3028
rect 34692 2994 34701 3005
rect 34701 2994 34735 3005
rect 34735 2994 34744 3005
rect 34692 2956 34744 2994
rect 34692 2953 34701 2956
rect 34701 2953 34735 2956
rect 34735 2953 34744 2956
rect 34692 2922 34701 2941
rect 34701 2922 34735 2941
rect 34735 2922 34744 2941
rect 34692 2889 34744 2922
rect 34692 2850 34701 2877
rect 34701 2850 34735 2877
rect 34735 2850 34744 2877
rect 34692 2825 34744 2850
rect 34692 2812 34744 2813
rect 34692 2778 34701 2812
rect 34701 2778 34735 2812
rect 34735 2778 34744 2812
rect 34692 2761 34744 2778
rect 34692 2740 34744 2749
rect 34692 2706 34701 2740
rect 34701 2706 34735 2740
rect 34735 2706 34744 2740
rect 34692 2697 34744 2706
rect 34692 2668 34744 2685
rect 34692 2634 34701 2668
rect 34701 2634 34735 2668
rect 34735 2634 34744 2668
rect 34692 2633 34744 2634
rect 34692 2596 34744 2621
rect 34692 2569 34701 2596
rect 34701 2569 34735 2596
rect 34735 2569 34744 2596
rect 34692 2524 34744 2557
rect 34692 2505 34701 2524
rect 34701 2505 34735 2524
rect 34735 2505 34744 2524
rect 34692 2490 34701 2493
rect 34701 2490 34735 2493
rect 34735 2490 34744 2493
rect 34692 2452 34744 2490
rect 34692 2441 34701 2452
rect 34701 2441 34735 2452
rect 34735 2441 34744 2452
rect 34692 2418 34701 2429
rect 34701 2418 34735 2429
rect 34735 2418 34744 2429
rect 34692 2380 34744 2418
rect 34692 2377 34701 2380
rect 34701 2377 34735 2380
rect 34735 2377 34744 2380
rect 34692 2346 34701 2365
rect 34701 2346 34735 2365
rect 34735 2346 34744 2365
rect 34692 2313 34744 2346
rect 34692 2274 34701 2301
rect 34701 2274 34735 2301
rect 34735 2274 34744 2301
rect 34692 2249 34744 2274
rect 34692 2236 34744 2237
rect 34692 2202 34701 2236
rect 34701 2202 34735 2236
rect 34735 2202 34744 2236
rect 34692 2185 34744 2202
rect 34692 2164 34744 2173
rect 34692 2130 34701 2164
rect 34701 2130 34735 2164
rect 34735 2130 34744 2164
rect 34692 2121 34744 2130
rect 34692 2092 34744 2109
rect 34692 2058 34701 2092
rect 34701 2058 34735 2092
rect 34735 2058 34744 2092
rect 34692 2057 34744 2058
rect 34692 2020 34744 2045
rect 34692 1993 34701 2020
rect 34701 1993 34735 2020
rect 34735 1993 34744 2020
rect 34692 1948 34744 1981
rect 34692 1929 34701 1948
rect 34701 1929 34735 1948
rect 34735 1929 34744 1948
rect 34692 1914 34701 1917
rect 34701 1914 34735 1917
rect 34735 1914 34744 1917
rect 34692 1876 34744 1914
rect 34692 1865 34701 1876
rect 34701 1865 34735 1876
rect 34735 1865 34744 1876
rect 34692 1842 34701 1853
rect 34701 1842 34735 1853
rect 34735 1842 34744 1853
rect 34692 1804 34744 1842
rect 34692 1801 34701 1804
rect 34701 1801 34735 1804
rect 34735 1801 34744 1804
rect 34692 1770 34701 1789
rect 34701 1770 34735 1789
rect 34735 1770 34744 1789
rect 34692 1737 34744 1770
rect 34692 1698 34701 1725
rect 34701 1698 34735 1725
rect 34735 1698 34744 1725
rect 34692 1673 34744 1698
rect 34692 1660 34744 1661
rect 34692 1626 34701 1660
rect 34701 1626 34735 1660
rect 34735 1626 34744 1660
rect 34692 1609 34744 1626
rect 34692 1588 34744 1597
rect 34692 1554 34701 1588
rect 34701 1554 34735 1588
rect 34735 1554 34744 1588
rect 34692 1545 34744 1554
rect 34692 1516 34744 1533
rect 34692 1482 34701 1516
rect 34701 1482 34735 1516
rect 34735 1482 34744 1516
rect 34692 1481 34744 1482
rect 34692 1444 34744 1469
rect 34692 1417 34701 1444
rect 34701 1417 34735 1444
rect 34735 1417 34744 1444
rect 34692 1372 34744 1405
rect 34692 1353 34701 1372
rect 34701 1353 34735 1372
rect 34735 1353 34744 1372
rect 34692 1338 34701 1341
rect 34701 1338 34735 1341
rect 34735 1338 34744 1341
rect 34692 1300 34744 1338
rect 34692 1289 34701 1300
rect 34701 1289 34735 1300
rect 34735 1289 34744 1300
rect 34692 1266 34701 1277
rect 34701 1266 34735 1277
rect 34735 1266 34744 1277
rect 34692 1228 34744 1266
rect 34692 1225 34701 1228
rect 34701 1225 34735 1228
rect 34735 1225 34744 1228
rect 34692 1194 34701 1213
rect 34701 1194 34735 1213
rect 34735 1194 34744 1213
rect 34692 1161 34744 1194
rect 34788 3100 34840 3133
rect 34788 3081 34797 3100
rect 34797 3081 34831 3100
rect 34831 3081 34840 3100
rect 34788 3066 34797 3069
rect 34797 3066 34831 3069
rect 34831 3066 34840 3069
rect 34788 3028 34840 3066
rect 34788 3017 34797 3028
rect 34797 3017 34831 3028
rect 34831 3017 34840 3028
rect 34788 2994 34797 3005
rect 34797 2994 34831 3005
rect 34831 2994 34840 3005
rect 34788 2956 34840 2994
rect 34788 2953 34797 2956
rect 34797 2953 34831 2956
rect 34831 2953 34840 2956
rect 34788 2922 34797 2941
rect 34797 2922 34831 2941
rect 34831 2922 34840 2941
rect 34788 2889 34840 2922
rect 34788 2850 34797 2877
rect 34797 2850 34831 2877
rect 34831 2850 34840 2877
rect 34788 2825 34840 2850
rect 34788 2812 34840 2813
rect 34788 2778 34797 2812
rect 34797 2778 34831 2812
rect 34831 2778 34840 2812
rect 34788 2761 34840 2778
rect 34788 2740 34840 2749
rect 34788 2706 34797 2740
rect 34797 2706 34831 2740
rect 34831 2706 34840 2740
rect 34788 2697 34840 2706
rect 34788 2668 34840 2685
rect 34788 2634 34797 2668
rect 34797 2634 34831 2668
rect 34831 2634 34840 2668
rect 34788 2633 34840 2634
rect 34788 2596 34840 2621
rect 34788 2569 34797 2596
rect 34797 2569 34831 2596
rect 34831 2569 34840 2596
rect 34788 2524 34840 2557
rect 34788 2505 34797 2524
rect 34797 2505 34831 2524
rect 34831 2505 34840 2524
rect 34788 2490 34797 2493
rect 34797 2490 34831 2493
rect 34831 2490 34840 2493
rect 34788 2452 34840 2490
rect 34788 2441 34797 2452
rect 34797 2441 34831 2452
rect 34831 2441 34840 2452
rect 34788 2418 34797 2429
rect 34797 2418 34831 2429
rect 34831 2418 34840 2429
rect 34788 2380 34840 2418
rect 34788 2377 34797 2380
rect 34797 2377 34831 2380
rect 34831 2377 34840 2380
rect 34788 2346 34797 2365
rect 34797 2346 34831 2365
rect 34831 2346 34840 2365
rect 34788 2313 34840 2346
rect 34788 2274 34797 2301
rect 34797 2274 34831 2301
rect 34831 2274 34840 2301
rect 34788 2249 34840 2274
rect 34788 2236 34840 2237
rect 34788 2202 34797 2236
rect 34797 2202 34831 2236
rect 34831 2202 34840 2236
rect 34788 2185 34840 2202
rect 34788 2164 34840 2173
rect 34788 2130 34797 2164
rect 34797 2130 34831 2164
rect 34831 2130 34840 2164
rect 34788 2121 34840 2130
rect 34788 2092 34840 2109
rect 34788 2058 34797 2092
rect 34797 2058 34831 2092
rect 34831 2058 34840 2092
rect 34788 2057 34840 2058
rect 34788 2020 34840 2045
rect 34788 1993 34797 2020
rect 34797 1993 34831 2020
rect 34831 1993 34840 2020
rect 34788 1948 34840 1981
rect 34788 1929 34797 1948
rect 34797 1929 34831 1948
rect 34831 1929 34840 1948
rect 34788 1914 34797 1917
rect 34797 1914 34831 1917
rect 34831 1914 34840 1917
rect 34788 1876 34840 1914
rect 34788 1865 34797 1876
rect 34797 1865 34831 1876
rect 34831 1865 34840 1876
rect 34788 1842 34797 1853
rect 34797 1842 34831 1853
rect 34831 1842 34840 1853
rect 34788 1804 34840 1842
rect 34788 1801 34797 1804
rect 34797 1801 34831 1804
rect 34831 1801 34840 1804
rect 34788 1770 34797 1789
rect 34797 1770 34831 1789
rect 34831 1770 34840 1789
rect 34788 1737 34840 1770
rect 34788 1698 34797 1725
rect 34797 1698 34831 1725
rect 34831 1698 34840 1725
rect 34788 1673 34840 1698
rect 34788 1660 34840 1661
rect 34788 1626 34797 1660
rect 34797 1626 34831 1660
rect 34831 1626 34840 1660
rect 34788 1609 34840 1626
rect 34788 1588 34840 1597
rect 34788 1554 34797 1588
rect 34797 1554 34831 1588
rect 34831 1554 34840 1588
rect 34788 1545 34840 1554
rect 34788 1516 34840 1533
rect 34788 1482 34797 1516
rect 34797 1482 34831 1516
rect 34831 1482 34840 1516
rect 34788 1481 34840 1482
rect 34788 1444 34840 1469
rect 34788 1417 34797 1444
rect 34797 1417 34831 1444
rect 34831 1417 34840 1444
rect 34788 1372 34840 1405
rect 34788 1353 34797 1372
rect 34797 1353 34831 1372
rect 34831 1353 34840 1372
rect 34788 1338 34797 1341
rect 34797 1338 34831 1341
rect 34831 1338 34840 1341
rect 34788 1300 34840 1338
rect 34788 1289 34797 1300
rect 34797 1289 34831 1300
rect 34831 1289 34840 1300
rect 34788 1266 34797 1277
rect 34797 1266 34831 1277
rect 34831 1266 34840 1277
rect 34788 1228 34840 1266
rect 34788 1225 34797 1228
rect 34797 1225 34831 1228
rect 34831 1225 34840 1228
rect 34788 1194 34797 1213
rect 34797 1194 34831 1213
rect 34831 1194 34840 1213
rect 34788 1161 34840 1194
rect 34884 3100 34936 3133
rect 34884 3081 34893 3100
rect 34893 3081 34927 3100
rect 34927 3081 34936 3100
rect 34884 3066 34893 3069
rect 34893 3066 34927 3069
rect 34927 3066 34936 3069
rect 34884 3028 34936 3066
rect 34884 3017 34893 3028
rect 34893 3017 34927 3028
rect 34927 3017 34936 3028
rect 34884 2994 34893 3005
rect 34893 2994 34927 3005
rect 34927 2994 34936 3005
rect 34884 2956 34936 2994
rect 34884 2953 34893 2956
rect 34893 2953 34927 2956
rect 34927 2953 34936 2956
rect 34884 2922 34893 2941
rect 34893 2922 34927 2941
rect 34927 2922 34936 2941
rect 34884 2889 34936 2922
rect 34884 2850 34893 2877
rect 34893 2850 34927 2877
rect 34927 2850 34936 2877
rect 34884 2825 34936 2850
rect 34884 2812 34936 2813
rect 34884 2778 34893 2812
rect 34893 2778 34927 2812
rect 34927 2778 34936 2812
rect 34884 2761 34936 2778
rect 34884 2740 34936 2749
rect 34884 2706 34893 2740
rect 34893 2706 34927 2740
rect 34927 2706 34936 2740
rect 34884 2697 34936 2706
rect 34884 2668 34936 2685
rect 34884 2634 34893 2668
rect 34893 2634 34927 2668
rect 34927 2634 34936 2668
rect 34884 2633 34936 2634
rect 34884 2596 34936 2621
rect 34884 2569 34893 2596
rect 34893 2569 34927 2596
rect 34927 2569 34936 2596
rect 34884 2524 34936 2557
rect 34884 2505 34893 2524
rect 34893 2505 34927 2524
rect 34927 2505 34936 2524
rect 34884 2490 34893 2493
rect 34893 2490 34927 2493
rect 34927 2490 34936 2493
rect 34884 2452 34936 2490
rect 34884 2441 34893 2452
rect 34893 2441 34927 2452
rect 34927 2441 34936 2452
rect 34884 2418 34893 2429
rect 34893 2418 34927 2429
rect 34927 2418 34936 2429
rect 34884 2380 34936 2418
rect 34884 2377 34893 2380
rect 34893 2377 34927 2380
rect 34927 2377 34936 2380
rect 34884 2346 34893 2365
rect 34893 2346 34927 2365
rect 34927 2346 34936 2365
rect 34884 2313 34936 2346
rect 34884 2274 34893 2301
rect 34893 2274 34927 2301
rect 34927 2274 34936 2301
rect 34884 2249 34936 2274
rect 34884 2236 34936 2237
rect 34884 2202 34893 2236
rect 34893 2202 34927 2236
rect 34927 2202 34936 2236
rect 34884 2185 34936 2202
rect 34884 2164 34936 2173
rect 34884 2130 34893 2164
rect 34893 2130 34927 2164
rect 34927 2130 34936 2164
rect 34884 2121 34936 2130
rect 34884 2092 34936 2109
rect 34884 2058 34893 2092
rect 34893 2058 34927 2092
rect 34927 2058 34936 2092
rect 34884 2057 34936 2058
rect 34884 2020 34936 2045
rect 34884 1993 34893 2020
rect 34893 1993 34927 2020
rect 34927 1993 34936 2020
rect 34884 1948 34936 1981
rect 34884 1929 34893 1948
rect 34893 1929 34927 1948
rect 34927 1929 34936 1948
rect 34884 1914 34893 1917
rect 34893 1914 34927 1917
rect 34927 1914 34936 1917
rect 34884 1876 34936 1914
rect 34884 1865 34893 1876
rect 34893 1865 34927 1876
rect 34927 1865 34936 1876
rect 34884 1842 34893 1853
rect 34893 1842 34927 1853
rect 34927 1842 34936 1853
rect 34884 1804 34936 1842
rect 34884 1801 34893 1804
rect 34893 1801 34927 1804
rect 34927 1801 34936 1804
rect 34884 1770 34893 1789
rect 34893 1770 34927 1789
rect 34927 1770 34936 1789
rect 34884 1737 34936 1770
rect 34884 1698 34893 1725
rect 34893 1698 34927 1725
rect 34927 1698 34936 1725
rect 34884 1673 34936 1698
rect 34884 1660 34936 1661
rect 34884 1626 34893 1660
rect 34893 1626 34927 1660
rect 34927 1626 34936 1660
rect 34884 1609 34936 1626
rect 34884 1588 34936 1597
rect 34884 1554 34893 1588
rect 34893 1554 34927 1588
rect 34927 1554 34936 1588
rect 34884 1545 34936 1554
rect 34884 1516 34936 1533
rect 34884 1482 34893 1516
rect 34893 1482 34927 1516
rect 34927 1482 34936 1516
rect 34884 1481 34936 1482
rect 34884 1444 34936 1469
rect 34884 1417 34893 1444
rect 34893 1417 34927 1444
rect 34927 1417 34936 1444
rect 34884 1372 34936 1405
rect 34884 1353 34893 1372
rect 34893 1353 34927 1372
rect 34927 1353 34936 1372
rect 34884 1338 34893 1341
rect 34893 1338 34927 1341
rect 34927 1338 34936 1341
rect 34884 1300 34936 1338
rect 34884 1289 34893 1300
rect 34893 1289 34927 1300
rect 34927 1289 34936 1300
rect 34884 1266 34893 1277
rect 34893 1266 34927 1277
rect 34927 1266 34936 1277
rect 34884 1228 34936 1266
rect 34884 1225 34893 1228
rect 34893 1225 34927 1228
rect 34927 1225 34936 1228
rect 34884 1194 34893 1213
rect 34893 1194 34927 1213
rect 34927 1194 34936 1213
rect 34884 1161 34936 1194
rect 34980 3100 35032 3133
rect 34980 3081 34989 3100
rect 34989 3081 35023 3100
rect 35023 3081 35032 3100
rect 34980 3066 34989 3069
rect 34989 3066 35023 3069
rect 35023 3066 35032 3069
rect 34980 3028 35032 3066
rect 34980 3017 34989 3028
rect 34989 3017 35023 3028
rect 35023 3017 35032 3028
rect 34980 2994 34989 3005
rect 34989 2994 35023 3005
rect 35023 2994 35032 3005
rect 34980 2956 35032 2994
rect 34980 2953 34989 2956
rect 34989 2953 35023 2956
rect 35023 2953 35032 2956
rect 34980 2922 34989 2941
rect 34989 2922 35023 2941
rect 35023 2922 35032 2941
rect 34980 2889 35032 2922
rect 34980 2850 34989 2877
rect 34989 2850 35023 2877
rect 35023 2850 35032 2877
rect 34980 2825 35032 2850
rect 34980 2812 35032 2813
rect 34980 2778 34989 2812
rect 34989 2778 35023 2812
rect 35023 2778 35032 2812
rect 34980 2761 35032 2778
rect 34980 2740 35032 2749
rect 34980 2706 34989 2740
rect 34989 2706 35023 2740
rect 35023 2706 35032 2740
rect 34980 2697 35032 2706
rect 34980 2668 35032 2685
rect 34980 2634 34989 2668
rect 34989 2634 35023 2668
rect 35023 2634 35032 2668
rect 34980 2633 35032 2634
rect 34980 2596 35032 2621
rect 34980 2569 34989 2596
rect 34989 2569 35023 2596
rect 35023 2569 35032 2596
rect 34980 2524 35032 2557
rect 34980 2505 34989 2524
rect 34989 2505 35023 2524
rect 35023 2505 35032 2524
rect 34980 2490 34989 2493
rect 34989 2490 35023 2493
rect 35023 2490 35032 2493
rect 34980 2452 35032 2490
rect 34980 2441 34989 2452
rect 34989 2441 35023 2452
rect 35023 2441 35032 2452
rect 34980 2418 34989 2429
rect 34989 2418 35023 2429
rect 35023 2418 35032 2429
rect 34980 2380 35032 2418
rect 34980 2377 34989 2380
rect 34989 2377 35023 2380
rect 35023 2377 35032 2380
rect 34980 2346 34989 2365
rect 34989 2346 35023 2365
rect 35023 2346 35032 2365
rect 34980 2313 35032 2346
rect 34980 2274 34989 2301
rect 34989 2274 35023 2301
rect 35023 2274 35032 2301
rect 34980 2249 35032 2274
rect 34980 2236 35032 2237
rect 34980 2202 34989 2236
rect 34989 2202 35023 2236
rect 35023 2202 35032 2236
rect 34980 2185 35032 2202
rect 34980 2164 35032 2173
rect 34980 2130 34989 2164
rect 34989 2130 35023 2164
rect 35023 2130 35032 2164
rect 34980 2121 35032 2130
rect 34980 2092 35032 2109
rect 34980 2058 34989 2092
rect 34989 2058 35023 2092
rect 35023 2058 35032 2092
rect 34980 2057 35032 2058
rect 34980 2020 35032 2045
rect 34980 1993 34989 2020
rect 34989 1993 35023 2020
rect 35023 1993 35032 2020
rect 34980 1948 35032 1981
rect 34980 1929 34989 1948
rect 34989 1929 35023 1948
rect 35023 1929 35032 1948
rect 34980 1914 34989 1917
rect 34989 1914 35023 1917
rect 35023 1914 35032 1917
rect 34980 1876 35032 1914
rect 34980 1865 34989 1876
rect 34989 1865 35023 1876
rect 35023 1865 35032 1876
rect 34980 1842 34989 1853
rect 34989 1842 35023 1853
rect 35023 1842 35032 1853
rect 34980 1804 35032 1842
rect 34980 1801 34989 1804
rect 34989 1801 35023 1804
rect 35023 1801 35032 1804
rect 34980 1770 34989 1789
rect 34989 1770 35023 1789
rect 35023 1770 35032 1789
rect 34980 1737 35032 1770
rect 34980 1698 34989 1725
rect 34989 1698 35023 1725
rect 35023 1698 35032 1725
rect 34980 1673 35032 1698
rect 34980 1660 35032 1661
rect 34980 1626 34989 1660
rect 34989 1626 35023 1660
rect 35023 1626 35032 1660
rect 34980 1609 35032 1626
rect 34980 1588 35032 1597
rect 34980 1554 34989 1588
rect 34989 1554 35023 1588
rect 35023 1554 35032 1588
rect 34980 1545 35032 1554
rect 34980 1516 35032 1533
rect 34980 1482 34989 1516
rect 34989 1482 35023 1516
rect 35023 1482 35032 1516
rect 34980 1481 35032 1482
rect 34980 1444 35032 1469
rect 34980 1417 34989 1444
rect 34989 1417 35023 1444
rect 35023 1417 35032 1444
rect 34980 1372 35032 1405
rect 34980 1353 34989 1372
rect 34989 1353 35023 1372
rect 35023 1353 35032 1372
rect 34980 1338 34989 1341
rect 34989 1338 35023 1341
rect 35023 1338 35032 1341
rect 34980 1300 35032 1338
rect 34980 1289 34989 1300
rect 34989 1289 35023 1300
rect 35023 1289 35032 1300
rect 34980 1266 34989 1277
rect 34989 1266 35023 1277
rect 35023 1266 35032 1277
rect 34980 1228 35032 1266
rect 34980 1225 34989 1228
rect 34989 1225 35023 1228
rect 35023 1225 35032 1228
rect 34980 1194 34989 1213
rect 34989 1194 35023 1213
rect 35023 1194 35032 1213
rect 34980 1161 35032 1194
rect 35076 3100 35128 3133
rect 35076 3081 35085 3100
rect 35085 3081 35119 3100
rect 35119 3081 35128 3100
rect 35076 3066 35085 3069
rect 35085 3066 35119 3069
rect 35119 3066 35128 3069
rect 35076 3028 35128 3066
rect 35076 3017 35085 3028
rect 35085 3017 35119 3028
rect 35119 3017 35128 3028
rect 35076 2994 35085 3005
rect 35085 2994 35119 3005
rect 35119 2994 35128 3005
rect 35076 2956 35128 2994
rect 35076 2953 35085 2956
rect 35085 2953 35119 2956
rect 35119 2953 35128 2956
rect 35076 2922 35085 2941
rect 35085 2922 35119 2941
rect 35119 2922 35128 2941
rect 35076 2889 35128 2922
rect 35076 2850 35085 2877
rect 35085 2850 35119 2877
rect 35119 2850 35128 2877
rect 35076 2825 35128 2850
rect 35076 2812 35128 2813
rect 35076 2778 35085 2812
rect 35085 2778 35119 2812
rect 35119 2778 35128 2812
rect 35076 2761 35128 2778
rect 35076 2740 35128 2749
rect 35076 2706 35085 2740
rect 35085 2706 35119 2740
rect 35119 2706 35128 2740
rect 35076 2697 35128 2706
rect 35076 2668 35128 2685
rect 35076 2634 35085 2668
rect 35085 2634 35119 2668
rect 35119 2634 35128 2668
rect 35076 2633 35128 2634
rect 35076 2596 35128 2621
rect 35076 2569 35085 2596
rect 35085 2569 35119 2596
rect 35119 2569 35128 2596
rect 35076 2524 35128 2557
rect 35076 2505 35085 2524
rect 35085 2505 35119 2524
rect 35119 2505 35128 2524
rect 35076 2490 35085 2493
rect 35085 2490 35119 2493
rect 35119 2490 35128 2493
rect 35076 2452 35128 2490
rect 35076 2441 35085 2452
rect 35085 2441 35119 2452
rect 35119 2441 35128 2452
rect 35076 2418 35085 2429
rect 35085 2418 35119 2429
rect 35119 2418 35128 2429
rect 35076 2380 35128 2418
rect 35076 2377 35085 2380
rect 35085 2377 35119 2380
rect 35119 2377 35128 2380
rect 35076 2346 35085 2365
rect 35085 2346 35119 2365
rect 35119 2346 35128 2365
rect 35076 2313 35128 2346
rect 35076 2274 35085 2301
rect 35085 2274 35119 2301
rect 35119 2274 35128 2301
rect 35076 2249 35128 2274
rect 35076 2236 35128 2237
rect 35076 2202 35085 2236
rect 35085 2202 35119 2236
rect 35119 2202 35128 2236
rect 35076 2185 35128 2202
rect 35076 2164 35128 2173
rect 35076 2130 35085 2164
rect 35085 2130 35119 2164
rect 35119 2130 35128 2164
rect 35076 2121 35128 2130
rect 35076 2092 35128 2109
rect 35076 2058 35085 2092
rect 35085 2058 35119 2092
rect 35119 2058 35128 2092
rect 35076 2057 35128 2058
rect 35076 2020 35128 2045
rect 35076 1993 35085 2020
rect 35085 1993 35119 2020
rect 35119 1993 35128 2020
rect 35076 1948 35128 1981
rect 35076 1929 35085 1948
rect 35085 1929 35119 1948
rect 35119 1929 35128 1948
rect 35076 1914 35085 1917
rect 35085 1914 35119 1917
rect 35119 1914 35128 1917
rect 35076 1876 35128 1914
rect 35076 1865 35085 1876
rect 35085 1865 35119 1876
rect 35119 1865 35128 1876
rect 35076 1842 35085 1853
rect 35085 1842 35119 1853
rect 35119 1842 35128 1853
rect 35076 1804 35128 1842
rect 35076 1801 35085 1804
rect 35085 1801 35119 1804
rect 35119 1801 35128 1804
rect 35076 1770 35085 1789
rect 35085 1770 35119 1789
rect 35119 1770 35128 1789
rect 35076 1737 35128 1770
rect 35076 1698 35085 1725
rect 35085 1698 35119 1725
rect 35119 1698 35128 1725
rect 35076 1673 35128 1698
rect 35076 1660 35128 1661
rect 35076 1626 35085 1660
rect 35085 1626 35119 1660
rect 35119 1626 35128 1660
rect 35076 1609 35128 1626
rect 35076 1588 35128 1597
rect 35076 1554 35085 1588
rect 35085 1554 35119 1588
rect 35119 1554 35128 1588
rect 35076 1545 35128 1554
rect 35076 1516 35128 1533
rect 35076 1482 35085 1516
rect 35085 1482 35119 1516
rect 35119 1482 35128 1516
rect 35076 1481 35128 1482
rect 35076 1444 35128 1469
rect 35076 1417 35085 1444
rect 35085 1417 35119 1444
rect 35119 1417 35128 1444
rect 35076 1372 35128 1405
rect 35076 1353 35085 1372
rect 35085 1353 35119 1372
rect 35119 1353 35128 1372
rect 35076 1338 35085 1341
rect 35085 1338 35119 1341
rect 35119 1338 35128 1341
rect 35076 1300 35128 1338
rect 35076 1289 35085 1300
rect 35085 1289 35119 1300
rect 35119 1289 35128 1300
rect 35076 1266 35085 1277
rect 35085 1266 35119 1277
rect 35119 1266 35128 1277
rect 35076 1228 35128 1266
rect 35076 1225 35085 1228
rect 35085 1225 35119 1228
rect 35119 1225 35128 1228
rect 35076 1194 35085 1213
rect 35085 1194 35119 1213
rect 35119 1194 35128 1213
rect 35076 1161 35128 1194
rect 35172 3100 35224 3133
rect 35172 3081 35181 3100
rect 35181 3081 35215 3100
rect 35215 3081 35224 3100
rect 35172 3066 35181 3069
rect 35181 3066 35215 3069
rect 35215 3066 35224 3069
rect 35172 3028 35224 3066
rect 35172 3017 35181 3028
rect 35181 3017 35215 3028
rect 35215 3017 35224 3028
rect 35172 2994 35181 3005
rect 35181 2994 35215 3005
rect 35215 2994 35224 3005
rect 35172 2956 35224 2994
rect 35172 2953 35181 2956
rect 35181 2953 35215 2956
rect 35215 2953 35224 2956
rect 35172 2922 35181 2941
rect 35181 2922 35215 2941
rect 35215 2922 35224 2941
rect 35172 2889 35224 2922
rect 35172 2850 35181 2877
rect 35181 2850 35215 2877
rect 35215 2850 35224 2877
rect 35172 2825 35224 2850
rect 35172 2812 35224 2813
rect 35172 2778 35181 2812
rect 35181 2778 35215 2812
rect 35215 2778 35224 2812
rect 35172 2761 35224 2778
rect 35172 2740 35224 2749
rect 35172 2706 35181 2740
rect 35181 2706 35215 2740
rect 35215 2706 35224 2740
rect 35172 2697 35224 2706
rect 35172 2668 35224 2685
rect 35172 2634 35181 2668
rect 35181 2634 35215 2668
rect 35215 2634 35224 2668
rect 35172 2633 35224 2634
rect 35172 2596 35224 2621
rect 35172 2569 35181 2596
rect 35181 2569 35215 2596
rect 35215 2569 35224 2596
rect 35172 2524 35224 2557
rect 35172 2505 35181 2524
rect 35181 2505 35215 2524
rect 35215 2505 35224 2524
rect 35172 2490 35181 2493
rect 35181 2490 35215 2493
rect 35215 2490 35224 2493
rect 35172 2452 35224 2490
rect 35172 2441 35181 2452
rect 35181 2441 35215 2452
rect 35215 2441 35224 2452
rect 35172 2418 35181 2429
rect 35181 2418 35215 2429
rect 35215 2418 35224 2429
rect 35172 2380 35224 2418
rect 35172 2377 35181 2380
rect 35181 2377 35215 2380
rect 35215 2377 35224 2380
rect 35172 2346 35181 2365
rect 35181 2346 35215 2365
rect 35215 2346 35224 2365
rect 35172 2313 35224 2346
rect 35172 2274 35181 2301
rect 35181 2274 35215 2301
rect 35215 2274 35224 2301
rect 35172 2249 35224 2274
rect 35172 2236 35224 2237
rect 35172 2202 35181 2236
rect 35181 2202 35215 2236
rect 35215 2202 35224 2236
rect 35172 2185 35224 2202
rect 35172 2164 35224 2173
rect 35172 2130 35181 2164
rect 35181 2130 35215 2164
rect 35215 2130 35224 2164
rect 35172 2121 35224 2130
rect 35172 2092 35224 2109
rect 35172 2058 35181 2092
rect 35181 2058 35215 2092
rect 35215 2058 35224 2092
rect 35172 2057 35224 2058
rect 35172 2020 35224 2045
rect 35172 1993 35181 2020
rect 35181 1993 35215 2020
rect 35215 1993 35224 2020
rect 35172 1948 35224 1981
rect 35172 1929 35181 1948
rect 35181 1929 35215 1948
rect 35215 1929 35224 1948
rect 35172 1914 35181 1917
rect 35181 1914 35215 1917
rect 35215 1914 35224 1917
rect 35172 1876 35224 1914
rect 35172 1865 35181 1876
rect 35181 1865 35215 1876
rect 35215 1865 35224 1876
rect 35172 1842 35181 1853
rect 35181 1842 35215 1853
rect 35215 1842 35224 1853
rect 35172 1804 35224 1842
rect 35172 1801 35181 1804
rect 35181 1801 35215 1804
rect 35215 1801 35224 1804
rect 35172 1770 35181 1789
rect 35181 1770 35215 1789
rect 35215 1770 35224 1789
rect 35172 1737 35224 1770
rect 35172 1698 35181 1725
rect 35181 1698 35215 1725
rect 35215 1698 35224 1725
rect 35172 1673 35224 1698
rect 35172 1660 35224 1661
rect 35172 1626 35181 1660
rect 35181 1626 35215 1660
rect 35215 1626 35224 1660
rect 35172 1609 35224 1626
rect 35172 1588 35224 1597
rect 35172 1554 35181 1588
rect 35181 1554 35215 1588
rect 35215 1554 35224 1588
rect 35172 1545 35224 1554
rect 35172 1516 35224 1533
rect 35172 1482 35181 1516
rect 35181 1482 35215 1516
rect 35215 1482 35224 1516
rect 35172 1481 35224 1482
rect 35172 1444 35224 1469
rect 35172 1417 35181 1444
rect 35181 1417 35215 1444
rect 35215 1417 35224 1444
rect 35172 1372 35224 1405
rect 35172 1353 35181 1372
rect 35181 1353 35215 1372
rect 35215 1353 35224 1372
rect 35172 1338 35181 1341
rect 35181 1338 35215 1341
rect 35215 1338 35224 1341
rect 35172 1300 35224 1338
rect 35172 1289 35181 1300
rect 35181 1289 35215 1300
rect 35215 1289 35224 1300
rect 35172 1266 35181 1277
rect 35181 1266 35215 1277
rect 35215 1266 35224 1277
rect 35172 1228 35224 1266
rect 35172 1225 35181 1228
rect 35181 1225 35215 1228
rect 35215 1225 35224 1228
rect 35172 1194 35181 1213
rect 35181 1194 35215 1213
rect 35215 1194 35224 1213
rect 35172 1161 35224 1194
rect 35268 3100 35320 3133
rect 35268 3081 35277 3100
rect 35277 3081 35311 3100
rect 35311 3081 35320 3100
rect 35268 3066 35277 3069
rect 35277 3066 35311 3069
rect 35311 3066 35320 3069
rect 35268 3028 35320 3066
rect 35268 3017 35277 3028
rect 35277 3017 35311 3028
rect 35311 3017 35320 3028
rect 35268 2994 35277 3005
rect 35277 2994 35311 3005
rect 35311 2994 35320 3005
rect 35268 2956 35320 2994
rect 35268 2953 35277 2956
rect 35277 2953 35311 2956
rect 35311 2953 35320 2956
rect 35268 2922 35277 2941
rect 35277 2922 35311 2941
rect 35311 2922 35320 2941
rect 35268 2889 35320 2922
rect 35268 2850 35277 2877
rect 35277 2850 35311 2877
rect 35311 2850 35320 2877
rect 35268 2825 35320 2850
rect 35268 2812 35320 2813
rect 35268 2778 35277 2812
rect 35277 2778 35311 2812
rect 35311 2778 35320 2812
rect 35268 2761 35320 2778
rect 35268 2740 35320 2749
rect 35268 2706 35277 2740
rect 35277 2706 35311 2740
rect 35311 2706 35320 2740
rect 35268 2697 35320 2706
rect 35268 2668 35320 2685
rect 35268 2634 35277 2668
rect 35277 2634 35311 2668
rect 35311 2634 35320 2668
rect 35268 2633 35320 2634
rect 35268 2596 35320 2621
rect 35268 2569 35277 2596
rect 35277 2569 35311 2596
rect 35311 2569 35320 2596
rect 35268 2524 35320 2557
rect 35268 2505 35277 2524
rect 35277 2505 35311 2524
rect 35311 2505 35320 2524
rect 35268 2490 35277 2493
rect 35277 2490 35311 2493
rect 35311 2490 35320 2493
rect 35268 2452 35320 2490
rect 35268 2441 35277 2452
rect 35277 2441 35311 2452
rect 35311 2441 35320 2452
rect 35268 2418 35277 2429
rect 35277 2418 35311 2429
rect 35311 2418 35320 2429
rect 35268 2380 35320 2418
rect 35268 2377 35277 2380
rect 35277 2377 35311 2380
rect 35311 2377 35320 2380
rect 35268 2346 35277 2365
rect 35277 2346 35311 2365
rect 35311 2346 35320 2365
rect 35268 2313 35320 2346
rect 35268 2274 35277 2301
rect 35277 2274 35311 2301
rect 35311 2274 35320 2301
rect 35268 2249 35320 2274
rect 35268 2236 35320 2237
rect 35268 2202 35277 2236
rect 35277 2202 35311 2236
rect 35311 2202 35320 2236
rect 35268 2185 35320 2202
rect 35268 2164 35320 2173
rect 35268 2130 35277 2164
rect 35277 2130 35311 2164
rect 35311 2130 35320 2164
rect 35268 2121 35320 2130
rect 35268 2092 35320 2109
rect 35268 2058 35277 2092
rect 35277 2058 35311 2092
rect 35311 2058 35320 2092
rect 35268 2057 35320 2058
rect 35268 2020 35320 2045
rect 35268 1993 35277 2020
rect 35277 1993 35311 2020
rect 35311 1993 35320 2020
rect 35268 1948 35320 1981
rect 35268 1929 35277 1948
rect 35277 1929 35311 1948
rect 35311 1929 35320 1948
rect 35268 1914 35277 1917
rect 35277 1914 35311 1917
rect 35311 1914 35320 1917
rect 35268 1876 35320 1914
rect 35268 1865 35277 1876
rect 35277 1865 35311 1876
rect 35311 1865 35320 1876
rect 35268 1842 35277 1853
rect 35277 1842 35311 1853
rect 35311 1842 35320 1853
rect 35268 1804 35320 1842
rect 35268 1801 35277 1804
rect 35277 1801 35311 1804
rect 35311 1801 35320 1804
rect 35268 1770 35277 1789
rect 35277 1770 35311 1789
rect 35311 1770 35320 1789
rect 35268 1737 35320 1770
rect 35268 1698 35277 1725
rect 35277 1698 35311 1725
rect 35311 1698 35320 1725
rect 35268 1673 35320 1698
rect 35268 1660 35320 1661
rect 35268 1626 35277 1660
rect 35277 1626 35311 1660
rect 35311 1626 35320 1660
rect 35268 1609 35320 1626
rect 35268 1588 35320 1597
rect 35268 1554 35277 1588
rect 35277 1554 35311 1588
rect 35311 1554 35320 1588
rect 35268 1545 35320 1554
rect 35268 1516 35320 1533
rect 35268 1482 35277 1516
rect 35277 1482 35311 1516
rect 35311 1482 35320 1516
rect 35268 1481 35320 1482
rect 35268 1444 35320 1469
rect 35268 1417 35277 1444
rect 35277 1417 35311 1444
rect 35311 1417 35320 1444
rect 35268 1372 35320 1405
rect 35268 1353 35277 1372
rect 35277 1353 35311 1372
rect 35311 1353 35320 1372
rect 35268 1338 35277 1341
rect 35277 1338 35311 1341
rect 35311 1338 35320 1341
rect 35268 1300 35320 1338
rect 35268 1289 35277 1300
rect 35277 1289 35311 1300
rect 35311 1289 35320 1300
rect 35268 1266 35277 1277
rect 35277 1266 35311 1277
rect 35311 1266 35320 1277
rect 35268 1228 35320 1266
rect 35268 1225 35277 1228
rect 35277 1225 35311 1228
rect 35311 1225 35320 1228
rect 35268 1194 35277 1213
rect 35277 1194 35311 1213
rect 35311 1194 35320 1213
rect 35268 1161 35320 1194
rect 35364 3100 35416 3133
rect 35364 3081 35373 3100
rect 35373 3081 35407 3100
rect 35407 3081 35416 3100
rect 35364 3066 35373 3069
rect 35373 3066 35407 3069
rect 35407 3066 35416 3069
rect 35364 3028 35416 3066
rect 35364 3017 35373 3028
rect 35373 3017 35407 3028
rect 35407 3017 35416 3028
rect 35364 2994 35373 3005
rect 35373 2994 35407 3005
rect 35407 2994 35416 3005
rect 35364 2956 35416 2994
rect 35364 2953 35373 2956
rect 35373 2953 35407 2956
rect 35407 2953 35416 2956
rect 35364 2922 35373 2941
rect 35373 2922 35407 2941
rect 35407 2922 35416 2941
rect 35364 2889 35416 2922
rect 35364 2850 35373 2877
rect 35373 2850 35407 2877
rect 35407 2850 35416 2877
rect 35364 2825 35416 2850
rect 35364 2812 35416 2813
rect 35364 2778 35373 2812
rect 35373 2778 35407 2812
rect 35407 2778 35416 2812
rect 35364 2761 35416 2778
rect 35364 2740 35416 2749
rect 35364 2706 35373 2740
rect 35373 2706 35407 2740
rect 35407 2706 35416 2740
rect 35364 2697 35416 2706
rect 35364 2668 35416 2685
rect 35364 2634 35373 2668
rect 35373 2634 35407 2668
rect 35407 2634 35416 2668
rect 35364 2633 35416 2634
rect 35364 2596 35416 2621
rect 35364 2569 35373 2596
rect 35373 2569 35407 2596
rect 35407 2569 35416 2596
rect 35364 2524 35416 2557
rect 35364 2505 35373 2524
rect 35373 2505 35407 2524
rect 35407 2505 35416 2524
rect 35364 2490 35373 2493
rect 35373 2490 35407 2493
rect 35407 2490 35416 2493
rect 35364 2452 35416 2490
rect 35364 2441 35373 2452
rect 35373 2441 35407 2452
rect 35407 2441 35416 2452
rect 35364 2418 35373 2429
rect 35373 2418 35407 2429
rect 35407 2418 35416 2429
rect 35364 2380 35416 2418
rect 35364 2377 35373 2380
rect 35373 2377 35407 2380
rect 35407 2377 35416 2380
rect 35364 2346 35373 2365
rect 35373 2346 35407 2365
rect 35407 2346 35416 2365
rect 35364 2313 35416 2346
rect 35364 2274 35373 2301
rect 35373 2274 35407 2301
rect 35407 2274 35416 2301
rect 35364 2249 35416 2274
rect 35364 2236 35416 2237
rect 35364 2202 35373 2236
rect 35373 2202 35407 2236
rect 35407 2202 35416 2236
rect 35364 2185 35416 2202
rect 35364 2164 35416 2173
rect 35364 2130 35373 2164
rect 35373 2130 35407 2164
rect 35407 2130 35416 2164
rect 35364 2121 35416 2130
rect 35364 2092 35416 2109
rect 35364 2058 35373 2092
rect 35373 2058 35407 2092
rect 35407 2058 35416 2092
rect 35364 2057 35416 2058
rect 35364 2020 35416 2045
rect 35364 1993 35373 2020
rect 35373 1993 35407 2020
rect 35407 1993 35416 2020
rect 35364 1948 35416 1981
rect 35364 1929 35373 1948
rect 35373 1929 35407 1948
rect 35407 1929 35416 1948
rect 35364 1914 35373 1917
rect 35373 1914 35407 1917
rect 35407 1914 35416 1917
rect 35364 1876 35416 1914
rect 35364 1865 35373 1876
rect 35373 1865 35407 1876
rect 35407 1865 35416 1876
rect 35364 1842 35373 1853
rect 35373 1842 35407 1853
rect 35407 1842 35416 1853
rect 35364 1804 35416 1842
rect 35364 1801 35373 1804
rect 35373 1801 35407 1804
rect 35407 1801 35416 1804
rect 35364 1770 35373 1789
rect 35373 1770 35407 1789
rect 35407 1770 35416 1789
rect 35364 1737 35416 1770
rect 35364 1698 35373 1725
rect 35373 1698 35407 1725
rect 35407 1698 35416 1725
rect 35364 1673 35416 1698
rect 35364 1660 35416 1661
rect 35364 1626 35373 1660
rect 35373 1626 35407 1660
rect 35407 1626 35416 1660
rect 35364 1609 35416 1626
rect 35364 1588 35416 1597
rect 35364 1554 35373 1588
rect 35373 1554 35407 1588
rect 35407 1554 35416 1588
rect 35364 1545 35416 1554
rect 35364 1516 35416 1533
rect 35364 1482 35373 1516
rect 35373 1482 35407 1516
rect 35407 1482 35416 1516
rect 35364 1481 35416 1482
rect 35364 1444 35416 1469
rect 35364 1417 35373 1444
rect 35373 1417 35407 1444
rect 35407 1417 35416 1444
rect 35364 1372 35416 1405
rect 35364 1353 35373 1372
rect 35373 1353 35407 1372
rect 35407 1353 35416 1372
rect 35364 1338 35373 1341
rect 35373 1338 35407 1341
rect 35407 1338 35416 1341
rect 35364 1300 35416 1338
rect 35364 1289 35373 1300
rect 35373 1289 35407 1300
rect 35407 1289 35416 1300
rect 35364 1266 35373 1277
rect 35373 1266 35407 1277
rect 35407 1266 35416 1277
rect 35364 1228 35416 1266
rect 35364 1225 35373 1228
rect 35373 1225 35407 1228
rect 35407 1225 35416 1228
rect 35364 1194 35373 1213
rect 35373 1194 35407 1213
rect 35407 1194 35416 1213
rect 35364 1161 35416 1194
rect 35460 3100 35512 3133
rect 35460 3081 35469 3100
rect 35469 3081 35503 3100
rect 35503 3081 35512 3100
rect 35460 3066 35469 3069
rect 35469 3066 35503 3069
rect 35503 3066 35512 3069
rect 35460 3028 35512 3066
rect 35460 3017 35469 3028
rect 35469 3017 35503 3028
rect 35503 3017 35512 3028
rect 35460 2994 35469 3005
rect 35469 2994 35503 3005
rect 35503 2994 35512 3005
rect 35460 2956 35512 2994
rect 35460 2953 35469 2956
rect 35469 2953 35503 2956
rect 35503 2953 35512 2956
rect 35460 2922 35469 2941
rect 35469 2922 35503 2941
rect 35503 2922 35512 2941
rect 35460 2889 35512 2922
rect 35460 2850 35469 2877
rect 35469 2850 35503 2877
rect 35503 2850 35512 2877
rect 35460 2825 35512 2850
rect 35460 2812 35512 2813
rect 35460 2778 35469 2812
rect 35469 2778 35503 2812
rect 35503 2778 35512 2812
rect 35460 2761 35512 2778
rect 35460 2740 35512 2749
rect 35460 2706 35469 2740
rect 35469 2706 35503 2740
rect 35503 2706 35512 2740
rect 35460 2697 35512 2706
rect 35460 2668 35512 2685
rect 35460 2634 35469 2668
rect 35469 2634 35503 2668
rect 35503 2634 35512 2668
rect 35460 2633 35512 2634
rect 35460 2596 35512 2621
rect 35460 2569 35469 2596
rect 35469 2569 35503 2596
rect 35503 2569 35512 2596
rect 35460 2524 35512 2557
rect 35460 2505 35469 2524
rect 35469 2505 35503 2524
rect 35503 2505 35512 2524
rect 35460 2490 35469 2493
rect 35469 2490 35503 2493
rect 35503 2490 35512 2493
rect 35460 2452 35512 2490
rect 35460 2441 35469 2452
rect 35469 2441 35503 2452
rect 35503 2441 35512 2452
rect 35460 2418 35469 2429
rect 35469 2418 35503 2429
rect 35503 2418 35512 2429
rect 35460 2380 35512 2418
rect 35460 2377 35469 2380
rect 35469 2377 35503 2380
rect 35503 2377 35512 2380
rect 35460 2346 35469 2365
rect 35469 2346 35503 2365
rect 35503 2346 35512 2365
rect 35460 2313 35512 2346
rect 35460 2274 35469 2301
rect 35469 2274 35503 2301
rect 35503 2274 35512 2301
rect 35460 2249 35512 2274
rect 35460 2236 35512 2237
rect 35460 2202 35469 2236
rect 35469 2202 35503 2236
rect 35503 2202 35512 2236
rect 35460 2185 35512 2202
rect 35460 2164 35512 2173
rect 35460 2130 35469 2164
rect 35469 2130 35503 2164
rect 35503 2130 35512 2164
rect 35460 2121 35512 2130
rect 35460 2092 35512 2109
rect 35460 2058 35469 2092
rect 35469 2058 35503 2092
rect 35503 2058 35512 2092
rect 35460 2057 35512 2058
rect 35460 2020 35512 2045
rect 35460 1993 35469 2020
rect 35469 1993 35503 2020
rect 35503 1993 35512 2020
rect 35460 1948 35512 1981
rect 35460 1929 35469 1948
rect 35469 1929 35503 1948
rect 35503 1929 35512 1948
rect 35460 1914 35469 1917
rect 35469 1914 35503 1917
rect 35503 1914 35512 1917
rect 35460 1876 35512 1914
rect 35460 1865 35469 1876
rect 35469 1865 35503 1876
rect 35503 1865 35512 1876
rect 35460 1842 35469 1853
rect 35469 1842 35503 1853
rect 35503 1842 35512 1853
rect 35460 1804 35512 1842
rect 35460 1801 35469 1804
rect 35469 1801 35503 1804
rect 35503 1801 35512 1804
rect 35460 1770 35469 1789
rect 35469 1770 35503 1789
rect 35503 1770 35512 1789
rect 35460 1737 35512 1770
rect 35460 1698 35469 1725
rect 35469 1698 35503 1725
rect 35503 1698 35512 1725
rect 35460 1673 35512 1698
rect 35460 1660 35512 1661
rect 35460 1626 35469 1660
rect 35469 1626 35503 1660
rect 35503 1626 35512 1660
rect 35460 1609 35512 1626
rect 35460 1588 35512 1597
rect 35460 1554 35469 1588
rect 35469 1554 35503 1588
rect 35503 1554 35512 1588
rect 35460 1545 35512 1554
rect 35460 1516 35512 1533
rect 35460 1482 35469 1516
rect 35469 1482 35503 1516
rect 35503 1482 35512 1516
rect 35460 1481 35512 1482
rect 35460 1444 35512 1469
rect 35460 1417 35469 1444
rect 35469 1417 35503 1444
rect 35503 1417 35512 1444
rect 35460 1372 35512 1405
rect 35460 1353 35469 1372
rect 35469 1353 35503 1372
rect 35503 1353 35512 1372
rect 35460 1338 35469 1341
rect 35469 1338 35503 1341
rect 35503 1338 35512 1341
rect 35460 1300 35512 1338
rect 35460 1289 35469 1300
rect 35469 1289 35503 1300
rect 35503 1289 35512 1300
rect 35460 1266 35469 1277
rect 35469 1266 35503 1277
rect 35503 1266 35512 1277
rect 35460 1228 35512 1266
rect 35460 1225 35469 1228
rect 35469 1225 35503 1228
rect 35503 1225 35512 1228
rect 35460 1194 35469 1213
rect 35469 1194 35503 1213
rect 35503 1194 35512 1213
rect 35460 1161 35512 1194
rect 35556 3100 35608 3133
rect 35556 3081 35565 3100
rect 35565 3081 35599 3100
rect 35599 3081 35608 3100
rect 35556 3066 35565 3069
rect 35565 3066 35599 3069
rect 35599 3066 35608 3069
rect 35556 3028 35608 3066
rect 35556 3017 35565 3028
rect 35565 3017 35599 3028
rect 35599 3017 35608 3028
rect 35556 2994 35565 3005
rect 35565 2994 35599 3005
rect 35599 2994 35608 3005
rect 35556 2956 35608 2994
rect 35556 2953 35565 2956
rect 35565 2953 35599 2956
rect 35599 2953 35608 2956
rect 35556 2922 35565 2941
rect 35565 2922 35599 2941
rect 35599 2922 35608 2941
rect 35556 2889 35608 2922
rect 35556 2850 35565 2877
rect 35565 2850 35599 2877
rect 35599 2850 35608 2877
rect 35556 2825 35608 2850
rect 35556 2812 35608 2813
rect 35556 2778 35565 2812
rect 35565 2778 35599 2812
rect 35599 2778 35608 2812
rect 35556 2761 35608 2778
rect 35556 2740 35608 2749
rect 35556 2706 35565 2740
rect 35565 2706 35599 2740
rect 35599 2706 35608 2740
rect 35556 2697 35608 2706
rect 35556 2668 35608 2685
rect 35556 2634 35565 2668
rect 35565 2634 35599 2668
rect 35599 2634 35608 2668
rect 35556 2633 35608 2634
rect 35556 2596 35608 2621
rect 35556 2569 35565 2596
rect 35565 2569 35599 2596
rect 35599 2569 35608 2596
rect 35556 2524 35608 2557
rect 35556 2505 35565 2524
rect 35565 2505 35599 2524
rect 35599 2505 35608 2524
rect 35556 2490 35565 2493
rect 35565 2490 35599 2493
rect 35599 2490 35608 2493
rect 35556 2452 35608 2490
rect 35556 2441 35565 2452
rect 35565 2441 35599 2452
rect 35599 2441 35608 2452
rect 35556 2418 35565 2429
rect 35565 2418 35599 2429
rect 35599 2418 35608 2429
rect 35556 2380 35608 2418
rect 35556 2377 35565 2380
rect 35565 2377 35599 2380
rect 35599 2377 35608 2380
rect 35556 2346 35565 2365
rect 35565 2346 35599 2365
rect 35599 2346 35608 2365
rect 35556 2313 35608 2346
rect 35556 2274 35565 2301
rect 35565 2274 35599 2301
rect 35599 2274 35608 2301
rect 35556 2249 35608 2274
rect 35556 2236 35608 2237
rect 35556 2202 35565 2236
rect 35565 2202 35599 2236
rect 35599 2202 35608 2236
rect 35556 2185 35608 2202
rect 35556 2164 35608 2173
rect 35556 2130 35565 2164
rect 35565 2130 35599 2164
rect 35599 2130 35608 2164
rect 35556 2121 35608 2130
rect 35556 2092 35608 2109
rect 35556 2058 35565 2092
rect 35565 2058 35599 2092
rect 35599 2058 35608 2092
rect 35556 2057 35608 2058
rect 35556 2020 35608 2045
rect 35556 1993 35565 2020
rect 35565 1993 35599 2020
rect 35599 1993 35608 2020
rect 35556 1948 35608 1981
rect 35556 1929 35565 1948
rect 35565 1929 35599 1948
rect 35599 1929 35608 1948
rect 35556 1914 35565 1917
rect 35565 1914 35599 1917
rect 35599 1914 35608 1917
rect 35556 1876 35608 1914
rect 35556 1865 35565 1876
rect 35565 1865 35599 1876
rect 35599 1865 35608 1876
rect 35556 1842 35565 1853
rect 35565 1842 35599 1853
rect 35599 1842 35608 1853
rect 35556 1804 35608 1842
rect 35556 1801 35565 1804
rect 35565 1801 35599 1804
rect 35599 1801 35608 1804
rect 35556 1770 35565 1789
rect 35565 1770 35599 1789
rect 35599 1770 35608 1789
rect 35556 1737 35608 1770
rect 35556 1698 35565 1725
rect 35565 1698 35599 1725
rect 35599 1698 35608 1725
rect 35556 1673 35608 1698
rect 35556 1660 35608 1661
rect 35556 1626 35565 1660
rect 35565 1626 35599 1660
rect 35599 1626 35608 1660
rect 35556 1609 35608 1626
rect 35556 1588 35608 1597
rect 35556 1554 35565 1588
rect 35565 1554 35599 1588
rect 35599 1554 35608 1588
rect 35556 1545 35608 1554
rect 35556 1516 35608 1533
rect 35556 1482 35565 1516
rect 35565 1482 35599 1516
rect 35599 1482 35608 1516
rect 35556 1481 35608 1482
rect 35556 1444 35608 1469
rect 35556 1417 35565 1444
rect 35565 1417 35599 1444
rect 35599 1417 35608 1444
rect 35556 1372 35608 1405
rect 35556 1353 35565 1372
rect 35565 1353 35599 1372
rect 35599 1353 35608 1372
rect 35556 1338 35565 1341
rect 35565 1338 35599 1341
rect 35599 1338 35608 1341
rect 35556 1300 35608 1338
rect 35556 1289 35565 1300
rect 35565 1289 35599 1300
rect 35599 1289 35608 1300
rect 35556 1266 35565 1277
rect 35565 1266 35599 1277
rect 35599 1266 35608 1277
rect 35556 1228 35608 1266
rect 35556 1225 35565 1228
rect 35565 1225 35599 1228
rect 35599 1225 35608 1228
rect 35556 1194 35565 1213
rect 35565 1194 35599 1213
rect 35599 1194 35608 1213
rect 35556 1161 35608 1194
rect 35652 3100 35704 3133
rect 35652 3081 35661 3100
rect 35661 3081 35695 3100
rect 35695 3081 35704 3100
rect 35652 3066 35661 3069
rect 35661 3066 35695 3069
rect 35695 3066 35704 3069
rect 35652 3028 35704 3066
rect 35652 3017 35661 3028
rect 35661 3017 35695 3028
rect 35695 3017 35704 3028
rect 35652 2994 35661 3005
rect 35661 2994 35695 3005
rect 35695 2994 35704 3005
rect 35652 2956 35704 2994
rect 35652 2953 35661 2956
rect 35661 2953 35695 2956
rect 35695 2953 35704 2956
rect 35652 2922 35661 2941
rect 35661 2922 35695 2941
rect 35695 2922 35704 2941
rect 35652 2889 35704 2922
rect 35652 2850 35661 2877
rect 35661 2850 35695 2877
rect 35695 2850 35704 2877
rect 35652 2825 35704 2850
rect 35652 2812 35704 2813
rect 35652 2778 35661 2812
rect 35661 2778 35695 2812
rect 35695 2778 35704 2812
rect 35652 2761 35704 2778
rect 35652 2740 35704 2749
rect 35652 2706 35661 2740
rect 35661 2706 35695 2740
rect 35695 2706 35704 2740
rect 35652 2697 35704 2706
rect 35652 2668 35704 2685
rect 35652 2634 35661 2668
rect 35661 2634 35695 2668
rect 35695 2634 35704 2668
rect 35652 2633 35704 2634
rect 35652 2596 35704 2621
rect 35652 2569 35661 2596
rect 35661 2569 35695 2596
rect 35695 2569 35704 2596
rect 35652 2524 35704 2557
rect 35652 2505 35661 2524
rect 35661 2505 35695 2524
rect 35695 2505 35704 2524
rect 35652 2490 35661 2493
rect 35661 2490 35695 2493
rect 35695 2490 35704 2493
rect 35652 2452 35704 2490
rect 35652 2441 35661 2452
rect 35661 2441 35695 2452
rect 35695 2441 35704 2452
rect 35652 2418 35661 2429
rect 35661 2418 35695 2429
rect 35695 2418 35704 2429
rect 35652 2380 35704 2418
rect 35652 2377 35661 2380
rect 35661 2377 35695 2380
rect 35695 2377 35704 2380
rect 35652 2346 35661 2365
rect 35661 2346 35695 2365
rect 35695 2346 35704 2365
rect 35652 2313 35704 2346
rect 35652 2274 35661 2301
rect 35661 2274 35695 2301
rect 35695 2274 35704 2301
rect 35652 2249 35704 2274
rect 35652 2236 35704 2237
rect 35652 2202 35661 2236
rect 35661 2202 35695 2236
rect 35695 2202 35704 2236
rect 35652 2185 35704 2202
rect 35652 2164 35704 2173
rect 35652 2130 35661 2164
rect 35661 2130 35695 2164
rect 35695 2130 35704 2164
rect 35652 2121 35704 2130
rect 35652 2092 35704 2109
rect 35652 2058 35661 2092
rect 35661 2058 35695 2092
rect 35695 2058 35704 2092
rect 35652 2057 35704 2058
rect 35652 2020 35704 2045
rect 35652 1993 35661 2020
rect 35661 1993 35695 2020
rect 35695 1993 35704 2020
rect 35652 1948 35704 1981
rect 35652 1929 35661 1948
rect 35661 1929 35695 1948
rect 35695 1929 35704 1948
rect 35652 1914 35661 1917
rect 35661 1914 35695 1917
rect 35695 1914 35704 1917
rect 35652 1876 35704 1914
rect 35652 1865 35661 1876
rect 35661 1865 35695 1876
rect 35695 1865 35704 1876
rect 35652 1842 35661 1853
rect 35661 1842 35695 1853
rect 35695 1842 35704 1853
rect 35652 1804 35704 1842
rect 35652 1801 35661 1804
rect 35661 1801 35695 1804
rect 35695 1801 35704 1804
rect 35652 1770 35661 1789
rect 35661 1770 35695 1789
rect 35695 1770 35704 1789
rect 35652 1737 35704 1770
rect 35652 1698 35661 1725
rect 35661 1698 35695 1725
rect 35695 1698 35704 1725
rect 35652 1673 35704 1698
rect 35652 1660 35704 1661
rect 35652 1626 35661 1660
rect 35661 1626 35695 1660
rect 35695 1626 35704 1660
rect 35652 1609 35704 1626
rect 35652 1588 35704 1597
rect 35652 1554 35661 1588
rect 35661 1554 35695 1588
rect 35695 1554 35704 1588
rect 35652 1545 35704 1554
rect 35652 1516 35704 1533
rect 35652 1482 35661 1516
rect 35661 1482 35695 1516
rect 35695 1482 35704 1516
rect 35652 1481 35704 1482
rect 35652 1444 35704 1469
rect 35652 1417 35661 1444
rect 35661 1417 35695 1444
rect 35695 1417 35704 1444
rect 35652 1372 35704 1405
rect 35652 1353 35661 1372
rect 35661 1353 35695 1372
rect 35695 1353 35704 1372
rect 35652 1338 35661 1341
rect 35661 1338 35695 1341
rect 35695 1338 35704 1341
rect 35652 1300 35704 1338
rect 35652 1289 35661 1300
rect 35661 1289 35695 1300
rect 35695 1289 35704 1300
rect 35652 1266 35661 1277
rect 35661 1266 35695 1277
rect 35695 1266 35704 1277
rect 35652 1228 35704 1266
rect 35652 1225 35661 1228
rect 35661 1225 35695 1228
rect 35695 1225 35704 1228
rect 35652 1194 35661 1213
rect 35661 1194 35695 1213
rect 35695 1194 35704 1213
rect 35652 1161 35704 1194
rect 35748 3100 35800 3133
rect 35748 3081 35757 3100
rect 35757 3081 35791 3100
rect 35791 3081 35800 3100
rect 35748 3066 35757 3069
rect 35757 3066 35791 3069
rect 35791 3066 35800 3069
rect 35748 3028 35800 3066
rect 35748 3017 35757 3028
rect 35757 3017 35791 3028
rect 35791 3017 35800 3028
rect 35748 2994 35757 3005
rect 35757 2994 35791 3005
rect 35791 2994 35800 3005
rect 35748 2956 35800 2994
rect 35748 2953 35757 2956
rect 35757 2953 35791 2956
rect 35791 2953 35800 2956
rect 35748 2922 35757 2941
rect 35757 2922 35791 2941
rect 35791 2922 35800 2941
rect 35748 2889 35800 2922
rect 35748 2850 35757 2877
rect 35757 2850 35791 2877
rect 35791 2850 35800 2877
rect 35748 2825 35800 2850
rect 35748 2812 35800 2813
rect 35748 2778 35757 2812
rect 35757 2778 35791 2812
rect 35791 2778 35800 2812
rect 35748 2761 35800 2778
rect 35748 2740 35800 2749
rect 35748 2706 35757 2740
rect 35757 2706 35791 2740
rect 35791 2706 35800 2740
rect 35748 2697 35800 2706
rect 35748 2668 35800 2685
rect 35748 2634 35757 2668
rect 35757 2634 35791 2668
rect 35791 2634 35800 2668
rect 35748 2633 35800 2634
rect 35748 2596 35800 2621
rect 35748 2569 35757 2596
rect 35757 2569 35791 2596
rect 35791 2569 35800 2596
rect 35748 2524 35800 2557
rect 35748 2505 35757 2524
rect 35757 2505 35791 2524
rect 35791 2505 35800 2524
rect 35748 2490 35757 2493
rect 35757 2490 35791 2493
rect 35791 2490 35800 2493
rect 35748 2452 35800 2490
rect 35748 2441 35757 2452
rect 35757 2441 35791 2452
rect 35791 2441 35800 2452
rect 35748 2418 35757 2429
rect 35757 2418 35791 2429
rect 35791 2418 35800 2429
rect 35748 2380 35800 2418
rect 35748 2377 35757 2380
rect 35757 2377 35791 2380
rect 35791 2377 35800 2380
rect 35748 2346 35757 2365
rect 35757 2346 35791 2365
rect 35791 2346 35800 2365
rect 35748 2313 35800 2346
rect 35748 2274 35757 2301
rect 35757 2274 35791 2301
rect 35791 2274 35800 2301
rect 35748 2249 35800 2274
rect 35748 2236 35800 2237
rect 35748 2202 35757 2236
rect 35757 2202 35791 2236
rect 35791 2202 35800 2236
rect 35748 2185 35800 2202
rect 35748 2164 35800 2173
rect 35748 2130 35757 2164
rect 35757 2130 35791 2164
rect 35791 2130 35800 2164
rect 35748 2121 35800 2130
rect 35748 2092 35800 2109
rect 35748 2058 35757 2092
rect 35757 2058 35791 2092
rect 35791 2058 35800 2092
rect 35748 2057 35800 2058
rect 35748 2020 35800 2045
rect 35748 1993 35757 2020
rect 35757 1993 35791 2020
rect 35791 1993 35800 2020
rect 35748 1948 35800 1981
rect 35748 1929 35757 1948
rect 35757 1929 35791 1948
rect 35791 1929 35800 1948
rect 35748 1914 35757 1917
rect 35757 1914 35791 1917
rect 35791 1914 35800 1917
rect 35748 1876 35800 1914
rect 35748 1865 35757 1876
rect 35757 1865 35791 1876
rect 35791 1865 35800 1876
rect 35748 1842 35757 1853
rect 35757 1842 35791 1853
rect 35791 1842 35800 1853
rect 35748 1804 35800 1842
rect 35748 1801 35757 1804
rect 35757 1801 35791 1804
rect 35791 1801 35800 1804
rect 35748 1770 35757 1789
rect 35757 1770 35791 1789
rect 35791 1770 35800 1789
rect 35748 1737 35800 1770
rect 35748 1698 35757 1725
rect 35757 1698 35791 1725
rect 35791 1698 35800 1725
rect 35748 1673 35800 1698
rect 35748 1660 35800 1661
rect 35748 1626 35757 1660
rect 35757 1626 35791 1660
rect 35791 1626 35800 1660
rect 35748 1609 35800 1626
rect 35748 1588 35800 1597
rect 35748 1554 35757 1588
rect 35757 1554 35791 1588
rect 35791 1554 35800 1588
rect 35748 1545 35800 1554
rect 35748 1516 35800 1533
rect 35748 1482 35757 1516
rect 35757 1482 35791 1516
rect 35791 1482 35800 1516
rect 35748 1481 35800 1482
rect 35748 1444 35800 1469
rect 35748 1417 35757 1444
rect 35757 1417 35791 1444
rect 35791 1417 35800 1444
rect 35748 1372 35800 1405
rect 35748 1353 35757 1372
rect 35757 1353 35791 1372
rect 35791 1353 35800 1372
rect 35748 1338 35757 1341
rect 35757 1338 35791 1341
rect 35791 1338 35800 1341
rect 35748 1300 35800 1338
rect 35748 1289 35757 1300
rect 35757 1289 35791 1300
rect 35791 1289 35800 1300
rect 35748 1266 35757 1277
rect 35757 1266 35791 1277
rect 35791 1266 35800 1277
rect 35748 1228 35800 1266
rect 35748 1225 35757 1228
rect 35757 1225 35791 1228
rect 35791 1225 35800 1228
rect 35748 1194 35757 1213
rect 35757 1194 35791 1213
rect 35791 1194 35800 1213
rect 35748 1161 35800 1194
rect 35844 3100 35896 3133
rect 35844 3081 35853 3100
rect 35853 3081 35887 3100
rect 35887 3081 35896 3100
rect 35844 3066 35853 3069
rect 35853 3066 35887 3069
rect 35887 3066 35896 3069
rect 35844 3028 35896 3066
rect 35844 3017 35853 3028
rect 35853 3017 35887 3028
rect 35887 3017 35896 3028
rect 35844 2994 35853 3005
rect 35853 2994 35887 3005
rect 35887 2994 35896 3005
rect 35844 2956 35896 2994
rect 35844 2953 35853 2956
rect 35853 2953 35887 2956
rect 35887 2953 35896 2956
rect 35844 2922 35853 2941
rect 35853 2922 35887 2941
rect 35887 2922 35896 2941
rect 35844 2889 35896 2922
rect 35844 2850 35853 2877
rect 35853 2850 35887 2877
rect 35887 2850 35896 2877
rect 35844 2825 35896 2850
rect 35844 2812 35896 2813
rect 35844 2778 35853 2812
rect 35853 2778 35887 2812
rect 35887 2778 35896 2812
rect 35844 2761 35896 2778
rect 35844 2740 35896 2749
rect 35844 2706 35853 2740
rect 35853 2706 35887 2740
rect 35887 2706 35896 2740
rect 35844 2697 35896 2706
rect 35844 2668 35896 2685
rect 35844 2634 35853 2668
rect 35853 2634 35887 2668
rect 35887 2634 35896 2668
rect 35844 2633 35896 2634
rect 35844 2596 35896 2621
rect 35844 2569 35853 2596
rect 35853 2569 35887 2596
rect 35887 2569 35896 2596
rect 35844 2524 35896 2557
rect 35844 2505 35853 2524
rect 35853 2505 35887 2524
rect 35887 2505 35896 2524
rect 35844 2490 35853 2493
rect 35853 2490 35887 2493
rect 35887 2490 35896 2493
rect 35844 2452 35896 2490
rect 35844 2441 35853 2452
rect 35853 2441 35887 2452
rect 35887 2441 35896 2452
rect 35844 2418 35853 2429
rect 35853 2418 35887 2429
rect 35887 2418 35896 2429
rect 35844 2380 35896 2418
rect 35844 2377 35853 2380
rect 35853 2377 35887 2380
rect 35887 2377 35896 2380
rect 35844 2346 35853 2365
rect 35853 2346 35887 2365
rect 35887 2346 35896 2365
rect 35844 2313 35896 2346
rect 35844 2274 35853 2301
rect 35853 2274 35887 2301
rect 35887 2274 35896 2301
rect 35844 2249 35896 2274
rect 35844 2236 35896 2237
rect 35844 2202 35853 2236
rect 35853 2202 35887 2236
rect 35887 2202 35896 2236
rect 35844 2185 35896 2202
rect 35844 2164 35896 2173
rect 35844 2130 35853 2164
rect 35853 2130 35887 2164
rect 35887 2130 35896 2164
rect 35844 2121 35896 2130
rect 35844 2092 35896 2109
rect 35844 2058 35853 2092
rect 35853 2058 35887 2092
rect 35887 2058 35896 2092
rect 35844 2057 35896 2058
rect 35844 2020 35896 2045
rect 35844 1993 35853 2020
rect 35853 1993 35887 2020
rect 35887 1993 35896 2020
rect 35844 1948 35896 1981
rect 35844 1929 35853 1948
rect 35853 1929 35887 1948
rect 35887 1929 35896 1948
rect 35844 1914 35853 1917
rect 35853 1914 35887 1917
rect 35887 1914 35896 1917
rect 35844 1876 35896 1914
rect 35844 1865 35853 1876
rect 35853 1865 35887 1876
rect 35887 1865 35896 1876
rect 35844 1842 35853 1853
rect 35853 1842 35887 1853
rect 35887 1842 35896 1853
rect 35844 1804 35896 1842
rect 35844 1801 35853 1804
rect 35853 1801 35887 1804
rect 35887 1801 35896 1804
rect 35844 1770 35853 1789
rect 35853 1770 35887 1789
rect 35887 1770 35896 1789
rect 35844 1737 35896 1770
rect 35844 1698 35853 1725
rect 35853 1698 35887 1725
rect 35887 1698 35896 1725
rect 35844 1673 35896 1698
rect 35844 1660 35896 1661
rect 35844 1626 35853 1660
rect 35853 1626 35887 1660
rect 35887 1626 35896 1660
rect 35844 1609 35896 1626
rect 35844 1588 35896 1597
rect 35844 1554 35853 1588
rect 35853 1554 35887 1588
rect 35887 1554 35896 1588
rect 35844 1545 35896 1554
rect 35844 1516 35896 1533
rect 35844 1482 35853 1516
rect 35853 1482 35887 1516
rect 35887 1482 35896 1516
rect 35844 1481 35896 1482
rect 35844 1444 35896 1469
rect 35844 1417 35853 1444
rect 35853 1417 35887 1444
rect 35887 1417 35896 1444
rect 35844 1372 35896 1405
rect 35844 1353 35853 1372
rect 35853 1353 35887 1372
rect 35887 1353 35896 1372
rect 35844 1338 35853 1341
rect 35853 1338 35887 1341
rect 35887 1338 35896 1341
rect 35844 1300 35896 1338
rect 35844 1289 35853 1300
rect 35853 1289 35887 1300
rect 35887 1289 35896 1300
rect 35844 1266 35853 1277
rect 35853 1266 35887 1277
rect 35887 1266 35896 1277
rect 35844 1228 35896 1266
rect 35844 1225 35853 1228
rect 35853 1225 35887 1228
rect 35887 1225 35896 1228
rect 35844 1194 35853 1213
rect 35853 1194 35887 1213
rect 35887 1194 35896 1213
rect 35844 1161 35896 1194
rect 35940 3100 35992 3133
rect 35940 3081 35949 3100
rect 35949 3081 35983 3100
rect 35983 3081 35992 3100
rect 35940 3066 35949 3069
rect 35949 3066 35983 3069
rect 35983 3066 35992 3069
rect 35940 3028 35992 3066
rect 35940 3017 35949 3028
rect 35949 3017 35983 3028
rect 35983 3017 35992 3028
rect 35940 2994 35949 3005
rect 35949 2994 35983 3005
rect 35983 2994 35992 3005
rect 35940 2956 35992 2994
rect 35940 2953 35949 2956
rect 35949 2953 35983 2956
rect 35983 2953 35992 2956
rect 35940 2922 35949 2941
rect 35949 2922 35983 2941
rect 35983 2922 35992 2941
rect 35940 2889 35992 2922
rect 35940 2850 35949 2877
rect 35949 2850 35983 2877
rect 35983 2850 35992 2877
rect 35940 2825 35992 2850
rect 35940 2812 35992 2813
rect 35940 2778 35949 2812
rect 35949 2778 35983 2812
rect 35983 2778 35992 2812
rect 35940 2761 35992 2778
rect 35940 2740 35992 2749
rect 35940 2706 35949 2740
rect 35949 2706 35983 2740
rect 35983 2706 35992 2740
rect 35940 2697 35992 2706
rect 35940 2668 35992 2685
rect 35940 2634 35949 2668
rect 35949 2634 35983 2668
rect 35983 2634 35992 2668
rect 35940 2633 35992 2634
rect 35940 2596 35992 2621
rect 35940 2569 35949 2596
rect 35949 2569 35983 2596
rect 35983 2569 35992 2596
rect 35940 2524 35992 2557
rect 35940 2505 35949 2524
rect 35949 2505 35983 2524
rect 35983 2505 35992 2524
rect 35940 2490 35949 2493
rect 35949 2490 35983 2493
rect 35983 2490 35992 2493
rect 35940 2452 35992 2490
rect 35940 2441 35949 2452
rect 35949 2441 35983 2452
rect 35983 2441 35992 2452
rect 35940 2418 35949 2429
rect 35949 2418 35983 2429
rect 35983 2418 35992 2429
rect 35940 2380 35992 2418
rect 35940 2377 35949 2380
rect 35949 2377 35983 2380
rect 35983 2377 35992 2380
rect 35940 2346 35949 2365
rect 35949 2346 35983 2365
rect 35983 2346 35992 2365
rect 35940 2313 35992 2346
rect 35940 2274 35949 2301
rect 35949 2274 35983 2301
rect 35983 2274 35992 2301
rect 35940 2249 35992 2274
rect 35940 2236 35992 2237
rect 35940 2202 35949 2236
rect 35949 2202 35983 2236
rect 35983 2202 35992 2236
rect 35940 2185 35992 2202
rect 35940 2164 35992 2173
rect 35940 2130 35949 2164
rect 35949 2130 35983 2164
rect 35983 2130 35992 2164
rect 35940 2121 35992 2130
rect 35940 2092 35992 2109
rect 35940 2058 35949 2092
rect 35949 2058 35983 2092
rect 35983 2058 35992 2092
rect 35940 2057 35992 2058
rect 35940 2020 35992 2045
rect 35940 1993 35949 2020
rect 35949 1993 35983 2020
rect 35983 1993 35992 2020
rect 35940 1948 35992 1981
rect 35940 1929 35949 1948
rect 35949 1929 35983 1948
rect 35983 1929 35992 1948
rect 35940 1914 35949 1917
rect 35949 1914 35983 1917
rect 35983 1914 35992 1917
rect 35940 1876 35992 1914
rect 35940 1865 35949 1876
rect 35949 1865 35983 1876
rect 35983 1865 35992 1876
rect 35940 1842 35949 1853
rect 35949 1842 35983 1853
rect 35983 1842 35992 1853
rect 35940 1804 35992 1842
rect 35940 1801 35949 1804
rect 35949 1801 35983 1804
rect 35983 1801 35992 1804
rect 35940 1770 35949 1789
rect 35949 1770 35983 1789
rect 35983 1770 35992 1789
rect 35940 1737 35992 1770
rect 35940 1698 35949 1725
rect 35949 1698 35983 1725
rect 35983 1698 35992 1725
rect 35940 1673 35992 1698
rect 35940 1660 35992 1661
rect 35940 1626 35949 1660
rect 35949 1626 35983 1660
rect 35983 1626 35992 1660
rect 35940 1609 35992 1626
rect 35940 1588 35992 1597
rect 35940 1554 35949 1588
rect 35949 1554 35983 1588
rect 35983 1554 35992 1588
rect 35940 1545 35992 1554
rect 35940 1516 35992 1533
rect 35940 1482 35949 1516
rect 35949 1482 35983 1516
rect 35983 1482 35992 1516
rect 35940 1481 35992 1482
rect 35940 1444 35992 1469
rect 35940 1417 35949 1444
rect 35949 1417 35983 1444
rect 35983 1417 35992 1444
rect 35940 1372 35992 1405
rect 35940 1353 35949 1372
rect 35949 1353 35983 1372
rect 35983 1353 35992 1372
rect 35940 1338 35949 1341
rect 35949 1338 35983 1341
rect 35983 1338 35992 1341
rect 35940 1300 35992 1338
rect 35940 1289 35949 1300
rect 35949 1289 35983 1300
rect 35983 1289 35992 1300
rect 35940 1266 35949 1277
rect 35949 1266 35983 1277
rect 35983 1266 35992 1277
rect 35940 1228 35992 1266
rect 35940 1225 35949 1228
rect 35949 1225 35983 1228
rect 35983 1225 35992 1228
rect 35940 1194 35949 1213
rect 35949 1194 35983 1213
rect 35983 1194 35992 1213
rect 35940 1161 35992 1194
rect 36036 3100 36088 3133
rect 36036 3081 36045 3100
rect 36045 3081 36079 3100
rect 36079 3081 36088 3100
rect 36036 3066 36045 3069
rect 36045 3066 36079 3069
rect 36079 3066 36088 3069
rect 36036 3028 36088 3066
rect 36036 3017 36045 3028
rect 36045 3017 36079 3028
rect 36079 3017 36088 3028
rect 36036 2994 36045 3005
rect 36045 2994 36079 3005
rect 36079 2994 36088 3005
rect 36036 2956 36088 2994
rect 36036 2953 36045 2956
rect 36045 2953 36079 2956
rect 36079 2953 36088 2956
rect 36036 2922 36045 2941
rect 36045 2922 36079 2941
rect 36079 2922 36088 2941
rect 36036 2889 36088 2922
rect 36036 2850 36045 2877
rect 36045 2850 36079 2877
rect 36079 2850 36088 2877
rect 36036 2825 36088 2850
rect 36036 2812 36088 2813
rect 36036 2778 36045 2812
rect 36045 2778 36079 2812
rect 36079 2778 36088 2812
rect 36036 2761 36088 2778
rect 36036 2740 36088 2749
rect 36036 2706 36045 2740
rect 36045 2706 36079 2740
rect 36079 2706 36088 2740
rect 36036 2697 36088 2706
rect 36036 2668 36088 2685
rect 36036 2634 36045 2668
rect 36045 2634 36079 2668
rect 36079 2634 36088 2668
rect 36036 2633 36088 2634
rect 36036 2596 36088 2621
rect 36036 2569 36045 2596
rect 36045 2569 36079 2596
rect 36079 2569 36088 2596
rect 36036 2524 36088 2557
rect 36036 2505 36045 2524
rect 36045 2505 36079 2524
rect 36079 2505 36088 2524
rect 36036 2490 36045 2493
rect 36045 2490 36079 2493
rect 36079 2490 36088 2493
rect 36036 2452 36088 2490
rect 36036 2441 36045 2452
rect 36045 2441 36079 2452
rect 36079 2441 36088 2452
rect 36036 2418 36045 2429
rect 36045 2418 36079 2429
rect 36079 2418 36088 2429
rect 36036 2380 36088 2418
rect 36036 2377 36045 2380
rect 36045 2377 36079 2380
rect 36079 2377 36088 2380
rect 36036 2346 36045 2365
rect 36045 2346 36079 2365
rect 36079 2346 36088 2365
rect 36036 2313 36088 2346
rect 36036 2274 36045 2301
rect 36045 2274 36079 2301
rect 36079 2274 36088 2301
rect 36036 2249 36088 2274
rect 36036 2236 36088 2237
rect 36036 2202 36045 2236
rect 36045 2202 36079 2236
rect 36079 2202 36088 2236
rect 36036 2185 36088 2202
rect 36036 2164 36088 2173
rect 36036 2130 36045 2164
rect 36045 2130 36079 2164
rect 36079 2130 36088 2164
rect 36036 2121 36088 2130
rect 36036 2092 36088 2109
rect 36036 2058 36045 2092
rect 36045 2058 36079 2092
rect 36079 2058 36088 2092
rect 36036 2057 36088 2058
rect 36036 2020 36088 2045
rect 36036 1993 36045 2020
rect 36045 1993 36079 2020
rect 36079 1993 36088 2020
rect 36036 1948 36088 1981
rect 36036 1929 36045 1948
rect 36045 1929 36079 1948
rect 36079 1929 36088 1948
rect 36036 1914 36045 1917
rect 36045 1914 36079 1917
rect 36079 1914 36088 1917
rect 36036 1876 36088 1914
rect 36036 1865 36045 1876
rect 36045 1865 36079 1876
rect 36079 1865 36088 1876
rect 36036 1842 36045 1853
rect 36045 1842 36079 1853
rect 36079 1842 36088 1853
rect 36036 1804 36088 1842
rect 36036 1801 36045 1804
rect 36045 1801 36079 1804
rect 36079 1801 36088 1804
rect 36036 1770 36045 1789
rect 36045 1770 36079 1789
rect 36079 1770 36088 1789
rect 36036 1737 36088 1770
rect 36036 1698 36045 1725
rect 36045 1698 36079 1725
rect 36079 1698 36088 1725
rect 36036 1673 36088 1698
rect 36036 1660 36088 1661
rect 36036 1626 36045 1660
rect 36045 1626 36079 1660
rect 36079 1626 36088 1660
rect 36036 1609 36088 1626
rect 36036 1588 36088 1597
rect 36036 1554 36045 1588
rect 36045 1554 36079 1588
rect 36079 1554 36088 1588
rect 36036 1545 36088 1554
rect 36036 1516 36088 1533
rect 36036 1482 36045 1516
rect 36045 1482 36079 1516
rect 36079 1482 36088 1516
rect 36036 1481 36088 1482
rect 36036 1444 36088 1469
rect 36036 1417 36045 1444
rect 36045 1417 36079 1444
rect 36079 1417 36088 1444
rect 36036 1372 36088 1405
rect 36036 1353 36045 1372
rect 36045 1353 36079 1372
rect 36079 1353 36088 1372
rect 36036 1338 36045 1341
rect 36045 1338 36079 1341
rect 36079 1338 36088 1341
rect 36036 1300 36088 1338
rect 36036 1289 36045 1300
rect 36045 1289 36079 1300
rect 36079 1289 36088 1300
rect 36036 1266 36045 1277
rect 36045 1266 36079 1277
rect 36079 1266 36088 1277
rect 36036 1228 36088 1266
rect 36036 1225 36045 1228
rect 36045 1225 36079 1228
rect 36079 1225 36088 1228
rect 36036 1194 36045 1213
rect 36045 1194 36079 1213
rect 36079 1194 36088 1213
rect 36036 1161 36088 1194
rect 36132 3100 36184 3133
rect 36132 3081 36141 3100
rect 36141 3081 36175 3100
rect 36175 3081 36184 3100
rect 36132 3066 36141 3069
rect 36141 3066 36175 3069
rect 36175 3066 36184 3069
rect 36132 3028 36184 3066
rect 36132 3017 36141 3028
rect 36141 3017 36175 3028
rect 36175 3017 36184 3028
rect 36132 2994 36141 3005
rect 36141 2994 36175 3005
rect 36175 2994 36184 3005
rect 36132 2956 36184 2994
rect 36132 2953 36141 2956
rect 36141 2953 36175 2956
rect 36175 2953 36184 2956
rect 36132 2922 36141 2941
rect 36141 2922 36175 2941
rect 36175 2922 36184 2941
rect 36132 2889 36184 2922
rect 36132 2850 36141 2877
rect 36141 2850 36175 2877
rect 36175 2850 36184 2877
rect 36132 2825 36184 2850
rect 36132 2812 36184 2813
rect 36132 2778 36141 2812
rect 36141 2778 36175 2812
rect 36175 2778 36184 2812
rect 36132 2761 36184 2778
rect 36132 2740 36184 2749
rect 36132 2706 36141 2740
rect 36141 2706 36175 2740
rect 36175 2706 36184 2740
rect 36132 2697 36184 2706
rect 36132 2668 36184 2685
rect 36132 2634 36141 2668
rect 36141 2634 36175 2668
rect 36175 2634 36184 2668
rect 36132 2633 36184 2634
rect 36132 2596 36184 2621
rect 36132 2569 36141 2596
rect 36141 2569 36175 2596
rect 36175 2569 36184 2596
rect 36132 2524 36184 2557
rect 36132 2505 36141 2524
rect 36141 2505 36175 2524
rect 36175 2505 36184 2524
rect 36132 2490 36141 2493
rect 36141 2490 36175 2493
rect 36175 2490 36184 2493
rect 36132 2452 36184 2490
rect 36132 2441 36141 2452
rect 36141 2441 36175 2452
rect 36175 2441 36184 2452
rect 36132 2418 36141 2429
rect 36141 2418 36175 2429
rect 36175 2418 36184 2429
rect 36132 2380 36184 2418
rect 36132 2377 36141 2380
rect 36141 2377 36175 2380
rect 36175 2377 36184 2380
rect 36132 2346 36141 2365
rect 36141 2346 36175 2365
rect 36175 2346 36184 2365
rect 36132 2313 36184 2346
rect 36132 2274 36141 2301
rect 36141 2274 36175 2301
rect 36175 2274 36184 2301
rect 36132 2249 36184 2274
rect 36132 2236 36184 2237
rect 36132 2202 36141 2236
rect 36141 2202 36175 2236
rect 36175 2202 36184 2236
rect 36132 2185 36184 2202
rect 36132 2164 36184 2173
rect 36132 2130 36141 2164
rect 36141 2130 36175 2164
rect 36175 2130 36184 2164
rect 36132 2121 36184 2130
rect 36132 2092 36184 2109
rect 36132 2058 36141 2092
rect 36141 2058 36175 2092
rect 36175 2058 36184 2092
rect 36132 2057 36184 2058
rect 36132 2020 36184 2045
rect 36132 1993 36141 2020
rect 36141 1993 36175 2020
rect 36175 1993 36184 2020
rect 36132 1948 36184 1981
rect 36132 1929 36141 1948
rect 36141 1929 36175 1948
rect 36175 1929 36184 1948
rect 36132 1914 36141 1917
rect 36141 1914 36175 1917
rect 36175 1914 36184 1917
rect 36132 1876 36184 1914
rect 36132 1865 36141 1876
rect 36141 1865 36175 1876
rect 36175 1865 36184 1876
rect 36132 1842 36141 1853
rect 36141 1842 36175 1853
rect 36175 1842 36184 1853
rect 36132 1804 36184 1842
rect 36132 1801 36141 1804
rect 36141 1801 36175 1804
rect 36175 1801 36184 1804
rect 36132 1770 36141 1789
rect 36141 1770 36175 1789
rect 36175 1770 36184 1789
rect 36132 1737 36184 1770
rect 36132 1698 36141 1725
rect 36141 1698 36175 1725
rect 36175 1698 36184 1725
rect 36132 1673 36184 1698
rect 36132 1660 36184 1661
rect 36132 1626 36141 1660
rect 36141 1626 36175 1660
rect 36175 1626 36184 1660
rect 36132 1609 36184 1626
rect 36132 1588 36184 1597
rect 36132 1554 36141 1588
rect 36141 1554 36175 1588
rect 36175 1554 36184 1588
rect 36132 1545 36184 1554
rect 36132 1516 36184 1533
rect 36132 1482 36141 1516
rect 36141 1482 36175 1516
rect 36175 1482 36184 1516
rect 36132 1481 36184 1482
rect 36132 1444 36184 1469
rect 36132 1417 36141 1444
rect 36141 1417 36175 1444
rect 36175 1417 36184 1444
rect 36132 1372 36184 1405
rect 36132 1353 36141 1372
rect 36141 1353 36175 1372
rect 36175 1353 36184 1372
rect 36132 1338 36141 1341
rect 36141 1338 36175 1341
rect 36175 1338 36184 1341
rect 36132 1300 36184 1338
rect 36132 1289 36141 1300
rect 36141 1289 36175 1300
rect 36175 1289 36184 1300
rect 36132 1266 36141 1277
rect 36141 1266 36175 1277
rect 36175 1266 36184 1277
rect 36132 1228 36184 1266
rect 36132 1225 36141 1228
rect 36141 1225 36175 1228
rect 36175 1225 36184 1228
rect 36132 1194 36141 1213
rect 36141 1194 36175 1213
rect 36175 1194 36184 1213
rect 36132 1161 36184 1194
rect 36228 3100 36280 3133
rect 36228 3081 36237 3100
rect 36237 3081 36271 3100
rect 36271 3081 36280 3100
rect 36228 3066 36237 3069
rect 36237 3066 36271 3069
rect 36271 3066 36280 3069
rect 36228 3028 36280 3066
rect 36228 3017 36237 3028
rect 36237 3017 36271 3028
rect 36271 3017 36280 3028
rect 36228 2994 36237 3005
rect 36237 2994 36271 3005
rect 36271 2994 36280 3005
rect 36228 2956 36280 2994
rect 36228 2953 36237 2956
rect 36237 2953 36271 2956
rect 36271 2953 36280 2956
rect 36228 2922 36237 2941
rect 36237 2922 36271 2941
rect 36271 2922 36280 2941
rect 36228 2889 36280 2922
rect 36228 2850 36237 2877
rect 36237 2850 36271 2877
rect 36271 2850 36280 2877
rect 36228 2825 36280 2850
rect 36228 2812 36280 2813
rect 36228 2778 36237 2812
rect 36237 2778 36271 2812
rect 36271 2778 36280 2812
rect 36228 2761 36280 2778
rect 36228 2740 36280 2749
rect 36228 2706 36237 2740
rect 36237 2706 36271 2740
rect 36271 2706 36280 2740
rect 36228 2697 36280 2706
rect 36228 2668 36280 2685
rect 36228 2634 36237 2668
rect 36237 2634 36271 2668
rect 36271 2634 36280 2668
rect 36228 2633 36280 2634
rect 36228 2596 36280 2621
rect 36228 2569 36237 2596
rect 36237 2569 36271 2596
rect 36271 2569 36280 2596
rect 36228 2524 36280 2557
rect 36228 2505 36237 2524
rect 36237 2505 36271 2524
rect 36271 2505 36280 2524
rect 36228 2490 36237 2493
rect 36237 2490 36271 2493
rect 36271 2490 36280 2493
rect 36228 2452 36280 2490
rect 36228 2441 36237 2452
rect 36237 2441 36271 2452
rect 36271 2441 36280 2452
rect 36228 2418 36237 2429
rect 36237 2418 36271 2429
rect 36271 2418 36280 2429
rect 36228 2380 36280 2418
rect 36228 2377 36237 2380
rect 36237 2377 36271 2380
rect 36271 2377 36280 2380
rect 36228 2346 36237 2365
rect 36237 2346 36271 2365
rect 36271 2346 36280 2365
rect 36228 2313 36280 2346
rect 36228 2274 36237 2301
rect 36237 2274 36271 2301
rect 36271 2274 36280 2301
rect 36228 2249 36280 2274
rect 36228 2236 36280 2237
rect 36228 2202 36237 2236
rect 36237 2202 36271 2236
rect 36271 2202 36280 2236
rect 36228 2185 36280 2202
rect 36228 2164 36280 2173
rect 36228 2130 36237 2164
rect 36237 2130 36271 2164
rect 36271 2130 36280 2164
rect 36228 2121 36280 2130
rect 36228 2092 36280 2109
rect 36228 2058 36237 2092
rect 36237 2058 36271 2092
rect 36271 2058 36280 2092
rect 36228 2057 36280 2058
rect 36228 2020 36280 2045
rect 36228 1993 36237 2020
rect 36237 1993 36271 2020
rect 36271 1993 36280 2020
rect 36228 1948 36280 1981
rect 36228 1929 36237 1948
rect 36237 1929 36271 1948
rect 36271 1929 36280 1948
rect 36228 1914 36237 1917
rect 36237 1914 36271 1917
rect 36271 1914 36280 1917
rect 36228 1876 36280 1914
rect 36228 1865 36237 1876
rect 36237 1865 36271 1876
rect 36271 1865 36280 1876
rect 36228 1842 36237 1853
rect 36237 1842 36271 1853
rect 36271 1842 36280 1853
rect 36228 1804 36280 1842
rect 36228 1801 36237 1804
rect 36237 1801 36271 1804
rect 36271 1801 36280 1804
rect 36228 1770 36237 1789
rect 36237 1770 36271 1789
rect 36271 1770 36280 1789
rect 36228 1737 36280 1770
rect 36228 1698 36237 1725
rect 36237 1698 36271 1725
rect 36271 1698 36280 1725
rect 36228 1673 36280 1698
rect 36228 1660 36280 1661
rect 36228 1626 36237 1660
rect 36237 1626 36271 1660
rect 36271 1626 36280 1660
rect 36228 1609 36280 1626
rect 36228 1588 36280 1597
rect 36228 1554 36237 1588
rect 36237 1554 36271 1588
rect 36271 1554 36280 1588
rect 36228 1545 36280 1554
rect 36228 1516 36280 1533
rect 36228 1482 36237 1516
rect 36237 1482 36271 1516
rect 36271 1482 36280 1516
rect 36228 1481 36280 1482
rect 36228 1444 36280 1469
rect 36228 1417 36237 1444
rect 36237 1417 36271 1444
rect 36271 1417 36280 1444
rect 36228 1372 36280 1405
rect 36228 1353 36237 1372
rect 36237 1353 36271 1372
rect 36271 1353 36280 1372
rect 36228 1338 36237 1341
rect 36237 1338 36271 1341
rect 36271 1338 36280 1341
rect 36228 1300 36280 1338
rect 36228 1289 36237 1300
rect 36237 1289 36271 1300
rect 36271 1289 36280 1300
rect 36228 1266 36237 1277
rect 36237 1266 36271 1277
rect 36271 1266 36280 1277
rect 36228 1228 36280 1266
rect 36228 1225 36237 1228
rect 36237 1225 36271 1228
rect 36271 1225 36280 1228
rect 36228 1194 36237 1213
rect 36237 1194 36271 1213
rect 36271 1194 36280 1213
rect 36228 1161 36280 1194
rect 36324 3100 36376 3133
rect 36324 3081 36333 3100
rect 36333 3081 36367 3100
rect 36367 3081 36376 3100
rect 36324 3066 36333 3069
rect 36333 3066 36367 3069
rect 36367 3066 36376 3069
rect 36324 3028 36376 3066
rect 36324 3017 36333 3028
rect 36333 3017 36367 3028
rect 36367 3017 36376 3028
rect 36324 2994 36333 3005
rect 36333 2994 36367 3005
rect 36367 2994 36376 3005
rect 36324 2956 36376 2994
rect 36324 2953 36333 2956
rect 36333 2953 36367 2956
rect 36367 2953 36376 2956
rect 36324 2922 36333 2941
rect 36333 2922 36367 2941
rect 36367 2922 36376 2941
rect 36324 2889 36376 2922
rect 36324 2850 36333 2877
rect 36333 2850 36367 2877
rect 36367 2850 36376 2877
rect 36324 2825 36376 2850
rect 36324 2812 36376 2813
rect 36324 2778 36333 2812
rect 36333 2778 36367 2812
rect 36367 2778 36376 2812
rect 36324 2761 36376 2778
rect 36324 2740 36376 2749
rect 36324 2706 36333 2740
rect 36333 2706 36367 2740
rect 36367 2706 36376 2740
rect 36324 2697 36376 2706
rect 36324 2668 36376 2685
rect 36324 2634 36333 2668
rect 36333 2634 36367 2668
rect 36367 2634 36376 2668
rect 36324 2633 36376 2634
rect 36324 2596 36376 2621
rect 36324 2569 36333 2596
rect 36333 2569 36367 2596
rect 36367 2569 36376 2596
rect 36324 2524 36376 2557
rect 36324 2505 36333 2524
rect 36333 2505 36367 2524
rect 36367 2505 36376 2524
rect 36324 2490 36333 2493
rect 36333 2490 36367 2493
rect 36367 2490 36376 2493
rect 36324 2452 36376 2490
rect 36324 2441 36333 2452
rect 36333 2441 36367 2452
rect 36367 2441 36376 2452
rect 36324 2418 36333 2429
rect 36333 2418 36367 2429
rect 36367 2418 36376 2429
rect 36324 2380 36376 2418
rect 36324 2377 36333 2380
rect 36333 2377 36367 2380
rect 36367 2377 36376 2380
rect 36324 2346 36333 2365
rect 36333 2346 36367 2365
rect 36367 2346 36376 2365
rect 36324 2313 36376 2346
rect 36324 2274 36333 2301
rect 36333 2274 36367 2301
rect 36367 2274 36376 2301
rect 36324 2249 36376 2274
rect 36324 2236 36376 2237
rect 36324 2202 36333 2236
rect 36333 2202 36367 2236
rect 36367 2202 36376 2236
rect 36324 2185 36376 2202
rect 36324 2164 36376 2173
rect 36324 2130 36333 2164
rect 36333 2130 36367 2164
rect 36367 2130 36376 2164
rect 36324 2121 36376 2130
rect 36324 2092 36376 2109
rect 36324 2058 36333 2092
rect 36333 2058 36367 2092
rect 36367 2058 36376 2092
rect 36324 2057 36376 2058
rect 36324 2020 36376 2045
rect 36324 1993 36333 2020
rect 36333 1993 36367 2020
rect 36367 1993 36376 2020
rect 36324 1948 36376 1981
rect 36324 1929 36333 1948
rect 36333 1929 36367 1948
rect 36367 1929 36376 1948
rect 36324 1914 36333 1917
rect 36333 1914 36367 1917
rect 36367 1914 36376 1917
rect 36324 1876 36376 1914
rect 36324 1865 36333 1876
rect 36333 1865 36367 1876
rect 36367 1865 36376 1876
rect 36324 1842 36333 1853
rect 36333 1842 36367 1853
rect 36367 1842 36376 1853
rect 36324 1804 36376 1842
rect 36324 1801 36333 1804
rect 36333 1801 36367 1804
rect 36367 1801 36376 1804
rect 36324 1770 36333 1789
rect 36333 1770 36367 1789
rect 36367 1770 36376 1789
rect 36324 1737 36376 1770
rect 36324 1698 36333 1725
rect 36333 1698 36367 1725
rect 36367 1698 36376 1725
rect 36324 1673 36376 1698
rect 36324 1660 36376 1661
rect 36324 1626 36333 1660
rect 36333 1626 36367 1660
rect 36367 1626 36376 1660
rect 36324 1609 36376 1626
rect 36324 1588 36376 1597
rect 36324 1554 36333 1588
rect 36333 1554 36367 1588
rect 36367 1554 36376 1588
rect 36324 1545 36376 1554
rect 36324 1516 36376 1533
rect 36324 1482 36333 1516
rect 36333 1482 36367 1516
rect 36367 1482 36376 1516
rect 36324 1481 36376 1482
rect 36324 1444 36376 1469
rect 36324 1417 36333 1444
rect 36333 1417 36367 1444
rect 36367 1417 36376 1444
rect 36324 1372 36376 1405
rect 36324 1353 36333 1372
rect 36333 1353 36367 1372
rect 36367 1353 36376 1372
rect 36324 1338 36333 1341
rect 36333 1338 36367 1341
rect 36367 1338 36376 1341
rect 36324 1300 36376 1338
rect 36324 1289 36333 1300
rect 36333 1289 36367 1300
rect 36367 1289 36376 1300
rect 36324 1266 36333 1277
rect 36333 1266 36367 1277
rect 36367 1266 36376 1277
rect 36324 1228 36376 1266
rect 36324 1225 36333 1228
rect 36333 1225 36367 1228
rect 36367 1225 36376 1228
rect 36324 1194 36333 1213
rect 36333 1194 36367 1213
rect 36367 1194 36376 1213
rect 36324 1161 36376 1194
rect 36420 3100 36472 3133
rect 36420 3081 36429 3100
rect 36429 3081 36463 3100
rect 36463 3081 36472 3100
rect 36420 3066 36429 3069
rect 36429 3066 36463 3069
rect 36463 3066 36472 3069
rect 36420 3028 36472 3066
rect 36420 3017 36429 3028
rect 36429 3017 36463 3028
rect 36463 3017 36472 3028
rect 36420 2994 36429 3005
rect 36429 2994 36463 3005
rect 36463 2994 36472 3005
rect 36420 2956 36472 2994
rect 36420 2953 36429 2956
rect 36429 2953 36463 2956
rect 36463 2953 36472 2956
rect 36420 2922 36429 2941
rect 36429 2922 36463 2941
rect 36463 2922 36472 2941
rect 36420 2889 36472 2922
rect 36420 2850 36429 2877
rect 36429 2850 36463 2877
rect 36463 2850 36472 2877
rect 36420 2825 36472 2850
rect 36420 2812 36472 2813
rect 36420 2778 36429 2812
rect 36429 2778 36463 2812
rect 36463 2778 36472 2812
rect 36420 2761 36472 2778
rect 36420 2740 36472 2749
rect 36420 2706 36429 2740
rect 36429 2706 36463 2740
rect 36463 2706 36472 2740
rect 36420 2697 36472 2706
rect 36420 2668 36472 2685
rect 36420 2634 36429 2668
rect 36429 2634 36463 2668
rect 36463 2634 36472 2668
rect 36420 2633 36472 2634
rect 36420 2596 36472 2621
rect 36420 2569 36429 2596
rect 36429 2569 36463 2596
rect 36463 2569 36472 2596
rect 36420 2524 36472 2557
rect 36420 2505 36429 2524
rect 36429 2505 36463 2524
rect 36463 2505 36472 2524
rect 36420 2490 36429 2493
rect 36429 2490 36463 2493
rect 36463 2490 36472 2493
rect 36420 2452 36472 2490
rect 36420 2441 36429 2452
rect 36429 2441 36463 2452
rect 36463 2441 36472 2452
rect 36420 2418 36429 2429
rect 36429 2418 36463 2429
rect 36463 2418 36472 2429
rect 36420 2380 36472 2418
rect 36420 2377 36429 2380
rect 36429 2377 36463 2380
rect 36463 2377 36472 2380
rect 36420 2346 36429 2365
rect 36429 2346 36463 2365
rect 36463 2346 36472 2365
rect 36420 2313 36472 2346
rect 36420 2274 36429 2301
rect 36429 2274 36463 2301
rect 36463 2274 36472 2301
rect 36420 2249 36472 2274
rect 36420 2236 36472 2237
rect 36420 2202 36429 2236
rect 36429 2202 36463 2236
rect 36463 2202 36472 2236
rect 36420 2185 36472 2202
rect 36420 2164 36472 2173
rect 36420 2130 36429 2164
rect 36429 2130 36463 2164
rect 36463 2130 36472 2164
rect 36420 2121 36472 2130
rect 36420 2092 36472 2109
rect 36420 2058 36429 2092
rect 36429 2058 36463 2092
rect 36463 2058 36472 2092
rect 36420 2057 36472 2058
rect 36420 2020 36472 2045
rect 36420 1993 36429 2020
rect 36429 1993 36463 2020
rect 36463 1993 36472 2020
rect 36420 1948 36472 1981
rect 36420 1929 36429 1948
rect 36429 1929 36463 1948
rect 36463 1929 36472 1948
rect 36420 1914 36429 1917
rect 36429 1914 36463 1917
rect 36463 1914 36472 1917
rect 36420 1876 36472 1914
rect 36420 1865 36429 1876
rect 36429 1865 36463 1876
rect 36463 1865 36472 1876
rect 36420 1842 36429 1853
rect 36429 1842 36463 1853
rect 36463 1842 36472 1853
rect 36420 1804 36472 1842
rect 36420 1801 36429 1804
rect 36429 1801 36463 1804
rect 36463 1801 36472 1804
rect 36420 1770 36429 1789
rect 36429 1770 36463 1789
rect 36463 1770 36472 1789
rect 36420 1737 36472 1770
rect 36420 1698 36429 1725
rect 36429 1698 36463 1725
rect 36463 1698 36472 1725
rect 36420 1673 36472 1698
rect 36420 1660 36472 1661
rect 36420 1626 36429 1660
rect 36429 1626 36463 1660
rect 36463 1626 36472 1660
rect 36420 1609 36472 1626
rect 36420 1588 36472 1597
rect 36420 1554 36429 1588
rect 36429 1554 36463 1588
rect 36463 1554 36472 1588
rect 36420 1545 36472 1554
rect 36420 1516 36472 1533
rect 36420 1482 36429 1516
rect 36429 1482 36463 1516
rect 36463 1482 36472 1516
rect 36420 1481 36472 1482
rect 36420 1444 36472 1469
rect 36420 1417 36429 1444
rect 36429 1417 36463 1444
rect 36463 1417 36472 1444
rect 36420 1372 36472 1405
rect 36420 1353 36429 1372
rect 36429 1353 36463 1372
rect 36463 1353 36472 1372
rect 36420 1338 36429 1341
rect 36429 1338 36463 1341
rect 36463 1338 36472 1341
rect 36420 1300 36472 1338
rect 36420 1289 36429 1300
rect 36429 1289 36463 1300
rect 36463 1289 36472 1300
rect 36420 1266 36429 1277
rect 36429 1266 36463 1277
rect 36463 1266 36472 1277
rect 36420 1228 36472 1266
rect 36420 1225 36429 1228
rect 36429 1225 36463 1228
rect 36463 1225 36472 1228
rect 36420 1194 36429 1213
rect 36429 1194 36463 1213
rect 36463 1194 36472 1213
rect 36420 1161 36472 1194
rect 36516 3100 36568 3133
rect 36516 3081 36525 3100
rect 36525 3081 36559 3100
rect 36559 3081 36568 3100
rect 36516 3066 36525 3069
rect 36525 3066 36559 3069
rect 36559 3066 36568 3069
rect 36516 3028 36568 3066
rect 36516 3017 36525 3028
rect 36525 3017 36559 3028
rect 36559 3017 36568 3028
rect 36516 2994 36525 3005
rect 36525 2994 36559 3005
rect 36559 2994 36568 3005
rect 36516 2956 36568 2994
rect 36516 2953 36525 2956
rect 36525 2953 36559 2956
rect 36559 2953 36568 2956
rect 36516 2922 36525 2941
rect 36525 2922 36559 2941
rect 36559 2922 36568 2941
rect 36516 2889 36568 2922
rect 36516 2850 36525 2877
rect 36525 2850 36559 2877
rect 36559 2850 36568 2877
rect 36516 2825 36568 2850
rect 36516 2812 36568 2813
rect 36516 2778 36525 2812
rect 36525 2778 36559 2812
rect 36559 2778 36568 2812
rect 36516 2761 36568 2778
rect 36516 2740 36568 2749
rect 36516 2706 36525 2740
rect 36525 2706 36559 2740
rect 36559 2706 36568 2740
rect 36516 2697 36568 2706
rect 36516 2668 36568 2685
rect 36516 2634 36525 2668
rect 36525 2634 36559 2668
rect 36559 2634 36568 2668
rect 36516 2633 36568 2634
rect 36516 2596 36568 2621
rect 36516 2569 36525 2596
rect 36525 2569 36559 2596
rect 36559 2569 36568 2596
rect 36516 2524 36568 2557
rect 36516 2505 36525 2524
rect 36525 2505 36559 2524
rect 36559 2505 36568 2524
rect 36516 2490 36525 2493
rect 36525 2490 36559 2493
rect 36559 2490 36568 2493
rect 36516 2452 36568 2490
rect 36516 2441 36525 2452
rect 36525 2441 36559 2452
rect 36559 2441 36568 2452
rect 36516 2418 36525 2429
rect 36525 2418 36559 2429
rect 36559 2418 36568 2429
rect 36516 2380 36568 2418
rect 36516 2377 36525 2380
rect 36525 2377 36559 2380
rect 36559 2377 36568 2380
rect 36516 2346 36525 2365
rect 36525 2346 36559 2365
rect 36559 2346 36568 2365
rect 36516 2313 36568 2346
rect 36516 2274 36525 2301
rect 36525 2274 36559 2301
rect 36559 2274 36568 2301
rect 36516 2249 36568 2274
rect 36516 2236 36568 2237
rect 36516 2202 36525 2236
rect 36525 2202 36559 2236
rect 36559 2202 36568 2236
rect 36516 2185 36568 2202
rect 36516 2164 36568 2173
rect 36516 2130 36525 2164
rect 36525 2130 36559 2164
rect 36559 2130 36568 2164
rect 36516 2121 36568 2130
rect 36516 2092 36568 2109
rect 36516 2058 36525 2092
rect 36525 2058 36559 2092
rect 36559 2058 36568 2092
rect 36516 2057 36568 2058
rect 36516 2020 36568 2045
rect 36516 1993 36525 2020
rect 36525 1993 36559 2020
rect 36559 1993 36568 2020
rect 36516 1948 36568 1981
rect 36516 1929 36525 1948
rect 36525 1929 36559 1948
rect 36559 1929 36568 1948
rect 36516 1914 36525 1917
rect 36525 1914 36559 1917
rect 36559 1914 36568 1917
rect 36516 1876 36568 1914
rect 36516 1865 36525 1876
rect 36525 1865 36559 1876
rect 36559 1865 36568 1876
rect 36516 1842 36525 1853
rect 36525 1842 36559 1853
rect 36559 1842 36568 1853
rect 36516 1804 36568 1842
rect 36516 1801 36525 1804
rect 36525 1801 36559 1804
rect 36559 1801 36568 1804
rect 36516 1770 36525 1789
rect 36525 1770 36559 1789
rect 36559 1770 36568 1789
rect 36516 1737 36568 1770
rect 36516 1698 36525 1725
rect 36525 1698 36559 1725
rect 36559 1698 36568 1725
rect 36516 1673 36568 1698
rect 36516 1660 36568 1661
rect 36516 1626 36525 1660
rect 36525 1626 36559 1660
rect 36559 1626 36568 1660
rect 36516 1609 36568 1626
rect 36516 1588 36568 1597
rect 36516 1554 36525 1588
rect 36525 1554 36559 1588
rect 36559 1554 36568 1588
rect 36516 1545 36568 1554
rect 36516 1516 36568 1533
rect 36516 1482 36525 1516
rect 36525 1482 36559 1516
rect 36559 1482 36568 1516
rect 36516 1481 36568 1482
rect 36516 1444 36568 1469
rect 36516 1417 36525 1444
rect 36525 1417 36559 1444
rect 36559 1417 36568 1444
rect 36516 1372 36568 1405
rect 36516 1353 36525 1372
rect 36525 1353 36559 1372
rect 36559 1353 36568 1372
rect 36516 1338 36525 1341
rect 36525 1338 36559 1341
rect 36559 1338 36568 1341
rect 36516 1300 36568 1338
rect 36516 1289 36525 1300
rect 36525 1289 36559 1300
rect 36559 1289 36568 1300
rect 36516 1266 36525 1277
rect 36525 1266 36559 1277
rect 36559 1266 36568 1277
rect 36516 1228 36568 1266
rect 36516 1225 36525 1228
rect 36525 1225 36559 1228
rect 36559 1225 36568 1228
rect 36516 1194 36525 1213
rect 36525 1194 36559 1213
rect 36559 1194 36568 1213
rect 36516 1161 36568 1194
rect 36612 3100 36664 3133
rect 36612 3081 36621 3100
rect 36621 3081 36655 3100
rect 36655 3081 36664 3100
rect 36612 3066 36621 3069
rect 36621 3066 36655 3069
rect 36655 3066 36664 3069
rect 36612 3028 36664 3066
rect 36612 3017 36621 3028
rect 36621 3017 36655 3028
rect 36655 3017 36664 3028
rect 36612 2994 36621 3005
rect 36621 2994 36655 3005
rect 36655 2994 36664 3005
rect 36612 2956 36664 2994
rect 36612 2953 36621 2956
rect 36621 2953 36655 2956
rect 36655 2953 36664 2956
rect 36612 2922 36621 2941
rect 36621 2922 36655 2941
rect 36655 2922 36664 2941
rect 36612 2889 36664 2922
rect 36612 2850 36621 2877
rect 36621 2850 36655 2877
rect 36655 2850 36664 2877
rect 36612 2825 36664 2850
rect 36612 2812 36664 2813
rect 36612 2778 36621 2812
rect 36621 2778 36655 2812
rect 36655 2778 36664 2812
rect 36612 2761 36664 2778
rect 36612 2740 36664 2749
rect 36612 2706 36621 2740
rect 36621 2706 36655 2740
rect 36655 2706 36664 2740
rect 36612 2697 36664 2706
rect 36612 2668 36664 2685
rect 36612 2634 36621 2668
rect 36621 2634 36655 2668
rect 36655 2634 36664 2668
rect 36612 2633 36664 2634
rect 36612 2596 36664 2621
rect 36612 2569 36621 2596
rect 36621 2569 36655 2596
rect 36655 2569 36664 2596
rect 36612 2524 36664 2557
rect 36612 2505 36621 2524
rect 36621 2505 36655 2524
rect 36655 2505 36664 2524
rect 36612 2490 36621 2493
rect 36621 2490 36655 2493
rect 36655 2490 36664 2493
rect 36612 2452 36664 2490
rect 36612 2441 36621 2452
rect 36621 2441 36655 2452
rect 36655 2441 36664 2452
rect 36612 2418 36621 2429
rect 36621 2418 36655 2429
rect 36655 2418 36664 2429
rect 36612 2380 36664 2418
rect 36612 2377 36621 2380
rect 36621 2377 36655 2380
rect 36655 2377 36664 2380
rect 36612 2346 36621 2365
rect 36621 2346 36655 2365
rect 36655 2346 36664 2365
rect 36612 2313 36664 2346
rect 36612 2274 36621 2301
rect 36621 2274 36655 2301
rect 36655 2274 36664 2301
rect 36612 2249 36664 2274
rect 36612 2236 36664 2237
rect 36612 2202 36621 2236
rect 36621 2202 36655 2236
rect 36655 2202 36664 2236
rect 36612 2185 36664 2202
rect 36612 2164 36664 2173
rect 36612 2130 36621 2164
rect 36621 2130 36655 2164
rect 36655 2130 36664 2164
rect 36612 2121 36664 2130
rect 36612 2092 36664 2109
rect 36612 2058 36621 2092
rect 36621 2058 36655 2092
rect 36655 2058 36664 2092
rect 36612 2057 36664 2058
rect 36612 2020 36664 2045
rect 36612 1993 36621 2020
rect 36621 1993 36655 2020
rect 36655 1993 36664 2020
rect 36612 1948 36664 1981
rect 36612 1929 36621 1948
rect 36621 1929 36655 1948
rect 36655 1929 36664 1948
rect 36612 1914 36621 1917
rect 36621 1914 36655 1917
rect 36655 1914 36664 1917
rect 36612 1876 36664 1914
rect 36612 1865 36621 1876
rect 36621 1865 36655 1876
rect 36655 1865 36664 1876
rect 36612 1842 36621 1853
rect 36621 1842 36655 1853
rect 36655 1842 36664 1853
rect 36612 1804 36664 1842
rect 36612 1801 36621 1804
rect 36621 1801 36655 1804
rect 36655 1801 36664 1804
rect 36612 1770 36621 1789
rect 36621 1770 36655 1789
rect 36655 1770 36664 1789
rect 36612 1737 36664 1770
rect 36612 1698 36621 1725
rect 36621 1698 36655 1725
rect 36655 1698 36664 1725
rect 36612 1673 36664 1698
rect 36612 1660 36664 1661
rect 36612 1626 36621 1660
rect 36621 1626 36655 1660
rect 36655 1626 36664 1660
rect 36612 1609 36664 1626
rect 36612 1588 36664 1597
rect 36612 1554 36621 1588
rect 36621 1554 36655 1588
rect 36655 1554 36664 1588
rect 36612 1545 36664 1554
rect 36612 1516 36664 1533
rect 36612 1482 36621 1516
rect 36621 1482 36655 1516
rect 36655 1482 36664 1516
rect 36612 1481 36664 1482
rect 36612 1444 36664 1469
rect 36612 1417 36621 1444
rect 36621 1417 36655 1444
rect 36655 1417 36664 1444
rect 36612 1372 36664 1405
rect 36612 1353 36621 1372
rect 36621 1353 36655 1372
rect 36655 1353 36664 1372
rect 36612 1338 36621 1341
rect 36621 1338 36655 1341
rect 36655 1338 36664 1341
rect 36612 1300 36664 1338
rect 36612 1289 36621 1300
rect 36621 1289 36655 1300
rect 36655 1289 36664 1300
rect 36612 1266 36621 1277
rect 36621 1266 36655 1277
rect 36655 1266 36664 1277
rect 36612 1228 36664 1266
rect 36612 1225 36621 1228
rect 36621 1225 36655 1228
rect 36655 1225 36664 1228
rect 36612 1194 36621 1213
rect 36621 1194 36655 1213
rect 36655 1194 36664 1213
rect 36612 1161 36664 1194
rect 36708 3100 36760 3133
rect 36708 3081 36717 3100
rect 36717 3081 36751 3100
rect 36751 3081 36760 3100
rect 36708 3066 36717 3069
rect 36717 3066 36751 3069
rect 36751 3066 36760 3069
rect 36708 3028 36760 3066
rect 36708 3017 36717 3028
rect 36717 3017 36751 3028
rect 36751 3017 36760 3028
rect 36708 2994 36717 3005
rect 36717 2994 36751 3005
rect 36751 2994 36760 3005
rect 36708 2956 36760 2994
rect 36708 2953 36717 2956
rect 36717 2953 36751 2956
rect 36751 2953 36760 2956
rect 36708 2922 36717 2941
rect 36717 2922 36751 2941
rect 36751 2922 36760 2941
rect 36708 2889 36760 2922
rect 36708 2850 36717 2877
rect 36717 2850 36751 2877
rect 36751 2850 36760 2877
rect 36708 2825 36760 2850
rect 36708 2812 36760 2813
rect 36708 2778 36717 2812
rect 36717 2778 36751 2812
rect 36751 2778 36760 2812
rect 36708 2761 36760 2778
rect 36708 2740 36760 2749
rect 36708 2706 36717 2740
rect 36717 2706 36751 2740
rect 36751 2706 36760 2740
rect 36708 2697 36760 2706
rect 36708 2668 36760 2685
rect 36708 2634 36717 2668
rect 36717 2634 36751 2668
rect 36751 2634 36760 2668
rect 36708 2633 36760 2634
rect 36708 2596 36760 2621
rect 36708 2569 36717 2596
rect 36717 2569 36751 2596
rect 36751 2569 36760 2596
rect 36708 2524 36760 2557
rect 36708 2505 36717 2524
rect 36717 2505 36751 2524
rect 36751 2505 36760 2524
rect 36708 2490 36717 2493
rect 36717 2490 36751 2493
rect 36751 2490 36760 2493
rect 36708 2452 36760 2490
rect 36708 2441 36717 2452
rect 36717 2441 36751 2452
rect 36751 2441 36760 2452
rect 36708 2418 36717 2429
rect 36717 2418 36751 2429
rect 36751 2418 36760 2429
rect 36708 2380 36760 2418
rect 36708 2377 36717 2380
rect 36717 2377 36751 2380
rect 36751 2377 36760 2380
rect 36708 2346 36717 2365
rect 36717 2346 36751 2365
rect 36751 2346 36760 2365
rect 36708 2313 36760 2346
rect 36708 2274 36717 2301
rect 36717 2274 36751 2301
rect 36751 2274 36760 2301
rect 36708 2249 36760 2274
rect 36708 2236 36760 2237
rect 36708 2202 36717 2236
rect 36717 2202 36751 2236
rect 36751 2202 36760 2236
rect 36708 2185 36760 2202
rect 36708 2164 36760 2173
rect 36708 2130 36717 2164
rect 36717 2130 36751 2164
rect 36751 2130 36760 2164
rect 36708 2121 36760 2130
rect 36708 2092 36760 2109
rect 36708 2058 36717 2092
rect 36717 2058 36751 2092
rect 36751 2058 36760 2092
rect 36708 2057 36760 2058
rect 36708 2020 36760 2045
rect 36708 1993 36717 2020
rect 36717 1993 36751 2020
rect 36751 1993 36760 2020
rect 36708 1948 36760 1981
rect 36708 1929 36717 1948
rect 36717 1929 36751 1948
rect 36751 1929 36760 1948
rect 36708 1914 36717 1917
rect 36717 1914 36751 1917
rect 36751 1914 36760 1917
rect 36708 1876 36760 1914
rect 36708 1865 36717 1876
rect 36717 1865 36751 1876
rect 36751 1865 36760 1876
rect 36708 1842 36717 1853
rect 36717 1842 36751 1853
rect 36751 1842 36760 1853
rect 36708 1804 36760 1842
rect 36708 1801 36717 1804
rect 36717 1801 36751 1804
rect 36751 1801 36760 1804
rect 36708 1770 36717 1789
rect 36717 1770 36751 1789
rect 36751 1770 36760 1789
rect 36708 1737 36760 1770
rect 36708 1698 36717 1725
rect 36717 1698 36751 1725
rect 36751 1698 36760 1725
rect 36708 1673 36760 1698
rect 36708 1660 36760 1661
rect 36708 1626 36717 1660
rect 36717 1626 36751 1660
rect 36751 1626 36760 1660
rect 36708 1609 36760 1626
rect 36708 1588 36760 1597
rect 36708 1554 36717 1588
rect 36717 1554 36751 1588
rect 36751 1554 36760 1588
rect 36708 1545 36760 1554
rect 36708 1516 36760 1533
rect 36708 1482 36717 1516
rect 36717 1482 36751 1516
rect 36751 1482 36760 1516
rect 36708 1481 36760 1482
rect 36708 1444 36760 1469
rect 36708 1417 36717 1444
rect 36717 1417 36751 1444
rect 36751 1417 36760 1444
rect 36708 1372 36760 1405
rect 36708 1353 36717 1372
rect 36717 1353 36751 1372
rect 36751 1353 36760 1372
rect 36708 1338 36717 1341
rect 36717 1338 36751 1341
rect 36751 1338 36760 1341
rect 36708 1300 36760 1338
rect 36708 1289 36717 1300
rect 36717 1289 36751 1300
rect 36751 1289 36760 1300
rect 36708 1266 36717 1277
rect 36717 1266 36751 1277
rect 36751 1266 36760 1277
rect 36708 1228 36760 1266
rect 36708 1225 36717 1228
rect 36717 1225 36751 1228
rect 36751 1225 36760 1228
rect 36708 1194 36717 1213
rect 36717 1194 36751 1213
rect 36751 1194 36760 1213
rect 36708 1161 36760 1194
rect 36804 3100 36856 3133
rect 36804 3081 36813 3100
rect 36813 3081 36847 3100
rect 36847 3081 36856 3100
rect 36804 3066 36813 3069
rect 36813 3066 36847 3069
rect 36847 3066 36856 3069
rect 36804 3028 36856 3066
rect 36804 3017 36813 3028
rect 36813 3017 36847 3028
rect 36847 3017 36856 3028
rect 36804 2994 36813 3005
rect 36813 2994 36847 3005
rect 36847 2994 36856 3005
rect 36804 2956 36856 2994
rect 36804 2953 36813 2956
rect 36813 2953 36847 2956
rect 36847 2953 36856 2956
rect 36804 2922 36813 2941
rect 36813 2922 36847 2941
rect 36847 2922 36856 2941
rect 36804 2889 36856 2922
rect 36804 2850 36813 2877
rect 36813 2850 36847 2877
rect 36847 2850 36856 2877
rect 36804 2825 36856 2850
rect 36804 2812 36856 2813
rect 36804 2778 36813 2812
rect 36813 2778 36847 2812
rect 36847 2778 36856 2812
rect 36804 2761 36856 2778
rect 36804 2740 36856 2749
rect 36804 2706 36813 2740
rect 36813 2706 36847 2740
rect 36847 2706 36856 2740
rect 36804 2697 36856 2706
rect 36804 2668 36856 2685
rect 36804 2634 36813 2668
rect 36813 2634 36847 2668
rect 36847 2634 36856 2668
rect 36804 2633 36856 2634
rect 36804 2596 36856 2621
rect 36804 2569 36813 2596
rect 36813 2569 36847 2596
rect 36847 2569 36856 2596
rect 36804 2524 36856 2557
rect 36804 2505 36813 2524
rect 36813 2505 36847 2524
rect 36847 2505 36856 2524
rect 36804 2490 36813 2493
rect 36813 2490 36847 2493
rect 36847 2490 36856 2493
rect 36804 2452 36856 2490
rect 36804 2441 36813 2452
rect 36813 2441 36847 2452
rect 36847 2441 36856 2452
rect 36804 2418 36813 2429
rect 36813 2418 36847 2429
rect 36847 2418 36856 2429
rect 36804 2380 36856 2418
rect 36804 2377 36813 2380
rect 36813 2377 36847 2380
rect 36847 2377 36856 2380
rect 36804 2346 36813 2365
rect 36813 2346 36847 2365
rect 36847 2346 36856 2365
rect 36804 2313 36856 2346
rect 36804 2274 36813 2301
rect 36813 2274 36847 2301
rect 36847 2274 36856 2301
rect 36804 2249 36856 2274
rect 36804 2236 36856 2237
rect 36804 2202 36813 2236
rect 36813 2202 36847 2236
rect 36847 2202 36856 2236
rect 36804 2185 36856 2202
rect 36804 2164 36856 2173
rect 36804 2130 36813 2164
rect 36813 2130 36847 2164
rect 36847 2130 36856 2164
rect 36804 2121 36856 2130
rect 36804 2092 36856 2109
rect 36804 2058 36813 2092
rect 36813 2058 36847 2092
rect 36847 2058 36856 2092
rect 36804 2057 36856 2058
rect 36804 2020 36856 2045
rect 36804 1993 36813 2020
rect 36813 1993 36847 2020
rect 36847 1993 36856 2020
rect 36804 1948 36856 1981
rect 36804 1929 36813 1948
rect 36813 1929 36847 1948
rect 36847 1929 36856 1948
rect 36804 1914 36813 1917
rect 36813 1914 36847 1917
rect 36847 1914 36856 1917
rect 36804 1876 36856 1914
rect 36804 1865 36813 1876
rect 36813 1865 36847 1876
rect 36847 1865 36856 1876
rect 36804 1842 36813 1853
rect 36813 1842 36847 1853
rect 36847 1842 36856 1853
rect 36804 1804 36856 1842
rect 36804 1801 36813 1804
rect 36813 1801 36847 1804
rect 36847 1801 36856 1804
rect 36804 1770 36813 1789
rect 36813 1770 36847 1789
rect 36847 1770 36856 1789
rect 36804 1737 36856 1770
rect 36804 1698 36813 1725
rect 36813 1698 36847 1725
rect 36847 1698 36856 1725
rect 36804 1673 36856 1698
rect 36804 1660 36856 1661
rect 36804 1626 36813 1660
rect 36813 1626 36847 1660
rect 36847 1626 36856 1660
rect 36804 1609 36856 1626
rect 36804 1588 36856 1597
rect 36804 1554 36813 1588
rect 36813 1554 36847 1588
rect 36847 1554 36856 1588
rect 36804 1545 36856 1554
rect 36804 1516 36856 1533
rect 36804 1482 36813 1516
rect 36813 1482 36847 1516
rect 36847 1482 36856 1516
rect 36804 1481 36856 1482
rect 36804 1444 36856 1469
rect 36804 1417 36813 1444
rect 36813 1417 36847 1444
rect 36847 1417 36856 1444
rect 36804 1372 36856 1405
rect 36804 1353 36813 1372
rect 36813 1353 36847 1372
rect 36847 1353 36856 1372
rect 36804 1338 36813 1341
rect 36813 1338 36847 1341
rect 36847 1338 36856 1341
rect 36804 1300 36856 1338
rect 36804 1289 36813 1300
rect 36813 1289 36847 1300
rect 36847 1289 36856 1300
rect 36804 1266 36813 1277
rect 36813 1266 36847 1277
rect 36847 1266 36856 1277
rect 36804 1228 36856 1266
rect 36804 1225 36813 1228
rect 36813 1225 36847 1228
rect 36847 1225 36856 1228
rect 36804 1194 36813 1213
rect 36813 1194 36847 1213
rect 36847 1194 36856 1213
rect 36804 1161 36856 1194
rect 36900 3100 36952 3133
rect 36900 3081 36909 3100
rect 36909 3081 36943 3100
rect 36943 3081 36952 3100
rect 36900 3066 36909 3069
rect 36909 3066 36943 3069
rect 36943 3066 36952 3069
rect 36900 3028 36952 3066
rect 36900 3017 36909 3028
rect 36909 3017 36943 3028
rect 36943 3017 36952 3028
rect 36900 2994 36909 3005
rect 36909 2994 36943 3005
rect 36943 2994 36952 3005
rect 36900 2956 36952 2994
rect 36900 2953 36909 2956
rect 36909 2953 36943 2956
rect 36943 2953 36952 2956
rect 36900 2922 36909 2941
rect 36909 2922 36943 2941
rect 36943 2922 36952 2941
rect 36900 2889 36952 2922
rect 36900 2850 36909 2877
rect 36909 2850 36943 2877
rect 36943 2850 36952 2877
rect 36900 2825 36952 2850
rect 36900 2812 36952 2813
rect 36900 2778 36909 2812
rect 36909 2778 36943 2812
rect 36943 2778 36952 2812
rect 36900 2761 36952 2778
rect 36900 2740 36952 2749
rect 36900 2706 36909 2740
rect 36909 2706 36943 2740
rect 36943 2706 36952 2740
rect 36900 2697 36952 2706
rect 36900 2668 36952 2685
rect 36900 2634 36909 2668
rect 36909 2634 36943 2668
rect 36943 2634 36952 2668
rect 36900 2633 36952 2634
rect 36900 2596 36952 2621
rect 36900 2569 36909 2596
rect 36909 2569 36943 2596
rect 36943 2569 36952 2596
rect 36900 2524 36952 2557
rect 36900 2505 36909 2524
rect 36909 2505 36943 2524
rect 36943 2505 36952 2524
rect 36900 2490 36909 2493
rect 36909 2490 36943 2493
rect 36943 2490 36952 2493
rect 36900 2452 36952 2490
rect 36900 2441 36909 2452
rect 36909 2441 36943 2452
rect 36943 2441 36952 2452
rect 36900 2418 36909 2429
rect 36909 2418 36943 2429
rect 36943 2418 36952 2429
rect 36900 2380 36952 2418
rect 36900 2377 36909 2380
rect 36909 2377 36943 2380
rect 36943 2377 36952 2380
rect 36900 2346 36909 2365
rect 36909 2346 36943 2365
rect 36943 2346 36952 2365
rect 36900 2313 36952 2346
rect 36900 2274 36909 2301
rect 36909 2274 36943 2301
rect 36943 2274 36952 2301
rect 36900 2249 36952 2274
rect 36900 2236 36952 2237
rect 36900 2202 36909 2236
rect 36909 2202 36943 2236
rect 36943 2202 36952 2236
rect 36900 2185 36952 2202
rect 36900 2164 36952 2173
rect 36900 2130 36909 2164
rect 36909 2130 36943 2164
rect 36943 2130 36952 2164
rect 36900 2121 36952 2130
rect 36900 2092 36952 2109
rect 36900 2058 36909 2092
rect 36909 2058 36943 2092
rect 36943 2058 36952 2092
rect 36900 2057 36952 2058
rect 36900 2020 36952 2045
rect 36900 1993 36909 2020
rect 36909 1993 36943 2020
rect 36943 1993 36952 2020
rect 36900 1948 36952 1981
rect 36900 1929 36909 1948
rect 36909 1929 36943 1948
rect 36943 1929 36952 1948
rect 36900 1914 36909 1917
rect 36909 1914 36943 1917
rect 36943 1914 36952 1917
rect 36900 1876 36952 1914
rect 36900 1865 36909 1876
rect 36909 1865 36943 1876
rect 36943 1865 36952 1876
rect 36900 1842 36909 1853
rect 36909 1842 36943 1853
rect 36943 1842 36952 1853
rect 36900 1804 36952 1842
rect 36900 1801 36909 1804
rect 36909 1801 36943 1804
rect 36943 1801 36952 1804
rect 36900 1770 36909 1789
rect 36909 1770 36943 1789
rect 36943 1770 36952 1789
rect 36900 1737 36952 1770
rect 36900 1698 36909 1725
rect 36909 1698 36943 1725
rect 36943 1698 36952 1725
rect 36900 1673 36952 1698
rect 36900 1660 36952 1661
rect 36900 1626 36909 1660
rect 36909 1626 36943 1660
rect 36943 1626 36952 1660
rect 36900 1609 36952 1626
rect 36900 1588 36952 1597
rect 36900 1554 36909 1588
rect 36909 1554 36943 1588
rect 36943 1554 36952 1588
rect 36900 1545 36952 1554
rect 36900 1516 36952 1533
rect 36900 1482 36909 1516
rect 36909 1482 36943 1516
rect 36943 1482 36952 1516
rect 36900 1481 36952 1482
rect 36900 1444 36952 1469
rect 36900 1417 36909 1444
rect 36909 1417 36943 1444
rect 36943 1417 36952 1444
rect 36900 1372 36952 1405
rect 36900 1353 36909 1372
rect 36909 1353 36943 1372
rect 36943 1353 36952 1372
rect 36900 1338 36909 1341
rect 36909 1338 36943 1341
rect 36943 1338 36952 1341
rect 36900 1300 36952 1338
rect 36900 1289 36909 1300
rect 36909 1289 36943 1300
rect 36943 1289 36952 1300
rect 36900 1266 36909 1277
rect 36909 1266 36943 1277
rect 36943 1266 36952 1277
rect 36900 1228 36952 1266
rect 36900 1225 36909 1228
rect 36909 1225 36943 1228
rect 36943 1225 36952 1228
rect 36900 1194 36909 1213
rect 36909 1194 36943 1213
rect 36943 1194 36952 1213
rect 36900 1161 36952 1194
rect 36996 3100 37048 3133
rect 36996 3081 37005 3100
rect 37005 3081 37039 3100
rect 37039 3081 37048 3100
rect 36996 3066 37005 3069
rect 37005 3066 37039 3069
rect 37039 3066 37048 3069
rect 36996 3028 37048 3066
rect 36996 3017 37005 3028
rect 37005 3017 37039 3028
rect 37039 3017 37048 3028
rect 36996 2994 37005 3005
rect 37005 2994 37039 3005
rect 37039 2994 37048 3005
rect 36996 2956 37048 2994
rect 36996 2953 37005 2956
rect 37005 2953 37039 2956
rect 37039 2953 37048 2956
rect 36996 2922 37005 2941
rect 37005 2922 37039 2941
rect 37039 2922 37048 2941
rect 36996 2889 37048 2922
rect 36996 2850 37005 2877
rect 37005 2850 37039 2877
rect 37039 2850 37048 2877
rect 36996 2825 37048 2850
rect 36996 2812 37048 2813
rect 36996 2778 37005 2812
rect 37005 2778 37039 2812
rect 37039 2778 37048 2812
rect 36996 2761 37048 2778
rect 36996 2740 37048 2749
rect 36996 2706 37005 2740
rect 37005 2706 37039 2740
rect 37039 2706 37048 2740
rect 36996 2697 37048 2706
rect 36996 2668 37048 2685
rect 36996 2634 37005 2668
rect 37005 2634 37039 2668
rect 37039 2634 37048 2668
rect 36996 2633 37048 2634
rect 36996 2596 37048 2621
rect 36996 2569 37005 2596
rect 37005 2569 37039 2596
rect 37039 2569 37048 2596
rect 36996 2524 37048 2557
rect 36996 2505 37005 2524
rect 37005 2505 37039 2524
rect 37039 2505 37048 2524
rect 36996 2490 37005 2493
rect 37005 2490 37039 2493
rect 37039 2490 37048 2493
rect 36996 2452 37048 2490
rect 36996 2441 37005 2452
rect 37005 2441 37039 2452
rect 37039 2441 37048 2452
rect 36996 2418 37005 2429
rect 37005 2418 37039 2429
rect 37039 2418 37048 2429
rect 36996 2380 37048 2418
rect 36996 2377 37005 2380
rect 37005 2377 37039 2380
rect 37039 2377 37048 2380
rect 36996 2346 37005 2365
rect 37005 2346 37039 2365
rect 37039 2346 37048 2365
rect 36996 2313 37048 2346
rect 36996 2274 37005 2301
rect 37005 2274 37039 2301
rect 37039 2274 37048 2301
rect 36996 2249 37048 2274
rect 36996 2236 37048 2237
rect 36996 2202 37005 2236
rect 37005 2202 37039 2236
rect 37039 2202 37048 2236
rect 36996 2185 37048 2202
rect 36996 2164 37048 2173
rect 36996 2130 37005 2164
rect 37005 2130 37039 2164
rect 37039 2130 37048 2164
rect 36996 2121 37048 2130
rect 36996 2092 37048 2109
rect 36996 2058 37005 2092
rect 37005 2058 37039 2092
rect 37039 2058 37048 2092
rect 36996 2057 37048 2058
rect 36996 2020 37048 2045
rect 36996 1993 37005 2020
rect 37005 1993 37039 2020
rect 37039 1993 37048 2020
rect 36996 1948 37048 1981
rect 36996 1929 37005 1948
rect 37005 1929 37039 1948
rect 37039 1929 37048 1948
rect 36996 1914 37005 1917
rect 37005 1914 37039 1917
rect 37039 1914 37048 1917
rect 36996 1876 37048 1914
rect 36996 1865 37005 1876
rect 37005 1865 37039 1876
rect 37039 1865 37048 1876
rect 36996 1842 37005 1853
rect 37005 1842 37039 1853
rect 37039 1842 37048 1853
rect 36996 1804 37048 1842
rect 36996 1801 37005 1804
rect 37005 1801 37039 1804
rect 37039 1801 37048 1804
rect 36996 1770 37005 1789
rect 37005 1770 37039 1789
rect 37039 1770 37048 1789
rect 36996 1737 37048 1770
rect 36996 1698 37005 1725
rect 37005 1698 37039 1725
rect 37039 1698 37048 1725
rect 36996 1673 37048 1698
rect 36996 1660 37048 1661
rect 36996 1626 37005 1660
rect 37005 1626 37039 1660
rect 37039 1626 37048 1660
rect 36996 1609 37048 1626
rect 36996 1588 37048 1597
rect 36996 1554 37005 1588
rect 37005 1554 37039 1588
rect 37039 1554 37048 1588
rect 36996 1545 37048 1554
rect 36996 1516 37048 1533
rect 36996 1482 37005 1516
rect 37005 1482 37039 1516
rect 37039 1482 37048 1516
rect 36996 1481 37048 1482
rect 36996 1444 37048 1469
rect 36996 1417 37005 1444
rect 37005 1417 37039 1444
rect 37039 1417 37048 1444
rect 36996 1372 37048 1405
rect 36996 1353 37005 1372
rect 37005 1353 37039 1372
rect 37039 1353 37048 1372
rect 36996 1338 37005 1341
rect 37005 1338 37039 1341
rect 37039 1338 37048 1341
rect 36996 1300 37048 1338
rect 36996 1289 37005 1300
rect 37005 1289 37039 1300
rect 37039 1289 37048 1300
rect 36996 1266 37005 1277
rect 37005 1266 37039 1277
rect 37039 1266 37048 1277
rect 36996 1228 37048 1266
rect 36996 1225 37005 1228
rect 37005 1225 37039 1228
rect 37039 1225 37048 1228
rect 36996 1194 37005 1213
rect 37005 1194 37039 1213
rect 37039 1194 37048 1213
rect 36996 1161 37048 1194
rect 37092 3100 37144 3133
rect 37092 3081 37101 3100
rect 37101 3081 37135 3100
rect 37135 3081 37144 3100
rect 37092 3066 37101 3069
rect 37101 3066 37135 3069
rect 37135 3066 37144 3069
rect 37092 3028 37144 3066
rect 37092 3017 37101 3028
rect 37101 3017 37135 3028
rect 37135 3017 37144 3028
rect 37092 2994 37101 3005
rect 37101 2994 37135 3005
rect 37135 2994 37144 3005
rect 37092 2956 37144 2994
rect 37092 2953 37101 2956
rect 37101 2953 37135 2956
rect 37135 2953 37144 2956
rect 37092 2922 37101 2941
rect 37101 2922 37135 2941
rect 37135 2922 37144 2941
rect 37092 2889 37144 2922
rect 37092 2850 37101 2877
rect 37101 2850 37135 2877
rect 37135 2850 37144 2877
rect 37092 2825 37144 2850
rect 37092 2812 37144 2813
rect 37092 2778 37101 2812
rect 37101 2778 37135 2812
rect 37135 2778 37144 2812
rect 37092 2761 37144 2778
rect 37092 2740 37144 2749
rect 37092 2706 37101 2740
rect 37101 2706 37135 2740
rect 37135 2706 37144 2740
rect 37092 2697 37144 2706
rect 37092 2668 37144 2685
rect 37092 2634 37101 2668
rect 37101 2634 37135 2668
rect 37135 2634 37144 2668
rect 37092 2633 37144 2634
rect 37092 2596 37144 2621
rect 37092 2569 37101 2596
rect 37101 2569 37135 2596
rect 37135 2569 37144 2596
rect 37092 2524 37144 2557
rect 37092 2505 37101 2524
rect 37101 2505 37135 2524
rect 37135 2505 37144 2524
rect 37092 2490 37101 2493
rect 37101 2490 37135 2493
rect 37135 2490 37144 2493
rect 37092 2452 37144 2490
rect 37092 2441 37101 2452
rect 37101 2441 37135 2452
rect 37135 2441 37144 2452
rect 37092 2418 37101 2429
rect 37101 2418 37135 2429
rect 37135 2418 37144 2429
rect 37092 2380 37144 2418
rect 37092 2377 37101 2380
rect 37101 2377 37135 2380
rect 37135 2377 37144 2380
rect 37092 2346 37101 2365
rect 37101 2346 37135 2365
rect 37135 2346 37144 2365
rect 37092 2313 37144 2346
rect 37092 2274 37101 2301
rect 37101 2274 37135 2301
rect 37135 2274 37144 2301
rect 37092 2249 37144 2274
rect 37092 2236 37144 2237
rect 37092 2202 37101 2236
rect 37101 2202 37135 2236
rect 37135 2202 37144 2236
rect 37092 2185 37144 2202
rect 37092 2164 37144 2173
rect 37092 2130 37101 2164
rect 37101 2130 37135 2164
rect 37135 2130 37144 2164
rect 37092 2121 37144 2130
rect 37092 2092 37144 2109
rect 37092 2058 37101 2092
rect 37101 2058 37135 2092
rect 37135 2058 37144 2092
rect 37092 2057 37144 2058
rect 37092 2020 37144 2045
rect 37092 1993 37101 2020
rect 37101 1993 37135 2020
rect 37135 1993 37144 2020
rect 37092 1948 37144 1981
rect 37092 1929 37101 1948
rect 37101 1929 37135 1948
rect 37135 1929 37144 1948
rect 37092 1914 37101 1917
rect 37101 1914 37135 1917
rect 37135 1914 37144 1917
rect 37092 1876 37144 1914
rect 37092 1865 37101 1876
rect 37101 1865 37135 1876
rect 37135 1865 37144 1876
rect 37092 1842 37101 1853
rect 37101 1842 37135 1853
rect 37135 1842 37144 1853
rect 37092 1804 37144 1842
rect 37092 1801 37101 1804
rect 37101 1801 37135 1804
rect 37135 1801 37144 1804
rect 37092 1770 37101 1789
rect 37101 1770 37135 1789
rect 37135 1770 37144 1789
rect 37092 1737 37144 1770
rect 37092 1698 37101 1725
rect 37101 1698 37135 1725
rect 37135 1698 37144 1725
rect 37092 1673 37144 1698
rect 37092 1660 37144 1661
rect 37092 1626 37101 1660
rect 37101 1626 37135 1660
rect 37135 1626 37144 1660
rect 37092 1609 37144 1626
rect 37092 1588 37144 1597
rect 37092 1554 37101 1588
rect 37101 1554 37135 1588
rect 37135 1554 37144 1588
rect 37092 1545 37144 1554
rect 37092 1516 37144 1533
rect 37092 1482 37101 1516
rect 37101 1482 37135 1516
rect 37135 1482 37144 1516
rect 37092 1481 37144 1482
rect 37092 1444 37144 1469
rect 37092 1417 37101 1444
rect 37101 1417 37135 1444
rect 37135 1417 37144 1444
rect 37092 1372 37144 1405
rect 37092 1353 37101 1372
rect 37101 1353 37135 1372
rect 37135 1353 37144 1372
rect 37092 1338 37101 1341
rect 37101 1338 37135 1341
rect 37135 1338 37144 1341
rect 37092 1300 37144 1338
rect 37092 1289 37101 1300
rect 37101 1289 37135 1300
rect 37135 1289 37144 1300
rect 37092 1266 37101 1277
rect 37101 1266 37135 1277
rect 37135 1266 37144 1277
rect 37092 1228 37144 1266
rect 37092 1225 37101 1228
rect 37101 1225 37135 1228
rect 37135 1225 37144 1228
rect 37092 1194 37101 1213
rect 37101 1194 37135 1213
rect 37135 1194 37144 1213
rect 37092 1161 37144 1194
rect 37188 3100 37240 3133
rect 37188 3081 37197 3100
rect 37197 3081 37231 3100
rect 37231 3081 37240 3100
rect 37188 3066 37197 3069
rect 37197 3066 37231 3069
rect 37231 3066 37240 3069
rect 37188 3028 37240 3066
rect 37188 3017 37197 3028
rect 37197 3017 37231 3028
rect 37231 3017 37240 3028
rect 37188 2994 37197 3005
rect 37197 2994 37231 3005
rect 37231 2994 37240 3005
rect 37188 2956 37240 2994
rect 37188 2953 37197 2956
rect 37197 2953 37231 2956
rect 37231 2953 37240 2956
rect 37188 2922 37197 2941
rect 37197 2922 37231 2941
rect 37231 2922 37240 2941
rect 37188 2889 37240 2922
rect 37188 2850 37197 2877
rect 37197 2850 37231 2877
rect 37231 2850 37240 2877
rect 37188 2825 37240 2850
rect 37188 2812 37240 2813
rect 37188 2778 37197 2812
rect 37197 2778 37231 2812
rect 37231 2778 37240 2812
rect 37188 2761 37240 2778
rect 37188 2740 37240 2749
rect 37188 2706 37197 2740
rect 37197 2706 37231 2740
rect 37231 2706 37240 2740
rect 37188 2697 37240 2706
rect 37188 2668 37240 2685
rect 37188 2634 37197 2668
rect 37197 2634 37231 2668
rect 37231 2634 37240 2668
rect 37188 2633 37240 2634
rect 37188 2596 37240 2621
rect 37188 2569 37197 2596
rect 37197 2569 37231 2596
rect 37231 2569 37240 2596
rect 37188 2524 37240 2557
rect 37188 2505 37197 2524
rect 37197 2505 37231 2524
rect 37231 2505 37240 2524
rect 37188 2490 37197 2493
rect 37197 2490 37231 2493
rect 37231 2490 37240 2493
rect 37188 2452 37240 2490
rect 37188 2441 37197 2452
rect 37197 2441 37231 2452
rect 37231 2441 37240 2452
rect 37188 2418 37197 2429
rect 37197 2418 37231 2429
rect 37231 2418 37240 2429
rect 37188 2380 37240 2418
rect 37188 2377 37197 2380
rect 37197 2377 37231 2380
rect 37231 2377 37240 2380
rect 37188 2346 37197 2365
rect 37197 2346 37231 2365
rect 37231 2346 37240 2365
rect 37188 2313 37240 2346
rect 37188 2274 37197 2301
rect 37197 2274 37231 2301
rect 37231 2274 37240 2301
rect 37188 2249 37240 2274
rect 37188 2236 37240 2237
rect 37188 2202 37197 2236
rect 37197 2202 37231 2236
rect 37231 2202 37240 2236
rect 37188 2185 37240 2202
rect 37188 2164 37240 2173
rect 37188 2130 37197 2164
rect 37197 2130 37231 2164
rect 37231 2130 37240 2164
rect 37188 2121 37240 2130
rect 37188 2092 37240 2109
rect 37188 2058 37197 2092
rect 37197 2058 37231 2092
rect 37231 2058 37240 2092
rect 37188 2057 37240 2058
rect 37188 2020 37240 2045
rect 37188 1993 37197 2020
rect 37197 1993 37231 2020
rect 37231 1993 37240 2020
rect 37188 1948 37240 1981
rect 37188 1929 37197 1948
rect 37197 1929 37231 1948
rect 37231 1929 37240 1948
rect 37188 1914 37197 1917
rect 37197 1914 37231 1917
rect 37231 1914 37240 1917
rect 37188 1876 37240 1914
rect 37188 1865 37197 1876
rect 37197 1865 37231 1876
rect 37231 1865 37240 1876
rect 37188 1842 37197 1853
rect 37197 1842 37231 1853
rect 37231 1842 37240 1853
rect 37188 1804 37240 1842
rect 37188 1801 37197 1804
rect 37197 1801 37231 1804
rect 37231 1801 37240 1804
rect 37188 1770 37197 1789
rect 37197 1770 37231 1789
rect 37231 1770 37240 1789
rect 37188 1737 37240 1770
rect 37188 1698 37197 1725
rect 37197 1698 37231 1725
rect 37231 1698 37240 1725
rect 37188 1673 37240 1698
rect 37188 1660 37240 1661
rect 37188 1626 37197 1660
rect 37197 1626 37231 1660
rect 37231 1626 37240 1660
rect 37188 1609 37240 1626
rect 37188 1588 37240 1597
rect 37188 1554 37197 1588
rect 37197 1554 37231 1588
rect 37231 1554 37240 1588
rect 37188 1545 37240 1554
rect 37188 1516 37240 1533
rect 37188 1482 37197 1516
rect 37197 1482 37231 1516
rect 37231 1482 37240 1516
rect 37188 1481 37240 1482
rect 37188 1444 37240 1469
rect 37188 1417 37197 1444
rect 37197 1417 37231 1444
rect 37231 1417 37240 1444
rect 37188 1372 37240 1405
rect 37188 1353 37197 1372
rect 37197 1353 37231 1372
rect 37231 1353 37240 1372
rect 37188 1338 37197 1341
rect 37197 1338 37231 1341
rect 37231 1338 37240 1341
rect 37188 1300 37240 1338
rect 37188 1289 37197 1300
rect 37197 1289 37231 1300
rect 37231 1289 37240 1300
rect 37188 1266 37197 1277
rect 37197 1266 37231 1277
rect 37231 1266 37240 1277
rect 37188 1228 37240 1266
rect 37188 1225 37197 1228
rect 37197 1225 37231 1228
rect 37231 1225 37240 1228
rect 37188 1194 37197 1213
rect 37197 1194 37231 1213
rect 37231 1194 37240 1213
rect 37188 1161 37240 1194
rect 37284 3100 37336 3133
rect 37284 3081 37293 3100
rect 37293 3081 37327 3100
rect 37327 3081 37336 3100
rect 37284 3066 37293 3069
rect 37293 3066 37327 3069
rect 37327 3066 37336 3069
rect 37284 3028 37336 3066
rect 37284 3017 37293 3028
rect 37293 3017 37327 3028
rect 37327 3017 37336 3028
rect 37284 2994 37293 3005
rect 37293 2994 37327 3005
rect 37327 2994 37336 3005
rect 37284 2956 37336 2994
rect 37284 2953 37293 2956
rect 37293 2953 37327 2956
rect 37327 2953 37336 2956
rect 37284 2922 37293 2941
rect 37293 2922 37327 2941
rect 37327 2922 37336 2941
rect 37284 2889 37336 2922
rect 37284 2850 37293 2877
rect 37293 2850 37327 2877
rect 37327 2850 37336 2877
rect 37284 2825 37336 2850
rect 37284 2812 37336 2813
rect 37284 2778 37293 2812
rect 37293 2778 37327 2812
rect 37327 2778 37336 2812
rect 37284 2761 37336 2778
rect 37284 2740 37336 2749
rect 37284 2706 37293 2740
rect 37293 2706 37327 2740
rect 37327 2706 37336 2740
rect 37284 2697 37336 2706
rect 37284 2668 37336 2685
rect 37284 2634 37293 2668
rect 37293 2634 37327 2668
rect 37327 2634 37336 2668
rect 37284 2633 37336 2634
rect 37284 2596 37336 2621
rect 37284 2569 37293 2596
rect 37293 2569 37327 2596
rect 37327 2569 37336 2596
rect 37284 2524 37336 2557
rect 37284 2505 37293 2524
rect 37293 2505 37327 2524
rect 37327 2505 37336 2524
rect 37284 2490 37293 2493
rect 37293 2490 37327 2493
rect 37327 2490 37336 2493
rect 37284 2452 37336 2490
rect 37284 2441 37293 2452
rect 37293 2441 37327 2452
rect 37327 2441 37336 2452
rect 37284 2418 37293 2429
rect 37293 2418 37327 2429
rect 37327 2418 37336 2429
rect 37284 2380 37336 2418
rect 37284 2377 37293 2380
rect 37293 2377 37327 2380
rect 37327 2377 37336 2380
rect 37284 2346 37293 2365
rect 37293 2346 37327 2365
rect 37327 2346 37336 2365
rect 37284 2313 37336 2346
rect 37284 2274 37293 2301
rect 37293 2274 37327 2301
rect 37327 2274 37336 2301
rect 37284 2249 37336 2274
rect 37284 2236 37336 2237
rect 37284 2202 37293 2236
rect 37293 2202 37327 2236
rect 37327 2202 37336 2236
rect 37284 2185 37336 2202
rect 37284 2164 37336 2173
rect 37284 2130 37293 2164
rect 37293 2130 37327 2164
rect 37327 2130 37336 2164
rect 37284 2121 37336 2130
rect 37284 2092 37336 2109
rect 37284 2058 37293 2092
rect 37293 2058 37327 2092
rect 37327 2058 37336 2092
rect 37284 2057 37336 2058
rect 37284 2020 37336 2045
rect 37284 1993 37293 2020
rect 37293 1993 37327 2020
rect 37327 1993 37336 2020
rect 37284 1948 37336 1981
rect 37284 1929 37293 1948
rect 37293 1929 37327 1948
rect 37327 1929 37336 1948
rect 37284 1914 37293 1917
rect 37293 1914 37327 1917
rect 37327 1914 37336 1917
rect 37284 1876 37336 1914
rect 37284 1865 37293 1876
rect 37293 1865 37327 1876
rect 37327 1865 37336 1876
rect 37284 1842 37293 1853
rect 37293 1842 37327 1853
rect 37327 1842 37336 1853
rect 37284 1804 37336 1842
rect 37284 1801 37293 1804
rect 37293 1801 37327 1804
rect 37327 1801 37336 1804
rect 37284 1770 37293 1789
rect 37293 1770 37327 1789
rect 37327 1770 37336 1789
rect 37284 1737 37336 1770
rect 37284 1698 37293 1725
rect 37293 1698 37327 1725
rect 37327 1698 37336 1725
rect 37284 1673 37336 1698
rect 37284 1660 37336 1661
rect 37284 1626 37293 1660
rect 37293 1626 37327 1660
rect 37327 1626 37336 1660
rect 37284 1609 37336 1626
rect 37284 1588 37336 1597
rect 37284 1554 37293 1588
rect 37293 1554 37327 1588
rect 37327 1554 37336 1588
rect 37284 1545 37336 1554
rect 37284 1516 37336 1533
rect 37284 1482 37293 1516
rect 37293 1482 37327 1516
rect 37327 1482 37336 1516
rect 37284 1481 37336 1482
rect 37284 1444 37336 1469
rect 37284 1417 37293 1444
rect 37293 1417 37327 1444
rect 37327 1417 37336 1444
rect 37284 1372 37336 1405
rect 37284 1353 37293 1372
rect 37293 1353 37327 1372
rect 37327 1353 37336 1372
rect 37284 1338 37293 1341
rect 37293 1338 37327 1341
rect 37327 1338 37336 1341
rect 37284 1300 37336 1338
rect 37284 1289 37293 1300
rect 37293 1289 37327 1300
rect 37327 1289 37336 1300
rect 37284 1266 37293 1277
rect 37293 1266 37327 1277
rect 37327 1266 37336 1277
rect 37284 1228 37336 1266
rect 37284 1225 37293 1228
rect 37293 1225 37327 1228
rect 37327 1225 37336 1228
rect 37284 1194 37293 1213
rect 37293 1194 37327 1213
rect 37327 1194 37336 1213
rect 37284 1161 37336 1194
rect 37380 3100 37432 3133
rect 37380 3081 37389 3100
rect 37389 3081 37423 3100
rect 37423 3081 37432 3100
rect 37380 3066 37389 3069
rect 37389 3066 37423 3069
rect 37423 3066 37432 3069
rect 37380 3028 37432 3066
rect 37380 3017 37389 3028
rect 37389 3017 37423 3028
rect 37423 3017 37432 3028
rect 37380 2994 37389 3005
rect 37389 2994 37423 3005
rect 37423 2994 37432 3005
rect 37380 2956 37432 2994
rect 37380 2953 37389 2956
rect 37389 2953 37423 2956
rect 37423 2953 37432 2956
rect 37380 2922 37389 2941
rect 37389 2922 37423 2941
rect 37423 2922 37432 2941
rect 37380 2889 37432 2922
rect 37380 2850 37389 2877
rect 37389 2850 37423 2877
rect 37423 2850 37432 2877
rect 37380 2825 37432 2850
rect 37380 2812 37432 2813
rect 37380 2778 37389 2812
rect 37389 2778 37423 2812
rect 37423 2778 37432 2812
rect 37380 2761 37432 2778
rect 37380 2740 37432 2749
rect 37380 2706 37389 2740
rect 37389 2706 37423 2740
rect 37423 2706 37432 2740
rect 37380 2697 37432 2706
rect 37380 2668 37432 2685
rect 37380 2634 37389 2668
rect 37389 2634 37423 2668
rect 37423 2634 37432 2668
rect 37380 2633 37432 2634
rect 37380 2596 37432 2621
rect 37380 2569 37389 2596
rect 37389 2569 37423 2596
rect 37423 2569 37432 2596
rect 37380 2524 37432 2557
rect 37380 2505 37389 2524
rect 37389 2505 37423 2524
rect 37423 2505 37432 2524
rect 37380 2490 37389 2493
rect 37389 2490 37423 2493
rect 37423 2490 37432 2493
rect 37380 2452 37432 2490
rect 37380 2441 37389 2452
rect 37389 2441 37423 2452
rect 37423 2441 37432 2452
rect 37380 2418 37389 2429
rect 37389 2418 37423 2429
rect 37423 2418 37432 2429
rect 37380 2380 37432 2418
rect 37380 2377 37389 2380
rect 37389 2377 37423 2380
rect 37423 2377 37432 2380
rect 37380 2346 37389 2365
rect 37389 2346 37423 2365
rect 37423 2346 37432 2365
rect 37380 2313 37432 2346
rect 37380 2274 37389 2301
rect 37389 2274 37423 2301
rect 37423 2274 37432 2301
rect 37380 2249 37432 2274
rect 37380 2236 37432 2237
rect 37380 2202 37389 2236
rect 37389 2202 37423 2236
rect 37423 2202 37432 2236
rect 37380 2185 37432 2202
rect 37380 2164 37432 2173
rect 37380 2130 37389 2164
rect 37389 2130 37423 2164
rect 37423 2130 37432 2164
rect 37380 2121 37432 2130
rect 37380 2092 37432 2109
rect 37380 2058 37389 2092
rect 37389 2058 37423 2092
rect 37423 2058 37432 2092
rect 37380 2057 37432 2058
rect 37380 2020 37432 2045
rect 37380 1993 37389 2020
rect 37389 1993 37423 2020
rect 37423 1993 37432 2020
rect 37380 1948 37432 1981
rect 37380 1929 37389 1948
rect 37389 1929 37423 1948
rect 37423 1929 37432 1948
rect 37380 1914 37389 1917
rect 37389 1914 37423 1917
rect 37423 1914 37432 1917
rect 37380 1876 37432 1914
rect 37380 1865 37389 1876
rect 37389 1865 37423 1876
rect 37423 1865 37432 1876
rect 37380 1842 37389 1853
rect 37389 1842 37423 1853
rect 37423 1842 37432 1853
rect 37380 1804 37432 1842
rect 37380 1801 37389 1804
rect 37389 1801 37423 1804
rect 37423 1801 37432 1804
rect 37380 1770 37389 1789
rect 37389 1770 37423 1789
rect 37423 1770 37432 1789
rect 37380 1737 37432 1770
rect 37380 1698 37389 1725
rect 37389 1698 37423 1725
rect 37423 1698 37432 1725
rect 37380 1673 37432 1698
rect 37380 1660 37432 1661
rect 37380 1626 37389 1660
rect 37389 1626 37423 1660
rect 37423 1626 37432 1660
rect 37380 1609 37432 1626
rect 37380 1588 37432 1597
rect 37380 1554 37389 1588
rect 37389 1554 37423 1588
rect 37423 1554 37432 1588
rect 37380 1545 37432 1554
rect 37380 1516 37432 1533
rect 37380 1482 37389 1516
rect 37389 1482 37423 1516
rect 37423 1482 37432 1516
rect 37380 1481 37432 1482
rect 37380 1444 37432 1469
rect 37380 1417 37389 1444
rect 37389 1417 37423 1444
rect 37423 1417 37432 1444
rect 37380 1372 37432 1405
rect 37380 1353 37389 1372
rect 37389 1353 37423 1372
rect 37423 1353 37432 1372
rect 37380 1338 37389 1341
rect 37389 1338 37423 1341
rect 37423 1338 37432 1341
rect 37380 1300 37432 1338
rect 37380 1289 37389 1300
rect 37389 1289 37423 1300
rect 37423 1289 37432 1300
rect 37380 1266 37389 1277
rect 37389 1266 37423 1277
rect 37423 1266 37432 1277
rect 37380 1228 37432 1266
rect 37380 1225 37389 1228
rect 37389 1225 37423 1228
rect 37423 1225 37432 1228
rect 37380 1194 37389 1213
rect 37389 1194 37423 1213
rect 37423 1194 37432 1213
rect 37380 1161 37432 1194
rect 37476 3100 37528 3133
rect 37476 3081 37485 3100
rect 37485 3081 37519 3100
rect 37519 3081 37528 3100
rect 37476 3066 37485 3069
rect 37485 3066 37519 3069
rect 37519 3066 37528 3069
rect 37476 3028 37528 3066
rect 37476 3017 37485 3028
rect 37485 3017 37519 3028
rect 37519 3017 37528 3028
rect 37476 2994 37485 3005
rect 37485 2994 37519 3005
rect 37519 2994 37528 3005
rect 37476 2956 37528 2994
rect 37476 2953 37485 2956
rect 37485 2953 37519 2956
rect 37519 2953 37528 2956
rect 37476 2922 37485 2941
rect 37485 2922 37519 2941
rect 37519 2922 37528 2941
rect 37476 2889 37528 2922
rect 37476 2850 37485 2877
rect 37485 2850 37519 2877
rect 37519 2850 37528 2877
rect 37476 2825 37528 2850
rect 37476 2812 37528 2813
rect 37476 2778 37485 2812
rect 37485 2778 37519 2812
rect 37519 2778 37528 2812
rect 37476 2761 37528 2778
rect 37476 2740 37528 2749
rect 37476 2706 37485 2740
rect 37485 2706 37519 2740
rect 37519 2706 37528 2740
rect 37476 2697 37528 2706
rect 37476 2668 37528 2685
rect 37476 2634 37485 2668
rect 37485 2634 37519 2668
rect 37519 2634 37528 2668
rect 37476 2633 37528 2634
rect 37476 2596 37528 2621
rect 37476 2569 37485 2596
rect 37485 2569 37519 2596
rect 37519 2569 37528 2596
rect 37476 2524 37528 2557
rect 37476 2505 37485 2524
rect 37485 2505 37519 2524
rect 37519 2505 37528 2524
rect 37476 2490 37485 2493
rect 37485 2490 37519 2493
rect 37519 2490 37528 2493
rect 37476 2452 37528 2490
rect 37476 2441 37485 2452
rect 37485 2441 37519 2452
rect 37519 2441 37528 2452
rect 37476 2418 37485 2429
rect 37485 2418 37519 2429
rect 37519 2418 37528 2429
rect 37476 2380 37528 2418
rect 37476 2377 37485 2380
rect 37485 2377 37519 2380
rect 37519 2377 37528 2380
rect 37476 2346 37485 2365
rect 37485 2346 37519 2365
rect 37519 2346 37528 2365
rect 37476 2313 37528 2346
rect 37476 2274 37485 2301
rect 37485 2274 37519 2301
rect 37519 2274 37528 2301
rect 37476 2249 37528 2274
rect 37476 2236 37528 2237
rect 37476 2202 37485 2236
rect 37485 2202 37519 2236
rect 37519 2202 37528 2236
rect 37476 2185 37528 2202
rect 37476 2164 37528 2173
rect 37476 2130 37485 2164
rect 37485 2130 37519 2164
rect 37519 2130 37528 2164
rect 37476 2121 37528 2130
rect 37476 2092 37528 2109
rect 37476 2058 37485 2092
rect 37485 2058 37519 2092
rect 37519 2058 37528 2092
rect 37476 2057 37528 2058
rect 37476 2020 37528 2045
rect 37476 1993 37485 2020
rect 37485 1993 37519 2020
rect 37519 1993 37528 2020
rect 37476 1948 37528 1981
rect 37476 1929 37485 1948
rect 37485 1929 37519 1948
rect 37519 1929 37528 1948
rect 37476 1914 37485 1917
rect 37485 1914 37519 1917
rect 37519 1914 37528 1917
rect 37476 1876 37528 1914
rect 37476 1865 37485 1876
rect 37485 1865 37519 1876
rect 37519 1865 37528 1876
rect 37476 1842 37485 1853
rect 37485 1842 37519 1853
rect 37519 1842 37528 1853
rect 37476 1804 37528 1842
rect 37476 1801 37485 1804
rect 37485 1801 37519 1804
rect 37519 1801 37528 1804
rect 37476 1770 37485 1789
rect 37485 1770 37519 1789
rect 37519 1770 37528 1789
rect 37476 1737 37528 1770
rect 37476 1698 37485 1725
rect 37485 1698 37519 1725
rect 37519 1698 37528 1725
rect 37476 1673 37528 1698
rect 37476 1660 37528 1661
rect 37476 1626 37485 1660
rect 37485 1626 37519 1660
rect 37519 1626 37528 1660
rect 37476 1609 37528 1626
rect 37476 1588 37528 1597
rect 37476 1554 37485 1588
rect 37485 1554 37519 1588
rect 37519 1554 37528 1588
rect 37476 1545 37528 1554
rect 37476 1516 37528 1533
rect 37476 1482 37485 1516
rect 37485 1482 37519 1516
rect 37519 1482 37528 1516
rect 37476 1481 37528 1482
rect 37476 1444 37528 1469
rect 37476 1417 37485 1444
rect 37485 1417 37519 1444
rect 37519 1417 37528 1444
rect 37476 1372 37528 1405
rect 37476 1353 37485 1372
rect 37485 1353 37519 1372
rect 37519 1353 37528 1372
rect 37476 1338 37485 1341
rect 37485 1338 37519 1341
rect 37519 1338 37528 1341
rect 37476 1300 37528 1338
rect 37476 1289 37485 1300
rect 37485 1289 37519 1300
rect 37519 1289 37528 1300
rect 37476 1266 37485 1277
rect 37485 1266 37519 1277
rect 37519 1266 37528 1277
rect 37476 1228 37528 1266
rect 37476 1225 37485 1228
rect 37485 1225 37519 1228
rect 37519 1225 37528 1228
rect 37476 1194 37485 1213
rect 37485 1194 37519 1213
rect 37519 1194 37528 1213
rect 37476 1161 37528 1194
rect 37572 3100 37624 3133
rect 37572 3081 37581 3100
rect 37581 3081 37615 3100
rect 37615 3081 37624 3100
rect 37572 3066 37581 3069
rect 37581 3066 37615 3069
rect 37615 3066 37624 3069
rect 37572 3028 37624 3066
rect 37572 3017 37581 3028
rect 37581 3017 37615 3028
rect 37615 3017 37624 3028
rect 37572 2994 37581 3005
rect 37581 2994 37615 3005
rect 37615 2994 37624 3005
rect 37572 2956 37624 2994
rect 37572 2953 37581 2956
rect 37581 2953 37615 2956
rect 37615 2953 37624 2956
rect 37572 2922 37581 2941
rect 37581 2922 37615 2941
rect 37615 2922 37624 2941
rect 37572 2889 37624 2922
rect 37572 2850 37581 2877
rect 37581 2850 37615 2877
rect 37615 2850 37624 2877
rect 37572 2825 37624 2850
rect 37572 2812 37624 2813
rect 37572 2778 37581 2812
rect 37581 2778 37615 2812
rect 37615 2778 37624 2812
rect 37572 2761 37624 2778
rect 37572 2740 37624 2749
rect 37572 2706 37581 2740
rect 37581 2706 37615 2740
rect 37615 2706 37624 2740
rect 37572 2697 37624 2706
rect 37572 2668 37624 2685
rect 37572 2634 37581 2668
rect 37581 2634 37615 2668
rect 37615 2634 37624 2668
rect 37572 2633 37624 2634
rect 37572 2596 37624 2621
rect 37572 2569 37581 2596
rect 37581 2569 37615 2596
rect 37615 2569 37624 2596
rect 37572 2524 37624 2557
rect 37572 2505 37581 2524
rect 37581 2505 37615 2524
rect 37615 2505 37624 2524
rect 37572 2490 37581 2493
rect 37581 2490 37615 2493
rect 37615 2490 37624 2493
rect 37572 2452 37624 2490
rect 37572 2441 37581 2452
rect 37581 2441 37615 2452
rect 37615 2441 37624 2452
rect 37572 2418 37581 2429
rect 37581 2418 37615 2429
rect 37615 2418 37624 2429
rect 37572 2380 37624 2418
rect 37572 2377 37581 2380
rect 37581 2377 37615 2380
rect 37615 2377 37624 2380
rect 37572 2346 37581 2365
rect 37581 2346 37615 2365
rect 37615 2346 37624 2365
rect 37572 2313 37624 2346
rect 37572 2274 37581 2301
rect 37581 2274 37615 2301
rect 37615 2274 37624 2301
rect 37572 2249 37624 2274
rect 37572 2236 37624 2237
rect 37572 2202 37581 2236
rect 37581 2202 37615 2236
rect 37615 2202 37624 2236
rect 37572 2185 37624 2202
rect 37572 2164 37624 2173
rect 37572 2130 37581 2164
rect 37581 2130 37615 2164
rect 37615 2130 37624 2164
rect 37572 2121 37624 2130
rect 37572 2092 37624 2109
rect 37572 2058 37581 2092
rect 37581 2058 37615 2092
rect 37615 2058 37624 2092
rect 37572 2057 37624 2058
rect 37572 2020 37624 2045
rect 37572 1993 37581 2020
rect 37581 1993 37615 2020
rect 37615 1993 37624 2020
rect 37572 1948 37624 1981
rect 37572 1929 37581 1948
rect 37581 1929 37615 1948
rect 37615 1929 37624 1948
rect 37572 1914 37581 1917
rect 37581 1914 37615 1917
rect 37615 1914 37624 1917
rect 37572 1876 37624 1914
rect 37572 1865 37581 1876
rect 37581 1865 37615 1876
rect 37615 1865 37624 1876
rect 37572 1842 37581 1853
rect 37581 1842 37615 1853
rect 37615 1842 37624 1853
rect 37572 1804 37624 1842
rect 37572 1801 37581 1804
rect 37581 1801 37615 1804
rect 37615 1801 37624 1804
rect 37572 1770 37581 1789
rect 37581 1770 37615 1789
rect 37615 1770 37624 1789
rect 37572 1737 37624 1770
rect 37572 1698 37581 1725
rect 37581 1698 37615 1725
rect 37615 1698 37624 1725
rect 37572 1673 37624 1698
rect 37572 1660 37624 1661
rect 37572 1626 37581 1660
rect 37581 1626 37615 1660
rect 37615 1626 37624 1660
rect 37572 1609 37624 1626
rect 37572 1588 37624 1597
rect 37572 1554 37581 1588
rect 37581 1554 37615 1588
rect 37615 1554 37624 1588
rect 37572 1545 37624 1554
rect 37572 1516 37624 1533
rect 37572 1482 37581 1516
rect 37581 1482 37615 1516
rect 37615 1482 37624 1516
rect 37572 1481 37624 1482
rect 37572 1444 37624 1469
rect 37572 1417 37581 1444
rect 37581 1417 37615 1444
rect 37615 1417 37624 1444
rect 37572 1372 37624 1405
rect 37572 1353 37581 1372
rect 37581 1353 37615 1372
rect 37615 1353 37624 1372
rect 37572 1338 37581 1341
rect 37581 1338 37615 1341
rect 37615 1338 37624 1341
rect 37572 1300 37624 1338
rect 37572 1289 37581 1300
rect 37581 1289 37615 1300
rect 37615 1289 37624 1300
rect 37572 1266 37581 1277
rect 37581 1266 37615 1277
rect 37615 1266 37624 1277
rect 37572 1228 37624 1266
rect 37572 1225 37581 1228
rect 37581 1225 37615 1228
rect 37615 1225 37624 1228
rect 37572 1194 37581 1213
rect 37581 1194 37615 1213
rect 37615 1194 37624 1213
rect 37572 1161 37624 1194
rect 37668 3100 37720 3133
rect 37668 3081 37677 3100
rect 37677 3081 37711 3100
rect 37711 3081 37720 3100
rect 37668 3066 37677 3069
rect 37677 3066 37711 3069
rect 37711 3066 37720 3069
rect 37668 3028 37720 3066
rect 37668 3017 37677 3028
rect 37677 3017 37711 3028
rect 37711 3017 37720 3028
rect 37668 2994 37677 3005
rect 37677 2994 37711 3005
rect 37711 2994 37720 3005
rect 37668 2956 37720 2994
rect 37668 2953 37677 2956
rect 37677 2953 37711 2956
rect 37711 2953 37720 2956
rect 37668 2922 37677 2941
rect 37677 2922 37711 2941
rect 37711 2922 37720 2941
rect 37668 2889 37720 2922
rect 37668 2850 37677 2877
rect 37677 2850 37711 2877
rect 37711 2850 37720 2877
rect 37668 2825 37720 2850
rect 37668 2812 37720 2813
rect 37668 2778 37677 2812
rect 37677 2778 37711 2812
rect 37711 2778 37720 2812
rect 37668 2761 37720 2778
rect 37668 2740 37720 2749
rect 37668 2706 37677 2740
rect 37677 2706 37711 2740
rect 37711 2706 37720 2740
rect 37668 2697 37720 2706
rect 37668 2668 37720 2685
rect 37668 2634 37677 2668
rect 37677 2634 37711 2668
rect 37711 2634 37720 2668
rect 37668 2633 37720 2634
rect 37668 2596 37720 2621
rect 37668 2569 37677 2596
rect 37677 2569 37711 2596
rect 37711 2569 37720 2596
rect 37668 2524 37720 2557
rect 37668 2505 37677 2524
rect 37677 2505 37711 2524
rect 37711 2505 37720 2524
rect 37668 2490 37677 2493
rect 37677 2490 37711 2493
rect 37711 2490 37720 2493
rect 37668 2452 37720 2490
rect 37668 2441 37677 2452
rect 37677 2441 37711 2452
rect 37711 2441 37720 2452
rect 37668 2418 37677 2429
rect 37677 2418 37711 2429
rect 37711 2418 37720 2429
rect 37668 2380 37720 2418
rect 37668 2377 37677 2380
rect 37677 2377 37711 2380
rect 37711 2377 37720 2380
rect 37668 2346 37677 2365
rect 37677 2346 37711 2365
rect 37711 2346 37720 2365
rect 37668 2313 37720 2346
rect 37668 2274 37677 2301
rect 37677 2274 37711 2301
rect 37711 2274 37720 2301
rect 37668 2249 37720 2274
rect 37668 2236 37720 2237
rect 37668 2202 37677 2236
rect 37677 2202 37711 2236
rect 37711 2202 37720 2236
rect 37668 2185 37720 2202
rect 37668 2164 37720 2173
rect 37668 2130 37677 2164
rect 37677 2130 37711 2164
rect 37711 2130 37720 2164
rect 37668 2121 37720 2130
rect 37668 2092 37720 2109
rect 37668 2058 37677 2092
rect 37677 2058 37711 2092
rect 37711 2058 37720 2092
rect 37668 2057 37720 2058
rect 37668 2020 37720 2045
rect 37668 1993 37677 2020
rect 37677 1993 37711 2020
rect 37711 1993 37720 2020
rect 37668 1948 37720 1981
rect 37668 1929 37677 1948
rect 37677 1929 37711 1948
rect 37711 1929 37720 1948
rect 37668 1914 37677 1917
rect 37677 1914 37711 1917
rect 37711 1914 37720 1917
rect 37668 1876 37720 1914
rect 37668 1865 37677 1876
rect 37677 1865 37711 1876
rect 37711 1865 37720 1876
rect 37668 1842 37677 1853
rect 37677 1842 37711 1853
rect 37711 1842 37720 1853
rect 37668 1804 37720 1842
rect 37668 1801 37677 1804
rect 37677 1801 37711 1804
rect 37711 1801 37720 1804
rect 37668 1770 37677 1789
rect 37677 1770 37711 1789
rect 37711 1770 37720 1789
rect 37668 1737 37720 1770
rect 37668 1698 37677 1725
rect 37677 1698 37711 1725
rect 37711 1698 37720 1725
rect 37668 1673 37720 1698
rect 37668 1660 37720 1661
rect 37668 1626 37677 1660
rect 37677 1626 37711 1660
rect 37711 1626 37720 1660
rect 37668 1609 37720 1626
rect 37668 1588 37720 1597
rect 37668 1554 37677 1588
rect 37677 1554 37711 1588
rect 37711 1554 37720 1588
rect 37668 1545 37720 1554
rect 37668 1516 37720 1533
rect 37668 1482 37677 1516
rect 37677 1482 37711 1516
rect 37711 1482 37720 1516
rect 37668 1481 37720 1482
rect 37668 1444 37720 1469
rect 37668 1417 37677 1444
rect 37677 1417 37711 1444
rect 37711 1417 37720 1444
rect 37668 1372 37720 1405
rect 37668 1353 37677 1372
rect 37677 1353 37711 1372
rect 37711 1353 37720 1372
rect 37668 1338 37677 1341
rect 37677 1338 37711 1341
rect 37711 1338 37720 1341
rect 37668 1300 37720 1338
rect 37668 1289 37677 1300
rect 37677 1289 37711 1300
rect 37711 1289 37720 1300
rect 37668 1266 37677 1277
rect 37677 1266 37711 1277
rect 37711 1266 37720 1277
rect 37668 1228 37720 1266
rect 37668 1225 37677 1228
rect 37677 1225 37711 1228
rect 37711 1225 37720 1228
rect 37668 1194 37677 1213
rect 37677 1194 37711 1213
rect 37711 1194 37720 1213
rect 37668 1161 37720 1194
rect 37764 3100 37816 3133
rect 37764 3081 37773 3100
rect 37773 3081 37807 3100
rect 37807 3081 37816 3100
rect 37764 3066 37773 3069
rect 37773 3066 37807 3069
rect 37807 3066 37816 3069
rect 37764 3028 37816 3066
rect 37764 3017 37773 3028
rect 37773 3017 37807 3028
rect 37807 3017 37816 3028
rect 37764 2994 37773 3005
rect 37773 2994 37807 3005
rect 37807 2994 37816 3005
rect 37764 2956 37816 2994
rect 37764 2953 37773 2956
rect 37773 2953 37807 2956
rect 37807 2953 37816 2956
rect 37764 2922 37773 2941
rect 37773 2922 37807 2941
rect 37807 2922 37816 2941
rect 37764 2889 37816 2922
rect 37764 2850 37773 2877
rect 37773 2850 37807 2877
rect 37807 2850 37816 2877
rect 37764 2825 37816 2850
rect 37764 2812 37816 2813
rect 37764 2778 37773 2812
rect 37773 2778 37807 2812
rect 37807 2778 37816 2812
rect 37764 2761 37816 2778
rect 37764 2740 37816 2749
rect 37764 2706 37773 2740
rect 37773 2706 37807 2740
rect 37807 2706 37816 2740
rect 37764 2697 37816 2706
rect 37764 2668 37816 2685
rect 37764 2634 37773 2668
rect 37773 2634 37807 2668
rect 37807 2634 37816 2668
rect 37764 2633 37816 2634
rect 37764 2596 37816 2621
rect 37764 2569 37773 2596
rect 37773 2569 37807 2596
rect 37807 2569 37816 2596
rect 37764 2524 37816 2557
rect 37764 2505 37773 2524
rect 37773 2505 37807 2524
rect 37807 2505 37816 2524
rect 37764 2490 37773 2493
rect 37773 2490 37807 2493
rect 37807 2490 37816 2493
rect 37764 2452 37816 2490
rect 37764 2441 37773 2452
rect 37773 2441 37807 2452
rect 37807 2441 37816 2452
rect 37764 2418 37773 2429
rect 37773 2418 37807 2429
rect 37807 2418 37816 2429
rect 37764 2380 37816 2418
rect 37764 2377 37773 2380
rect 37773 2377 37807 2380
rect 37807 2377 37816 2380
rect 37764 2346 37773 2365
rect 37773 2346 37807 2365
rect 37807 2346 37816 2365
rect 37764 2313 37816 2346
rect 37764 2274 37773 2301
rect 37773 2274 37807 2301
rect 37807 2274 37816 2301
rect 37764 2249 37816 2274
rect 37764 2236 37816 2237
rect 37764 2202 37773 2236
rect 37773 2202 37807 2236
rect 37807 2202 37816 2236
rect 37764 2185 37816 2202
rect 37764 2164 37816 2173
rect 37764 2130 37773 2164
rect 37773 2130 37807 2164
rect 37807 2130 37816 2164
rect 37764 2121 37816 2130
rect 37764 2092 37816 2109
rect 37764 2058 37773 2092
rect 37773 2058 37807 2092
rect 37807 2058 37816 2092
rect 37764 2057 37816 2058
rect 37764 2020 37816 2045
rect 37764 1993 37773 2020
rect 37773 1993 37807 2020
rect 37807 1993 37816 2020
rect 37764 1948 37816 1981
rect 37764 1929 37773 1948
rect 37773 1929 37807 1948
rect 37807 1929 37816 1948
rect 37764 1914 37773 1917
rect 37773 1914 37807 1917
rect 37807 1914 37816 1917
rect 37764 1876 37816 1914
rect 37764 1865 37773 1876
rect 37773 1865 37807 1876
rect 37807 1865 37816 1876
rect 37764 1842 37773 1853
rect 37773 1842 37807 1853
rect 37807 1842 37816 1853
rect 37764 1804 37816 1842
rect 37764 1801 37773 1804
rect 37773 1801 37807 1804
rect 37807 1801 37816 1804
rect 37764 1770 37773 1789
rect 37773 1770 37807 1789
rect 37807 1770 37816 1789
rect 37764 1737 37816 1770
rect 37764 1698 37773 1725
rect 37773 1698 37807 1725
rect 37807 1698 37816 1725
rect 37764 1673 37816 1698
rect 37764 1660 37816 1661
rect 37764 1626 37773 1660
rect 37773 1626 37807 1660
rect 37807 1626 37816 1660
rect 37764 1609 37816 1626
rect 37764 1588 37816 1597
rect 37764 1554 37773 1588
rect 37773 1554 37807 1588
rect 37807 1554 37816 1588
rect 37764 1545 37816 1554
rect 37764 1516 37816 1533
rect 37764 1482 37773 1516
rect 37773 1482 37807 1516
rect 37807 1482 37816 1516
rect 37764 1481 37816 1482
rect 37764 1444 37816 1469
rect 37764 1417 37773 1444
rect 37773 1417 37807 1444
rect 37807 1417 37816 1444
rect 37764 1372 37816 1405
rect 37764 1353 37773 1372
rect 37773 1353 37807 1372
rect 37807 1353 37816 1372
rect 37764 1338 37773 1341
rect 37773 1338 37807 1341
rect 37807 1338 37816 1341
rect 37764 1300 37816 1338
rect 37764 1289 37773 1300
rect 37773 1289 37807 1300
rect 37807 1289 37816 1300
rect 37764 1266 37773 1277
rect 37773 1266 37807 1277
rect 37807 1266 37816 1277
rect 37764 1228 37816 1266
rect 37764 1225 37773 1228
rect 37773 1225 37807 1228
rect 37807 1225 37816 1228
rect 37764 1194 37773 1213
rect 37773 1194 37807 1213
rect 37807 1194 37816 1213
rect 37764 1161 37816 1194
rect 37860 3100 37912 3133
rect 37860 3081 37869 3100
rect 37869 3081 37903 3100
rect 37903 3081 37912 3100
rect 37860 3066 37869 3069
rect 37869 3066 37903 3069
rect 37903 3066 37912 3069
rect 37860 3028 37912 3066
rect 37860 3017 37869 3028
rect 37869 3017 37903 3028
rect 37903 3017 37912 3028
rect 37860 2994 37869 3005
rect 37869 2994 37903 3005
rect 37903 2994 37912 3005
rect 37860 2956 37912 2994
rect 37860 2953 37869 2956
rect 37869 2953 37903 2956
rect 37903 2953 37912 2956
rect 37860 2922 37869 2941
rect 37869 2922 37903 2941
rect 37903 2922 37912 2941
rect 37860 2889 37912 2922
rect 37860 2850 37869 2877
rect 37869 2850 37903 2877
rect 37903 2850 37912 2877
rect 37860 2825 37912 2850
rect 37860 2812 37912 2813
rect 37860 2778 37869 2812
rect 37869 2778 37903 2812
rect 37903 2778 37912 2812
rect 37860 2761 37912 2778
rect 37860 2740 37912 2749
rect 37860 2706 37869 2740
rect 37869 2706 37903 2740
rect 37903 2706 37912 2740
rect 37860 2697 37912 2706
rect 37860 2668 37912 2685
rect 37860 2634 37869 2668
rect 37869 2634 37903 2668
rect 37903 2634 37912 2668
rect 37860 2633 37912 2634
rect 37860 2596 37912 2621
rect 37860 2569 37869 2596
rect 37869 2569 37903 2596
rect 37903 2569 37912 2596
rect 37860 2524 37912 2557
rect 37860 2505 37869 2524
rect 37869 2505 37903 2524
rect 37903 2505 37912 2524
rect 37860 2490 37869 2493
rect 37869 2490 37903 2493
rect 37903 2490 37912 2493
rect 37860 2452 37912 2490
rect 37860 2441 37869 2452
rect 37869 2441 37903 2452
rect 37903 2441 37912 2452
rect 37860 2418 37869 2429
rect 37869 2418 37903 2429
rect 37903 2418 37912 2429
rect 37860 2380 37912 2418
rect 37860 2377 37869 2380
rect 37869 2377 37903 2380
rect 37903 2377 37912 2380
rect 37860 2346 37869 2365
rect 37869 2346 37903 2365
rect 37903 2346 37912 2365
rect 37860 2313 37912 2346
rect 37860 2274 37869 2301
rect 37869 2274 37903 2301
rect 37903 2274 37912 2301
rect 37860 2249 37912 2274
rect 37860 2236 37912 2237
rect 37860 2202 37869 2236
rect 37869 2202 37903 2236
rect 37903 2202 37912 2236
rect 37860 2185 37912 2202
rect 37860 2164 37912 2173
rect 37860 2130 37869 2164
rect 37869 2130 37903 2164
rect 37903 2130 37912 2164
rect 37860 2121 37912 2130
rect 37860 2092 37912 2109
rect 37860 2058 37869 2092
rect 37869 2058 37903 2092
rect 37903 2058 37912 2092
rect 37860 2057 37912 2058
rect 37860 2020 37912 2045
rect 37860 1993 37869 2020
rect 37869 1993 37903 2020
rect 37903 1993 37912 2020
rect 37860 1948 37912 1981
rect 37860 1929 37869 1948
rect 37869 1929 37903 1948
rect 37903 1929 37912 1948
rect 37860 1914 37869 1917
rect 37869 1914 37903 1917
rect 37903 1914 37912 1917
rect 37860 1876 37912 1914
rect 37860 1865 37869 1876
rect 37869 1865 37903 1876
rect 37903 1865 37912 1876
rect 37860 1842 37869 1853
rect 37869 1842 37903 1853
rect 37903 1842 37912 1853
rect 37860 1804 37912 1842
rect 37860 1801 37869 1804
rect 37869 1801 37903 1804
rect 37903 1801 37912 1804
rect 37860 1770 37869 1789
rect 37869 1770 37903 1789
rect 37903 1770 37912 1789
rect 37860 1737 37912 1770
rect 37860 1698 37869 1725
rect 37869 1698 37903 1725
rect 37903 1698 37912 1725
rect 37860 1673 37912 1698
rect 37860 1660 37912 1661
rect 37860 1626 37869 1660
rect 37869 1626 37903 1660
rect 37903 1626 37912 1660
rect 37860 1609 37912 1626
rect 37860 1588 37912 1597
rect 37860 1554 37869 1588
rect 37869 1554 37903 1588
rect 37903 1554 37912 1588
rect 37860 1545 37912 1554
rect 37860 1516 37912 1533
rect 37860 1482 37869 1516
rect 37869 1482 37903 1516
rect 37903 1482 37912 1516
rect 37860 1481 37912 1482
rect 37860 1444 37912 1469
rect 37860 1417 37869 1444
rect 37869 1417 37903 1444
rect 37903 1417 37912 1444
rect 37860 1372 37912 1405
rect 37860 1353 37869 1372
rect 37869 1353 37903 1372
rect 37903 1353 37912 1372
rect 37860 1338 37869 1341
rect 37869 1338 37903 1341
rect 37903 1338 37912 1341
rect 37860 1300 37912 1338
rect 37860 1289 37869 1300
rect 37869 1289 37903 1300
rect 37903 1289 37912 1300
rect 37860 1266 37869 1277
rect 37869 1266 37903 1277
rect 37903 1266 37912 1277
rect 37860 1228 37912 1266
rect 37860 1225 37869 1228
rect 37869 1225 37903 1228
rect 37903 1225 37912 1228
rect 37860 1194 37869 1213
rect 37869 1194 37903 1213
rect 37903 1194 37912 1213
rect 37860 1161 37912 1194
rect 37956 3100 38008 3133
rect 37956 3081 37965 3100
rect 37965 3081 37999 3100
rect 37999 3081 38008 3100
rect 37956 3066 37965 3069
rect 37965 3066 37999 3069
rect 37999 3066 38008 3069
rect 37956 3028 38008 3066
rect 37956 3017 37965 3028
rect 37965 3017 37999 3028
rect 37999 3017 38008 3028
rect 37956 2994 37965 3005
rect 37965 2994 37999 3005
rect 37999 2994 38008 3005
rect 37956 2956 38008 2994
rect 37956 2953 37965 2956
rect 37965 2953 37999 2956
rect 37999 2953 38008 2956
rect 37956 2922 37965 2941
rect 37965 2922 37999 2941
rect 37999 2922 38008 2941
rect 37956 2889 38008 2922
rect 37956 2850 37965 2877
rect 37965 2850 37999 2877
rect 37999 2850 38008 2877
rect 37956 2825 38008 2850
rect 37956 2812 38008 2813
rect 37956 2778 37965 2812
rect 37965 2778 37999 2812
rect 37999 2778 38008 2812
rect 37956 2761 38008 2778
rect 37956 2740 38008 2749
rect 37956 2706 37965 2740
rect 37965 2706 37999 2740
rect 37999 2706 38008 2740
rect 37956 2697 38008 2706
rect 37956 2668 38008 2685
rect 37956 2634 37965 2668
rect 37965 2634 37999 2668
rect 37999 2634 38008 2668
rect 37956 2633 38008 2634
rect 37956 2596 38008 2621
rect 37956 2569 37965 2596
rect 37965 2569 37999 2596
rect 37999 2569 38008 2596
rect 37956 2524 38008 2557
rect 37956 2505 37965 2524
rect 37965 2505 37999 2524
rect 37999 2505 38008 2524
rect 37956 2490 37965 2493
rect 37965 2490 37999 2493
rect 37999 2490 38008 2493
rect 37956 2452 38008 2490
rect 37956 2441 37965 2452
rect 37965 2441 37999 2452
rect 37999 2441 38008 2452
rect 37956 2418 37965 2429
rect 37965 2418 37999 2429
rect 37999 2418 38008 2429
rect 37956 2380 38008 2418
rect 37956 2377 37965 2380
rect 37965 2377 37999 2380
rect 37999 2377 38008 2380
rect 37956 2346 37965 2365
rect 37965 2346 37999 2365
rect 37999 2346 38008 2365
rect 37956 2313 38008 2346
rect 37956 2274 37965 2301
rect 37965 2274 37999 2301
rect 37999 2274 38008 2301
rect 37956 2249 38008 2274
rect 37956 2236 38008 2237
rect 37956 2202 37965 2236
rect 37965 2202 37999 2236
rect 37999 2202 38008 2236
rect 37956 2185 38008 2202
rect 37956 2164 38008 2173
rect 37956 2130 37965 2164
rect 37965 2130 37999 2164
rect 37999 2130 38008 2164
rect 37956 2121 38008 2130
rect 37956 2092 38008 2109
rect 37956 2058 37965 2092
rect 37965 2058 37999 2092
rect 37999 2058 38008 2092
rect 37956 2057 38008 2058
rect 37956 2020 38008 2045
rect 37956 1993 37965 2020
rect 37965 1993 37999 2020
rect 37999 1993 38008 2020
rect 37956 1948 38008 1981
rect 37956 1929 37965 1948
rect 37965 1929 37999 1948
rect 37999 1929 38008 1948
rect 37956 1914 37965 1917
rect 37965 1914 37999 1917
rect 37999 1914 38008 1917
rect 37956 1876 38008 1914
rect 37956 1865 37965 1876
rect 37965 1865 37999 1876
rect 37999 1865 38008 1876
rect 37956 1842 37965 1853
rect 37965 1842 37999 1853
rect 37999 1842 38008 1853
rect 37956 1804 38008 1842
rect 37956 1801 37965 1804
rect 37965 1801 37999 1804
rect 37999 1801 38008 1804
rect 37956 1770 37965 1789
rect 37965 1770 37999 1789
rect 37999 1770 38008 1789
rect 37956 1737 38008 1770
rect 37956 1698 37965 1725
rect 37965 1698 37999 1725
rect 37999 1698 38008 1725
rect 37956 1673 38008 1698
rect 37956 1660 38008 1661
rect 37956 1626 37965 1660
rect 37965 1626 37999 1660
rect 37999 1626 38008 1660
rect 37956 1609 38008 1626
rect 37956 1588 38008 1597
rect 37956 1554 37965 1588
rect 37965 1554 37999 1588
rect 37999 1554 38008 1588
rect 37956 1545 38008 1554
rect 37956 1516 38008 1533
rect 37956 1482 37965 1516
rect 37965 1482 37999 1516
rect 37999 1482 38008 1516
rect 37956 1481 38008 1482
rect 37956 1444 38008 1469
rect 37956 1417 37965 1444
rect 37965 1417 37999 1444
rect 37999 1417 38008 1444
rect 37956 1372 38008 1405
rect 37956 1353 37965 1372
rect 37965 1353 37999 1372
rect 37999 1353 38008 1372
rect 37956 1338 37965 1341
rect 37965 1338 37999 1341
rect 37999 1338 38008 1341
rect 37956 1300 38008 1338
rect 37956 1289 37965 1300
rect 37965 1289 37999 1300
rect 37999 1289 38008 1300
rect 37956 1266 37965 1277
rect 37965 1266 37999 1277
rect 37999 1266 38008 1277
rect 37956 1228 38008 1266
rect 37956 1225 37965 1228
rect 37965 1225 37999 1228
rect 37999 1225 38008 1228
rect 37956 1194 37965 1213
rect 37965 1194 37999 1213
rect 37999 1194 38008 1213
rect 37956 1161 38008 1194
rect 38052 3100 38104 3133
rect 38052 3081 38061 3100
rect 38061 3081 38095 3100
rect 38095 3081 38104 3100
rect 38052 3066 38061 3069
rect 38061 3066 38095 3069
rect 38095 3066 38104 3069
rect 38052 3028 38104 3066
rect 38052 3017 38061 3028
rect 38061 3017 38095 3028
rect 38095 3017 38104 3028
rect 38052 2994 38061 3005
rect 38061 2994 38095 3005
rect 38095 2994 38104 3005
rect 38052 2956 38104 2994
rect 38052 2953 38061 2956
rect 38061 2953 38095 2956
rect 38095 2953 38104 2956
rect 38052 2922 38061 2941
rect 38061 2922 38095 2941
rect 38095 2922 38104 2941
rect 38052 2889 38104 2922
rect 38052 2850 38061 2877
rect 38061 2850 38095 2877
rect 38095 2850 38104 2877
rect 38052 2825 38104 2850
rect 38052 2812 38104 2813
rect 38052 2778 38061 2812
rect 38061 2778 38095 2812
rect 38095 2778 38104 2812
rect 38052 2761 38104 2778
rect 38052 2740 38104 2749
rect 38052 2706 38061 2740
rect 38061 2706 38095 2740
rect 38095 2706 38104 2740
rect 38052 2697 38104 2706
rect 38052 2668 38104 2685
rect 38052 2634 38061 2668
rect 38061 2634 38095 2668
rect 38095 2634 38104 2668
rect 38052 2633 38104 2634
rect 38052 2596 38104 2621
rect 38052 2569 38061 2596
rect 38061 2569 38095 2596
rect 38095 2569 38104 2596
rect 38052 2524 38104 2557
rect 38052 2505 38061 2524
rect 38061 2505 38095 2524
rect 38095 2505 38104 2524
rect 38052 2490 38061 2493
rect 38061 2490 38095 2493
rect 38095 2490 38104 2493
rect 38052 2452 38104 2490
rect 38052 2441 38061 2452
rect 38061 2441 38095 2452
rect 38095 2441 38104 2452
rect 38052 2418 38061 2429
rect 38061 2418 38095 2429
rect 38095 2418 38104 2429
rect 38052 2380 38104 2418
rect 38052 2377 38061 2380
rect 38061 2377 38095 2380
rect 38095 2377 38104 2380
rect 38052 2346 38061 2365
rect 38061 2346 38095 2365
rect 38095 2346 38104 2365
rect 38052 2313 38104 2346
rect 38052 2274 38061 2301
rect 38061 2274 38095 2301
rect 38095 2274 38104 2301
rect 38052 2249 38104 2274
rect 38052 2236 38104 2237
rect 38052 2202 38061 2236
rect 38061 2202 38095 2236
rect 38095 2202 38104 2236
rect 38052 2185 38104 2202
rect 38052 2164 38104 2173
rect 38052 2130 38061 2164
rect 38061 2130 38095 2164
rect 38095 2130 38104 2164
rect 38052 2121 38104 2130
rect 38052 2092 38104 2109
rect 38052 2058 38061 2092
rect 38061 2058 38095 2092
rect 38095 2058 38104 2092
rect 38052 2057 38104 2058
rect 38052 2020 38104 2045
rect 38052 1993 38061 2020
rect 38061 1993 38095 2020
rect 38095 1993 38104 2020
rect 38052 1948 38104 1981
rect 38052 1929 38061 1948
rect 38061 1929 38095 1948
rect 38095 1929 38104 1948
rect 38052 1914 38061 1917
rect 38061 1914 38095 1917
rect 38095 1914 38104 1917
rect 38052 1876 38104 1914
rect 38052 1865 38061 1876
rect 38061 1865 38095 1876
rect 38095 1865 38104 1876
rect 38052 1842 38061 1853
rect 38061 1842 38095 1853
rect 38095 1842 38104 1853
rect 38052 1804 38104 1842
rect 38052 1801 38061 1804
rect 38061 1801 38095 1804
rect 38095 1801 38104 1804
rect 38052 1770 38061 1789
rect 38061 1770 38095 1789
rect 38095 1770 38104 1789
rect 38052 1737 38104 1770
rect 38052 1698 38061 1725
rect 38061 1698 38095 1725
rect 38095 1698 38104 1725
rect 38052 1673 38104 1698
rect 38052 1660 38104 1661
rect 38052 1626 38061 1660
rect 38061 1626 38095 1660
rect 38095 1626 38104 1660
rect 38052 1609 38104 1626
rect 38052 1588 38104 1597
rect 38052 1554 38061 1588
rect 38061 1554 38095 1588
rect 38095 1554 38104 1588
rect 38052 1545 38104 1554
rect 38052 1516 38104 1533
rect 38052 1482 38061 1516
rect 38061 1482 38095 1516
rect 38095 1482 38104 1516
rect 38052 1481 38104 1482
rect 38052 1444 38104 1469
rect 38052 1417 38061 1444
rect 38061 1417 38095 1444
rect 38095 1417 38104 1444
rect 38052 1372 38104 1405
rect 38052 1353 38061 1372
rect 38061 1353 38095 1372
rect 38095 1353 38104 1372
rect 38052 1338 38061 1341
rect 38061 1338 38095 1341
rect 38095 1338 38104 1341
rect 38052 1300 38104 1338
rect 38052 1289 38061 1300
rect 38061 1289 38095 1300
rect 38095 1289 38104 1300
rect 38052 1266 38061 1277
rect 38061 1266 38095 1277
rect 38095 1266 38104 1277
rect 38052 1228 38104 1266
rect 38052 1225 38061 1228
rect 38061 1225 38095 1228
rect 38095 1225 38104 1228
rect 38052 1194 38061 1213
rect 38061 1194 38095 1213
rect 38095 1194 38104 1213
rect 38052 1161 38104 1194
rect 38148 3100 38200 3133
rect 38148 3081 38157 3100
rect 38157 3081 38191 3100
rect 38191 3081 38200 3100
rect 38148 3066 38157 3069
rect 38157 3066 38191 3069
rect 38191 3066 38200 3069
rect 38148 3028 38200 3066
rect 38148 3017 38157 3028
rect 38157 3017 38191 3028
rect 38191 3017 38200 3028
rect 38148 2994 38157 3005
rect 38157 2994 38191 3005
rect 38191 2994 38200 3005
rect 38148 2956 38200 2994
rect 38148 2953 38157 2956
rect 38157 2953 38191 2956
rect 38191 2953 38200 2956
rect 38148 2922 38157 2941
rect 38157 2922 38191 2941
rect 38191 2922 38200 2941
rect 38148 2889 38200 2922
rect 38148 2850 38157 2877
rect 38157 2850 38191 2877
rect 38191 2850 38200 2877
rect 38148 2825 38200 2850
rect 38148 2812 38200 2813
rect 38148 2778 38157 2812
rect 38157 2778 38191 2812
rect 38191 2778 38200 2812
rect 38148 2761 38200 2778
rect 38148 2740 38200 2749
rect 38148 2706 38157 2740
rect 38157 2706 38191 2740
rect 38191 2706 38200 2740
rect 38148 2697 38200 2706
rect 38148 2668 38200 2685
rect 38148 2634 38157 2668
rect 38157 2634 38191 2668
rect 38191 2634 38200 2668
rect 38148 2633 38200 2634
rect 38148 2596 38200 2621
rect 38148 2569 38157 2596
rect 38157 2569 38191 2596
rect 38191 2569 38200 2596
rect 38148 2524 38200 2557
rect 38148 2505 38157 2524
rect 38157 2505 38191 2524
rect 38191 2505 38200 2524
rect 38148 2490 38157 2493
rect 38157 2490 38191 2493
rect 38191 2490 38200 2493
rect 38148 2452 38200 2490
rect 38148 2441 38157 2452
rect 38157 2441 38191 2452
rect 38191 2441 38200 2452
rect 38148 2418 38157 2429
rect 38157 2418 38191 2429
rect 38191 2418 38200 2429
rect 38148 2380 38200 2418
rect 38148 2377 38157 2380
rect 38157 2377 38191 2380
rect 38191 2377 38200 2380
rect 38148 2346 38157 2365
rect 38157 2346 38191 2365
rect 38191 2346 38200 2365
rect 38148 2313 38200 2346
rect 38148 2274 38157 2301
rect 38157 2274 38191 2301
rect 38191 2274 38200 2301
rect 38148 2249 38200 2274
rect 38148 2236 38200 2237
rect 38148 2202 38157 2236
rect 38157 2202 38191 2236
rect 38191 2202 38200 2236
rect 38148 2185 38200 2202
rect 38148 2164 38200 2173
rect 38148 2130 38157 2164
rect 38157 2130 38191 2164
rect 38191 2130 38200 2164
rect 38148 2121 38200 2130
rect 38148 2092 38200 2109
rect 38148 2058 38157 2092
rect 38157 2058 38191 2092
rect 38191 2058 38200 2092
rect 38148 2057 38200 2058
rect 38148 2020 38200 2045
rect 38148 1993 38157 2020
rect 38157 1993 38191 2020
rect 38191 1993 38200 2020
rect 38148 1948 38200 1981
rect 38148 1929 38157 1948
rect 38157 1929 38191 1948
rect 38191 1929 38200 1948
rect 38148 1914 38157 1917
rect 38157 1914 38191 1917
rect 38191 1914 38200 1917
rect 38148 1876 38200 1914
rect 38148 1865 38157 1876
rect 38157 1865 38191 1876
rect 38191 1865 38200 1876
rect 38148 1842 38157 1853
rect 38157 1842 38191 1853
rect 38191 1842 38200 1853
rect 38148 1804 38200 1842
rect 38148 1801 38157 1804
rect 38157 1801 38191 1804
rect 38191 1801 38200 1804
rect 38148 1770 38157 1789
rect 38157 1770 38191 1789
rect 38191 1770 38200 1789
rect 38148 1737 38200 1770
rect 38148 1698 38157 1725
rect 38157 1698 38191 1725
rect 38191 1698 38200 1725
rect 38148 1673 38200 1698
rect 38148 1660 38200 1661
rect 38148 1626 38157 1660
rect 38157 1626 38191 1660
rect 38191 1626 38200 1660
rect 38148 1609 38200 1626
rect 38148 1588 38200 1597
rect 38148 1554 38157 1588
rect 38157 1554 38191 1588
rect 38191 1554 38200 1588
rect 38148 1545 38200 1554
rect 38148 1516 38200 1533
rect 38148 1482 38157 1516
rect 38157 1482 38191 1516
rect 38191 1482 38200 1516
rect 38148 1481 38200 1482
rect 38148 1444 38200 1469
rect 38148 1417 38157 1444
rect 38157 1417 38191 1444
rect 38191 1417 38200 1444
rect 38148 1372 38200 1405
rect 38148 1353 38157 1372
rect 38157 1353 38191 1372
rect 38191 1353 38200 1372
rect 38148 1338 38157 1341
rect 38157 1338 38191 1341
rect 38191 1338 38200 1341
rect 38148 1300 38200 1338
rect 38148 1289 38157 1300
rect 38157 1289 38191 1300
rect 38191 1289 38200 1300
rect 38148 1266 38157 1277
rect 38157 1266 38191 1277
rect 38191 1266 38200 1277
rect 38148 1228 38200 1266
rect 38148 1225 38157 1228
rect 38157 1225 38191 1228
rect 38191 1225 38200 1228
rect 38148 1194 38157 1213
rect 38157 1194 38191 1213
rect 38191 1194 38200 1213
rect 38148 1161 38200 1194
rect 38244 3100 38296 3133
rect 38244 3081 38253 3100
rect 38253 3081 38287 3100
rect 38287 3081 38296 3100
rect 38244 3066 38253 3069
rect 38253 3066 38287 3069
rect 38287 3066 38296 3069
rect 38244 3028 38296 3066
rect 38244 3017 38253 3028
rect 38253 3017 38287 3028
rect 38287 3017 38296 3028
rect 38244 2994 38253 3005
rect 38253 2994 38287 3005
rect 38287 2994 38296 3005
rect 38244 2956 38296 2994
rect 38244 2953 38253 2956
rect 38253 2953 38287 2956
rect 38287 2953 38296 2956
rect 38244 2922 38253 2941
rect 38253 2922 38287 2941
rect 38287 2922 38296 2941
rect 38244 2889 38296 2922
rect 38244 2850 38253 2877
rect 38253 2850 38287 2877
rect 38287 2850 38296 2877
rect 38244 2825 38296 2850
rect 38244 2812 38296 2813
rect 38244 2778 38253 2812
rect 38253 2778 38287 2812
rect 38287 2778 38296 2812
rect 38244 2761 38296 2778
rect 38244 2740 38296 2749
rect 38244 2706 38253 2740
rect 38253 2706 38287 2740
rect 38287 2706 38296 2740
rect 38244 2697 38296 2706
rect 38244 2668 38296 2685
rect 38244 2634 38253 2668
rect 38253 2634 38287 2668
rect 38287 2634 38296 2668
rect 38244 2633 38296 2634
rect 38244 2596 38296 2621
rect 38244 2569 38253 2596
rect 38253 2569 38287 2596
rect 38287 2569 38296 2596
rect 38244 2524 38296 2557
rect 38244 2505 38253 2524
rect 38253 2505 38287 2524
rect 38287 2505 38296 2524
rect 38244 2490 38253 2493
rect 38253 2490 38287 2493
rect 38287 2490 38296 2493
rect 38244 2452 38296 2490
rect 38244 2441 38253 2452
rect 38253 2441 38287 2452
rect 38287 2441 38296 2452
rect 38244 2418 38253 2429
rect 38253 2418 38287 2429
rect 38287 2418 38296 2429
rect 38244 2380 38296 2418
rect 38244 2377 38253 2380
rect 38253 2377 38287 2380
rect 38287 2377 38296 2380
rect 38244 2346 38253 2365
rect 38253 2346 38287 2365
rect 38287 2346 38296 2365
rect 38244 2313 38296 2346
rect 38244 2274 38253 2301
rect 38253 2274 38287 2301
rect 38287 2274 38296 2301
rect 38244 2249 38296 2274
rect 38244 2236 38296 2237
rect 38244 2202 38253 2236
rect 38253 2202 38287 2236
rect 38287 2202 38296 2236
rect 38244 2185 38296 2202
rect 38244 2164 38296 2173
rect 38244 2130 38253 2164
rect 38253 2130 38287 2164
rect 38287 2130 38296 2164
rect 38244 2121 38296 2130
rect 38244 2092 38296 2109
rect 38244 2058 38253 2092
rect 38253 2058 38287 2092
rect 38287 2058 38296 2092
rect 38244 2057 38296 2058
rect 38244 2020 38296 2045
rect 38244 1993 38253 2020
rect 38253 1993 38287 2020
rect 38287 1993 38296 2020
rect 38244 1948 38296 1981
rect 38244 1929 38253 1948
rect 38253 1929 38287 1948
rect 38287 1929 38296 1948
rect 38244 1914 38253 1917
rect 38253 1914 38287 1917
rect 38287 1914 38296 1917
rect 38244 1876 38296 1914
rect 38244 1865 38253 1876
rect 38253 1865 38287 1876
rect 38287 1865 38296 1876
rect 38244 1842 38253 1853
rect 38253 1842 38287 1853
rect 38287 1842 38296 1853
rect 38244 1804 38296 1842
rect 38244 1801 38253 1804
rect 38253 1801 38287 1804
rect 38287 1801 38296 1804
rect 38244 1770 38253 1789
rect 38253 1770 38287 1789
rect 38287 1770 38296 1789
rect 38244 1737 38296 1770
rect 38244 1698 38253 1725
rect 38253 1698 38287 1725
rect 38287 1698 38296 1725
rect 38244 1673 38296 1698
rect 38244 1660 38296 1661
rect 38244 1626 38253 1660
rect 38253 1626 38287 1660
rect 38287 1626 38296 1660
rect 38244 1609 38296 1626
rect 38244 1588 38296 1597
rect 38244 1554 38253 1588
rect 38253 1554 38287 1588
rect 38287 1554 38296 1588
rect 38244 1545 38296 1554
rect 38244 1516 38296 1533
rect 38244 1482 38253 1516
rect 38253 1482 38287 1516
rect 38287 1482 38296 1516
rect 38244 1481 38296 1482
rect 38244 1444 38296 1469
rect 38244 1417 38253 1444
rect 38253 1417 38287 1444
rect 38287 1417 38296 1444
rect 38244 1372 38296 1405
rect 38244 1353 38253 1372
rect 38253 1353 38287 1372
rect 38287 1353 38296 1372
rect 38244 1338 38253 1341
rect 38253 1338 38287 1341
rect 38287 1338 38296 1341
rect 38244 1300 38296 1338
rect 38244 1289 38253 1300
rect 38253 1289 38287 1300
rect 38287 1289 38296 1300
rect 38244 1266 38253 1277
rect 38253 1266 38287 1277
rect 38287 1266 38296 1277
rect 38244 1228 38296 1266
rect 38244 1225 38253 1228
rect 38253 1225 38287 1228
rect 38287 1225 38296 1228
rect 38244 1194 38253 1213
rect 38253 1194 38287 1213
rect 38287 1194 38296 1213
rect 38244 1161 38296 1194
rect 38340 3100 38392 3133
rect 38340 3081 38349 3100
rect 38349 3081 38383 3100
rect 38383 3081 38392 3100
rect 38340 3066 38349 3069
rect 38349 3066 38383 3069
rect 38383 3066 38392 3069
rect 38340 3028 38392 3066
rect 38340 3017 38349 3028
rect 38349 3017 38383 3028
rect 38383 3017 38392 3028
rect 38340 2994 38349 3005
rect 38349 2994 38383 3005
rect 38383 2994 38392 3005
rect 38340 2956 38392 2994
rect 38340 2953 38349 2956
rect 38349 2953 38383 2956
rect 38383 2953 38392 2956
rect 38340 2922 38349 2941
rect 38349 2922 38383 2941
rect 38383 2922 38392 2941
rect 38340 2889 38392 2922
rect 38340 2850 38349 2877
rect 38349 2850 38383 2877
rect 38383 2850 38392 2877
rect 38340 2825 38392 2850
rect 38340 2812 38392 2813
rect 38340 2778 38349 2812
rect 38349 2778 38383 2812
rect 38383 2778 38392 2812
rect 38340 2761 38392 2778
rect 38340 2740 38392 2749
rect 38340 2706 38349 2740
rect 38349 2706 38383 2740
rect 38383 2706 38392 2740
rect 38340 2697 38392 2706
rect 38340 2668 38392 2685
rect 38340 2634 38349 2668
rect 38349 2634 38383 2668
rect 38383 2634 38392 2668
rect 38340 2633 38392 2634
rect 38340 2596 38392 2621
rect 38340 2569 38349 2596
rect 38349 2569 38383 2596
rect 38383 2569 38392 2596
rect 38340 2524 38392 2557
rect 38340 2505 38349 2524
rect 38349 2505 38383 2524
rect 38383 2505 38392 2524
rect 38340 2490 38349 2493
rect 38349 2490 38383 2493
rect 38383 2490 38392 2493
rect 38340 2452 38392 2490
rect 38340 2441 38349 2452
rect 38349 2441 38383 2452
rect 38383 2441 38392 2452
rect 38340 2418 38349 2429
rect 38349 2418 38383 2429
rect 38383 2418 38392 2429
rect 38340 2380 38392 2418
rect 38340 2377 38349 2380
rect 38349 2377 38383 2380
rect 38383 2377 38392 2380
rect 38340 2346 38349 2365
rect 38349 2346 38383 2365
rect 38383 2346 38392 2365
rect 38340 2313 38392 2346
rect 38340 2274 38349 2301
rect 38349 2274 38383 2301
rect 38383 2274 38392 2301
rect 38340 2249 38392 2274
rect 38340 2236 38392 2237
rect 38340 2202 38349 2236
rect 38349 2202 38383 2236
rect 38383 2202 38392 2236
rect 38340 2185 38392 2202
rect 38340 2164 38392 2173
rect 38340 2130 38349 2164
rect 38349 2130 38383 2164
rect 38383 2130 38392 2164
rect 38340 2121 38392 2130
rect 38340 2092 38392 2109
rect 38340 2058 38349 2092
rect 38349 2058 38383 2092
rect 38383 2058 38392 2092
rect 38340 2057 38392 2058
rect 38340 2020 38392 2045
rect 38340 1993 38349 2020
rect 38349 1993 38383 2020
rect 38383 1993 38392 2020
rect 38340 1948 38392 1981
rect 38340 1929 38349 1948
rect 38349 1929 38383 1948
rect 38383 1929 38392 1948
rect 38340 1914 38349 1917
rect 38349 1914 38383 1917
rect 38383 1914 38392 1917
rect 38340 1876 38392 1914
rect 38340 1865 38349 1876
rect 38349 1865 38383 1876
rect 38383 1865 38392 1876
rect 38340 1842 38349 1853
rect 38349 1842 38383 1853
rect 38383 1842 38392 1853
rect 38340 1804 38392 1842
rect 38340 1801 38349 1804
rect 38349 1801 38383 1804
rect 38383 1801 38392 1804
rect 38340 1770 38349 1789
rect 38349 1770 38383 1789
rect 38383 1770 38392 1789
rect 38340 1737 38392 1770
rect 38340 1698 38349 1725
rect 38349 1698 38383 1725
rect 38383 1698 38392 1725
rect 38340 1673 38392 1698
rect 38340 1660 38392 1661
rect 38340 1626 38349 1660
rect 38349 1626 38383 1660
rect 38383 1626 38392 1660
rect 38340 1609 38392 1626
rect 38340 1588 38392 1597
rect 38340 1554 38349 1588
rect 38349 1554 38383 1588
rect 38383 1554 38392 1588
rect 38340 1545 38392 1554
rect 38340 1516 38392 1533
rect 38340 1482 38349 1516
rect 38349 1482 38383 1516
rect 38383 1482 38392 1516
rect 38340 1481 38392 1482
rect 38340 1444 38392 1469
rect 38340 1417 38349 1444
rect 38349 1417 38383 1444
rect 38383 1417 38392 1444
rect 38340 1372 38392 1405
rect 38340 1353 38349 1372
rect 38349 1353 38383 1372
rect 38383 1353 38392 1372
rect 38340 1338 38349 1341
rect 38349 1338 38383 1341
rect 38383 1338 38392 1341
rect 38340 1300 38392 1338
rect 38340 1289 38349 1300
rect 38349 1289 38383 1300
rect 38383 1289 38392 1300
rect 38340 1266 38349 1277
rect 38349 1266 38383 1277
rect 38383 1266 38392 1277
rect 38340 1228 38392 1266
rect 38340 1225 38349 1228
rect 38349 1225 38383 1228
rect 38383 1225 38392 1228
rect 38340 1194 38349 1213
rect 38349 1194 38383 1213
rect 38383 1194 38392 1213
rect 38340 1161 38392 1194
rect 38436 3100 38488 3133
rect 38436 3081 38445 3100
rect 38445 3081 38479 3100
rect 38479 3081 38488 3100
rect 38436 3066 38445 3069
rect 38445 3066 38479 3069
rect 38479 3066 38488 3069
rect 38436 3028 38488 3066
rect 38436 3017 38445 3028
rect 38445 3017 38479 3028
rect 38479 3017 38488 3028
rect 38436 2994 38445 3005
rect 38445 2994 38479 3005
rect 38479 2994 38488 3005
rect 38436 2956 38488 2994
rect 38436 2953 38445 2956
rect 38445 2953 38479 2956
rect 38479 2953 38488 2956
rect 38436 2922 38445 2941
rect 38445 2922 38479 2941
rect 38479 2922 38488 2941
rect 38436 2889 38488 2922
rect 38436 2850 38445 2877
rect 38445 2850 38479 2877
rect 38479 2850 38488 2877
rect 38436 2825 38488 2850
rect 38436 2812 38488 2813
rect 38436 2778 38445 2812
rect 38445 2778 38479 2812
rect 38479 2778 38488 2812
rect 38436 2761 38488 2778
rect 38436 2740 38488 2749
rect 38436 2706 38445 2740
rect 38445 2706 38479 2740
rect 38479 2706 38488 2740
rect 38436 2697 38488 2706
rect 38436 2668 38488 2685
rect 38436 2634 38445 2668
rect 38445 2634 38479 2668
rect 38479 2634 38488 2668
rect 38436 2633 38488 2634
rect 38436 2596 38488 2621
rect 38436 2569 38445 2596
rect 38445 2569 38479 2596
rect 38479 2569 38488 2596
rect 38436 2524 38488 2557
rect 38436 2505 38445 2524
rect 38445 2505 38479 2524
rect 38479 2505 38488 2524
rect 38436 2490 38445 2493
rect 38445 2490 38479 2493
rect 38479 2490 38488 2493
rect 38436 2452 38488 2490
rect 38436 2441 38445 2452
rect 38445 2441 38479 2452
rect 38479 2441 38488 2452
rect 38436 2418 38445 2429
rect 38445 2418 38479 2429
rect 38479 2418 38488 2429
rect 38436 2380 38488 2418
rect 38436 2377 38445 2380
rect 38445 2377 38479 2380
rect 38479 2377 38488 2380
rect 38436 2346 38445 2365
rect 38445 2346 38479 2365
rect 38479 2346 38488 2365
rect 38436 2313 38488 2346
rect 38436 2274 38445 2301
rect 38445 2274 38479 2301
rect 38479 2274 38488 2301
rect 38436 2249 38488 2274
rect 38436 2236 38488 2237
rect 38436 2202 38445 2236
rect 38445 2202 38479 2236
rect 38479 2202 38488 2236
rect 38436 2185 38488 2202
rect 38436 2164 38488 2173
rect 38436 2130 38445 2164
rect 38445 2130 38479 2164
rect 38479 2130 38488 2164
rect 38436 2121 38488 2130
rect 38436 2092 38488 2109
rect 38436 2058 38445 2092
rect 38445 2058 38479 2092
rect 38479 2058 38488 2092
rect 38436 2057 38488 2058
rect 38436 2020 38488 2045
rect 38436 1993 38445 2020
rect 38445 1993 38479 2020
rect 38479 1993 38488 2020
rect 38436 1948 38488 1981
rect 38436 1929 38445 1948
rect 38445 1929 38479 1948
rect 38479 1929 38488 1948
rect 38436 1914 38445 1917
rect 38445 1914 38479 1917
rect 38479 1914 38488 1917
rect 38436 1876 38488 1914
rect 38436 1865 38445 1876
rect 38445 1865 38479 1876
rect 38479 1865 38488 1876
rect 38436 1842 38445 1853
rect 38445 1842 38479 1853
rect 38479 1842 38488 1853
rect 38436 1804 38488 1842
rect 38436 1801 38445 1804
rect 38445 1801 38479 1804
rect 38479 1801 38488 1804
rect 38436 1770 38445 1789
rect 38445 1770 38479 1789
rect 38479 1770 38488 1789
rect 38436 1737 38488 1770
rect 38436 1698 38445 1725
rect 38445 1698 38479 1725
rect 38479 1698 38488 1725
rect 38436 1673 38488 1698
rect 38436 1660 38488 1661
rect 38436 1626 38445 1660
rect 38445 1626 38479 1660
rect 38479 1626 38488 1660
rect 38436 1609 38488 1626
rect 38436 1588 38488 1597
rect 38436 1554 38445 1588
rect 38445 1554 38479 1588
rect 38479 1554 38488 1588
rect 38436 1545 38488 1554
rect 38436 1516 38488 1533
rect 38436 1482 38445 1516
rect 38445 1482 38479 1516
rect 38479 1482 38488 1516
rect 38436 1481 38488 1482
rect 38436 1444 38488 1469
rect 38436 1417 38445 1444
rect 38445 1417 38479 1444
rect 38479 1417 38488 1444
rect 38436 1372 38488 1405
rect 38436 1353 38445 1372
rect 38445 1353 38479 1372
rect 38479 1353 38488 1372
rect 38436 1338 38445 1341
rect 38445 1338 38479 1341
rect 38479 1338 38488 1341
rect 38436 1300 38488 1338
rect 38436 1289 38445 1300
rect 38445 1289 38479 1300
rect 38479 1289 38488 1300
rect 38436 1266 38445 1277
rect 38445 1266 38479 1277
rect 38479 1266 38488 1277
rect 38436 1228 38488 1266
rect 38436 1225 38445 1228
rect 38445 1225 38479 1228
rect 38479 1225 38488 1228
rect 38436 1194 38445 1213
rect 38445 1194 38479 1213
rect 38479 1194 38488 1213
rect 38436 1161 38488 1194
rect 38532 3100 38584 3133
rect 38532 3081 38541 3100
rect 38541 3081 38575 3100
rect 38575 3081 38584 3100
rect 38532 3066 38541 3069
rect 38541 3066 38575 3069
rect 38575 3066 38584 3069
rect 38532 3028 38584 3066
rect 38532 3017 38541 3028
rect 38541 3017 38575 3028
rect 38575 3017 38584 3028
rect 38532 2994 38541 3005
rect 38541 2994 38575 3005
rect 38575 2994 38584 3005
rect 38532 2956 38584 2994
rect 38532 2953 38541 2956
rect 38541 2953 38575 2956
rect 38575 2953 38584 2956
rect 38532 2922 38541 2941
rect 38541 2922 38575 2941
rect 38575 2922 38584 2941
rect 38532 2889 38584 2922
rect 38532 2850 38541 2877
rect 38541 2850 38575 2877
rect 38575 2850 38584 2877
rect 38532 2825 38584 2850
rect 38532 2812 38584 2813
rect 38532 2778 38541 2812
rect 38541 2778 38575 2812
rect 38575 2778 38584 2812
rect 38532 2761 38584 2778
rect 38532 2740 38584 2749
rect 38532 2706 38541 2740
rect 38541 2706 38575 2740
rect 38575 2706 38584 2740
rect 38532 2697 38584 2706
rect 38532 2668 38584 2685
rect 38532 2634 38541 2668
rect 38541 2634 38575 2668
rect 38575 2634 38584 2668
rect 38532 2633 38584 2634
rect 38532 2596 38584 2621
rect 38532 2569 38541 2596
rect 38541 2569 38575 2596
rect 38575 2569 38584 2596
rect 38532 2524 38584 2557
rect 38532 2505 38541 2524
rect 38541 2505 38575 2524
rect 38575 2505 38584 2524
rect 38532 2490 38541 2493
rect 38541 2490 38575 2493
rect 38575 2490 38584 2493
rect 38532 2452 38584 2490
rect 38532 2441 38541 2452
rect 38541 2441 38575 2452
rect 38575 2441 38584 2452
rect 38532 2418 38541 2429
rect 38541 2418 38575 2429
rect 38575 2418 38584 2429
rect 38532 2380 38584 2418
rect 38532 2377 38541 2380
rect 38541 2377 38575 2380
rect 38575 2377 38584 2380
rect 38532 2346 38541 2365
rect 38541 2346 38575 2365
rect 38575 2346 38584 2365
rect 38532 2313 38584 2346
rect 38532 2274 38541 2301
rect 38541 2274 38575 2301
rect 38575 2274 38584 2301
rect 38532 2249 38584 2274
rect 38532 2236 38584 2237
rect 38532 2202 38541 2236
rect 38541 2202 38575 2236
rect 38575 2202 38584 2236
rect 38532 2185 38584 2202
rect 38532 2164 38584 2173
rect 38532 2130 38541 2164
rect 38541 2130 38575 2164
rect 38575 2130 38584 2164
rect 38532 2121 38584 2130
rect 38532 2092 38584 2109
rect 38532 2058 38541 2092
rect 38541 2058 38575 2092
rect 38575 2058 38584 2092
rect 38532 2057 38584 2058
rect 38532 2020 38584 2045
rect 38532 1993 38541 2020
rect 38541 1993 38575 2020
rect 38575 1993 38584 2020
rect 38532 1948 38584 1981
rect 38532 1929 38541 1948
rect 38541 1929 38575 1948
rect 38575 1929 38584 1948
rect 38532 1914 38541 1917
rect 38541 1914 38575 1917
rect 38575 1914 38584 1917
rect 38532 1876 38584 1914
rect 38532 1865 38541 1876
rect 38541 1865 38575 1876
rect 38575 1865 38584 1876
rect 38532 1842 38541 1853
rect 38541 1842 38575 1853
rect 38575 1842 38584 1853
rect 38532 1804 38584 1842
rect 38532 1801 38541 1804
rect 38541 1801 38575 1804
rect 38575 1801 38584 1804
rect 38532 1770 38541 1789
rect 38541 1770 38575 1789
rect 38575 1770 38584 1789
rect 38532 1737 38584 1770
rect 38532 1698 38541 1725
rect 38541 1698 38575 1725
rect 38575 1698 38584 1725
rect 38532 1673 38584 1698
rect 38532 1660 38584 1661
rect 38532 1626 38541 1660
rect 38541 1626 38575 1660
rect 38575 1626 38584 1660
rect 38532 1609 38584 1626
rect 38532 1588 38584 1597
rect 38532 1554 38541 1588
rect 38541 1554 38575 1588
rect 38575 1554 38584 1588
rect 38532 1545 38584 1554
rect 38532 1516 38584 1533
rect 38532 1482 38541 1516
rect 38541 1482 38575 1516
rect 38575 1482 38584 1516
rect 38532 1481 38584 1482
rect 38532 1444 38584 1469
rect 38532 1417 38541 1444
rect 38541 1417 38575 1444
rect 38575 1417 38584 1444
rect 38532 1372 38584 1405
rect 38532 1353 38541 1372
rect 38541 1353 38575 1372
rect 38575 1353 38584 1372
rect 38532 1338 38541 1341
rect 38541 1338 38575 1341
rect 38575 1338 38584 1341
rect 38532 1300 38584 1338
rect 38532 1289 38541 1300
rect 38541 1289 38575 1300
rect 38575 1289 38584 1300
rect 38532 1266 38541 1277
rect 38541 1266 38575 1277
rect 38575 1266 38584 1277
rect 38532 1228 38584 1266
rect 38532 1225 38541 1228
rect 38541 1225 38575 1228
rect 38575 1225 38584 1228
rect 38532 1194 38541 1213
rect 38541 1194 38575 1213
rect 38575 1194 38584 1213
rect 38532 1161 38584 1194
rect 38628 3099 38680 3132
rect 38628 3080 38637 3099
rect 38637 3080 38671 3099
rect 38671 3080 38680 3099
rect 38628 3065 38637 3068
rect 38637 3065 38671 3068
rect 38671 3065 38680 3068
rect 38628 3027 38680 3065
rect 38628 3016 38637 3027
rect 38637 3016 38671 3027
rect 38671 3016 38680 3027
rect 38628 2993 38637 3004
rect 38637 2993 38671 3004
rect 38671 2993 38680 3004
rect 38628 2955 38680 2993
rect 38628 2952 38637 2955
rect 38637 2952 38671 2955
rect 38671 2952 38680 2955
rect 38628 2921 38637 2940
rect 38637 2921 38671 2940
rect 38671 2921 38680 2940
rect 38628 2888 38680 2921
rect 38628 2849 38637 2876
rect 38637 2849 38671 2876
rect 38671 2849 38680 2876
rect 38628 2824 38680 2849
rect 38628 2811 38680 2812
rect 38628 2777 38637 2811
rect 38637 2777 38671 2811
rect 38671 2777 38680 2811
rect 38628 2760 38680 2777
rect 38628 2739 38680 2748
rect 38628 2705 38637 2739
rect 38637 2705 38671 2739
rect 38671 2705 38680 2739
rect 38628 2696 38680 2705
rect 38628 2667 38680 2684
rect 38628 2633 38637 2667
rect 38637 2633 38671 2667
rect 38671 2633 38680 2667
rect 38628 2632 38680 2633
rect 38628 2595 38680 2620
rect 38628 2568 38637 2595
rect 38637 2568 38671 2595
rect 38671 2568 38680 2595
rect 38628 2523 38680 2556
rect 38628 2504 38637 2523
rect 38637 2504 38671 2523
rect 38671 2504 38680 2523
rect 38628 2489 38637 2492
rect 38637 2489 38671 2492
rect 38671 2489 38680 2492
rect 38628 2451 38680 2489
rect 38628 2440 38637 2451
rect 38637 2440 38671 2451
rect 38671 2440 38680 2451
rect 38628 2417 38637 2428
rect 38637 2417 38671 2428
rect 38671 2417 38680 2428
rect 38628 2379 38680 2417
rect 38628 2376 38637 2379
rect 38637 2376 38671 2379
rect 38671 2376 38680 2379
rect 38628 2345 38637 2364
rect 38637 2345 38671 2364
rect 38671 2345 38680 2364
rect 38628 2312 38680 2345
rect 38628 2273 38637 2300
rect 38637 2273 38671 2300
rect 38671 2273 38680 2300
rect 38628 2248 38680 2273
rect 38628 2235 38680 2236
rect 38628 2201 38637 2235
rect 38637 2201 38671 2235
rect 38671 2201 38680 2235
rect 38628 2184 38680 2201
rect 38628 2163 38680 2172
rect 38628 2129 38637 2163
rect 38637 2129 38671 2163
rect 38671 2129 38680 2163
rect 38628 2120 38680 2129
rect 38628 2091 38680 2108
rect 38628 2057 38637 2091
rect 38637 2057 38671 2091
rect 38671 2057 38680 2091
rect 38628 2056 38680 2057
rect 38628 2019 38680 2044
rect 38628 1992 38637 2019
rect 38637 1992 38671 2019
rect 38671 1992 38680 2019
rect 38628 1947 38680 1980
rect 38628 1928 38637 1947
rect 38637 1928 38671 1947
rect 38671 1928 38680 1947
rect 38628 1913 38637 1916
rect 38637 1913 38671 1916
rect 38671 1913 38680 1916
rect 38628 1875 38680 1913
rect 38628 1864 38637 1875
rect 38637 1864 38671 1875
rect 38671 1864 38680 1875
rect 38628 1841 38637 1852
rect 38637 1841 38671 1852
rect 38671 1841 38680 1852
rect 38628 1803 38680 1841
rect 38628 1800 38637 1803
rect 38637 1800 38671 1803
rect 38671 1800 38680 1803
rect 38628 1769 38637 1788
rect 38637 1769 38671 1788
rect 38671 1769 38680 1788
rect 38628 1736 38680 1769
rect 38628 1697 38637 1724
rect 38637 1697 38671 1724
rect 38671 1697 38680 1724
rect 38628 1672 38680 1697
rect 38628 1659 38680 1660
rect 38628 1625 38637 1659
rect 38637 1625 38671 1659
rect 38671 1625 38680 1659
rect 38628 1608 38680 1625
rect 38628 1587 38680 1596
rect 38628 1553 38637 1587
rect 38637 1553 38671 1587
rect 38671 1553 38680 1587
rect 38628 1544 38680 1553
rect 38628 1515 38680 1532
rect 38628 1481 38637 1515
rect 38637 1481 38671 1515
rect 38671 1481 38680 1515
rect 38628 1480 38680 1481
rect 38628 1443 38680 1468
rect 38628 1416 38637 1443
rect 38637 1416 38671 1443
rect 38671 1416 38680 1443
rect 38628 1371 38680 1404
rect 38628 1352 38637 1371
rect 38637 1352 38671 1371
rect 38671 1352 38680 1371
rect 38628 1337 38637 1340
rect 38637 1337 38671 1340
rect 38671 1337 38680 1340
rect 38628 1299 38680 1337
rect 38628 1288 38637 1299
rect 38637 1288 38671 1299
rect 38671 1288 38680 1299
rect 38628 1265 38637 1276
rect 38637 1265 38671 1276
rect 38671 1265 38680 1276
rect 38628 1227 38680 1265
rect 38628 1224 38637 1227
rect 38637 1224 38671 1227
rect 38671 1224 38680 1227
rect 38628 1193 38637 1212
rect 38637 1193 38671 1212
rect 38671 1193 38680 1212
rect 38628 1160 38680 1193
<< metal2 >>
rect 29025 3133 29083 3147
rect 29025 3081 29028 3133
rect 29080 3081 29083 3133
rect 29025 3069 29083 3081
rect 29025 3017 29028 3069
rect 29080 3017 29083 3069
rect 29025 3005 29083 3017
rect 29025 2953 29028 3005
rect 29080 2953 29083 3005
rect 29025 2941 29083 2953
rect 29025 2889 29028 2941
rect 29080 2889 29083 2941
rect 29025 2877 29083 2889
rect 29025 2825 29028 2877
rect 29080 2825 29083 2877
rect 29025 2813 29083 2825
rect 29025 2761 29028 2813
rect 29080 2761 29083 2813
rect 29025 2749 29083 2761
rect 29025 2697 29028 2749
rect 29080 2697 29083 2749
rect 29025 2685 29083 2697
rect 29025 2633 29028 2685
rect 29080 2633 29083 2685
rect 29025 2621 29083 2633
rect 29025 2569 29028 2621
rect 29080 2569 29083 2621
rect 29025 2557 29083 2569
rect 29025 2505 29028 2557
rect 29080 2505 29083 2557
rect 29025 2493 29083 2505
rect 29025 2441 29028 2493
rect 29080 2441 29083 2493
rect 29025 2429 29083 2441
rect 29025 2377 29028 2429
rect 29080 2377 29083 2429
rect 29025 2365 29083 2377
rect 29025 2313 29028 2365
rect 29080 2313 29083 2365
rect 29025 2301 29083 2313
rect 29025 2249 29028 2301
rect 29080 2249 29083 2301
rect 29025 2237 29083 2249
rect 29025 2185 29028 2237
rect 29080 2185 29083 2237
rect 29025 2173 29083 2185
rect 29025 2121 29028 2173
rect 29080 2121 29083 2173
rect 29025 2109 29083 2121
rect 29025 2057 29028 2109
rect 29080 2057 29083 2109
rect 29025 2045 29083 2057
rect 29025 1993 29028 2045
rect 29080 1993 29083 2045
rect 29025 1981 29083 1993
rect 29025 1929 29028 1981
rect 29080 1929 29083 1981
rect 29025 1917 29083 1929
rect 29025 1865 29028 1917
rect 29080 1865 29083 1917
rect 29025 1853 29083 1865
rect 29025 1801 29028 1853
rect 29080 1801 29083 1853
rect 29025 1789 29083 1801
rect 29025 1737 29028 1789
rect 29080 1737 29083 1789
rect 29025 1725 29083 1737
rect 29025 1673 29028 1725
rect 29080 1673 29083 1725
rect 29025 1661 29083 1673
rect 29025 1609 29028 1661
rect 29080 1609 29083 1661
rect 29025 1597 29083 1609
rect 29025 1545 29028 1597
rect 29080 1545 29083 1597
rect 29025 1533 29083 1545
rect 29025 1481 29028 1533
rect 29080 1481 29083 1533
rect 29025 1469 29083 1481
rect 29025 1417 29028 1469
rect 29080 1417 29083 1469
rect 29025 1405 29083 1417
rect 29025 1353 29028 1405
rect 29080 1353 29083 1405
rect 29025 1341 29083 1353
rect 29025 1289 29028 1341
rect 29080 1289 29083 1341
rect 29025 1277 29083 1289
rect 29025 1225 29028 1277
rect 29080 1225 29083 1277
rect 29025 1213 29083 1225
rect 29025 1161 29028 1213
rect 29080 1161 29083 1213
rect 29025 830 29083 1161
rect 29121 3135 29179 3147
rect 29121 3079 29122 3135
rect 29178 3079 29179 3135
rect 29121 3069 29179 3079
rect 29121 3055 29124 3069
rect 29176 3055 29179 3069
rect 29121 2999 29122 3055
rect 29178 2999 29179 3055
rect 29121 2975 29124 2999
rect 29176 2975 29179 2999
rect 29121 2919 29122 2975
rect 29178 2919 29179 2975
rect 29121 2895 29124 2919
rect 29176 2895 29179 2919
rect 29121 2839 29122 2895
rect 29178 2839 29179 2895
rect 29121 2825 29124 2839
rect 29176 2825 29179 2839
rect 29121 2815 29179 2825
rect 29121 2759 29122 2815
rect 29178 2759 29179 2815
rect 29121 2749 29179 2759
rect 29121 2735 29124 2749
rect 29176 2735 29179 2749
rect 29121 2679 29122 2735
rect 29178 2679 29179 2735
rect 29121 2655 29124 2679
rect 29176 2655 29179 2679
rect 29121 2599 29122 2655
rect 29178 2599 29179 2655
rect 29121 2575 29124 2599
rect 29176 2575 29179 2599
rect 29121 2519 29122 2575
rect 29178 2519 29179 2575
rect 29121 2505 29124 2519
rect 29176 2505 29179 2519
rect 29121 2495 29179 2505
rect 29121 2439 29122 2495
rect 29178 2439 29179 2495
rect 29121 2429 29179 2439
rect 29121 2415 29124 2429
rect 29176 2415 29179 2429
rect 29121 2359 29122 2415
rect 29178 2359 29179 2415
rect 29121 2335 29124 2359
rect 29176 2335 29179 2359
rect 29121 2279 29122 2335
rect 29178 2279 29179 2335
rect 29121 2255 29124 2279
rect 29176 2255 29179 2279
rect 29121 2199 29122 2255
rect 29178 2199 29179 2255
rect 29121 2185 29124 2199
rect 29176 2185 29179 2199
rect 29121 2175 29179 2185
rect 29121 2119 29122 2175
rect 29178 2119 29179 2175
rect 29121 2109 29179 2119
rect 29121 2095 29124 2109
rect 29176 2095 29179 2109
rect 29121 2039 29122 2095
rect 29178 2039 29179 2095
rect 29121 2015 29124 2039
rect 29176 2015 29179 2039
rect 29121 1959 29122 2015
rect 29178 1959 29179 2015
rect 29121 1935 29124 1959
rect 29176 1935 29179 1959
rect 29121 1879 29122 1935
rect 29178 1879 29179 1935
rect 29121 1865 29124 1879
rect 29176 1865 29179 1879
rect 29121 1855 29179 1865
rect 29121 1799 29122 1855
rect 29178 1799 29179 1855
rect 29121 1789 29179 1799
rect 29121 1775 29124 1789
rect 29176 1775 29179 1789
rect 29121 1719 29122 1775
rect 29178 1719 29179 1775
rect 29121 1695 29124 1719
rect 29176 1695 29179 1719
rect 29121 1639 29122 1695
rect 29178 1639 29179 1695
rect 29121 1615 29124 1639
rect 29176 1615 29179 1639
rect 29121 1559 29122 1615
rect 29178 1559 29179 1615
rect 29121 1545 29124 1559
rect 29176 1545 29179 1559
rect 29121 1535 29179 1545
rect 29121 1479 29122 1535
rect 29178 1479 29179 1535
rect 29121 1469 29179 1479
rect 29121 1455 29124 1469
rect 29176 1455 29179 1469
rect 29121 1399 29122 1455
rect 29178 1399 29179 1455
rect 29121 1375 29124 1399
rect 29176 1375 29179 1399
rect 29121 1319 29122 1375
rect 29178 1319 29179 1375
rect 29121 1295 29124 1319
rect 29176 1295 29179 1319
rect 29121 1239 29122 1295
rect 29178 1239 29179 1295
rect 29121 1225 29124 1239
rect 29176 1225 29179 1239
rect 29121 1215 29179 1225
rect 29121 1159 29122 1215
rect 29178 1159 29179 1215
rect 29121 1147 29179 1159
rect 29217 3133 29275 3147
rect 29217 3081 29220 3133
rect 29272 3081 29275 3133
rect 29217 3069 29275 3081
rect 29217 3017 29220 3069
rect 29272 3017 29275 3069
rect 29217 3005 29275 3017
rect 29217 2953 29220 3005
rect 29272 2953 29275 3005
rect 29217 2941 29275 2953
rect 29217 2889 29220 2941
rect 29272 2889 29275 2941
rect 29217 2877 29275 2889
rect 29217 2825 29220 2877
rect 29272 2825 29275 2877
rect 29217 2813 29275 2825
rect 29217 2761 29220 2813
rect 29272 2761 29275 2813
rect 29217 2749 29275 2761
rect 29217 2697 29220 2749
rect 29272 2697 29275 2749
rect 29217 2685 29275 2697
rect 29217 2633 29220 2685
rect 29272 2633 29275 2685
rect 29217 2621 29275 2633
rect 29217 2569 29220 2621
rect 29272 2569 29275 2621
rect 29217 2557 29275 2569
rect 29217 2505 29220 2557
rect 29272 2505 29275 2557
rect 29217 2493 29275 2505
rect 29217 2441 29220 2493
rect 29272 2441 29275 2493
rect 29217 2429 29275 2441
rect 29217 2377 29220 2429
rect 29272 2377 29275 2429
rect 29217 2365 29275 2377
rect 29217 2313 29220 2365
rect 29272 2313 29275 2365
rect 29217 2301 29275 2313
rect 29217 2249 29220 2301
rect 29272 2249 29275 2301
rect 29217 2237 29275 2249
rect 29217 2185 29220 2237
rect 29272 2185 29275 2237
rect 29217 2173 29275 2185
rect 29217 2121 29220 2173
rect 29272 2121 29275 2173
rect 29217 2109 29275 2121
rect 29217 2057 29220 2109
rect 29272 2057 29275 2109
rect 29217 2045 29275 2057
rect 29217 1993 29220 2045
rect 29272 1993 29275 2045
rect 29217 1981 29275 1993
rect 29217 1929 29220 1981
rect 29272 1929 29275 1981
rect 29217 1917 29275 1929
rect 29217 1865 29220 1917
rect 29272 1865 29275 1917
rect 29217 1853 29275 1865
rect 29217 1801 29220 1853
rect 29272 1801 29275 1853
rect 29217 1789 29275 1801
rect 29217 1737 29220 1789
rect 29272 1737 29275 1789
rect 29217 1725 29275 1737
rect 29217 1673 29220 1725
rect 29272 1673 29275 1725
rect 29217 1661 29275 1673
rect 29217 1609 29220 1661
rect 29272 1609 29275 1661
rect 29217 1597 29275 1609
rect 29217 1545 29220 1597
rect 29272 1545 29275 1597
rect 29217 1533 29275 1545
rect 29217 1481 29220 1533
rect 29272 1481 29275 1533
rect 29217 1469 29275 1481
rect 29217 1417 29220 1469
rect 29272 1417 29275 1469
rect 29217 1405 29275 1417
rect 29217 1353 29220 1405
rect 29272 1353 29275 1405
rect 29217 1341 29275 1353
rect 29217 1289 29220 1341
rect 29272 1289 29275 1341
rect 29217 1277 29275 1289
rect 29217 1225 29220 1277
rect 29272 1225 29275 1277
rect 29217 1213 29275 1225
rect 29217 1161 29220 1213
rect 29272 1161 29275 1213
rect 29217 830 29275 1161
rect 29313 3135 29371 3147
rect 29313 3079 29314 3135
rect 29370 3079 29371 3135
rect 29313 3069 29371 3079
rect 29313 3055 29316 3069
rect 29368 3055 29371 3069
rect 29313 2999 29314 3055
rect 29370 2999 29371 3055
rect 29313 2975 29316 2999
rect 29368 2975 29371 2999
rect 29313 2919 29314 2975
rect 29370 2919 29371 2975
rect 29313 2895 29316 2919
rect 29368 2895 29371 2919
rect 29313 2839 29314 2895
rect 29370 2839 29371 2895
rect 29313 2825 29316 2839
rect 29368 2825 29371 2839
rect 29313 2815 29371 2825
rect 29313 2759 29314 2815
rect 29370 2759 29371 2815
rect 29313 2749 29371 2759
rect 29313 2735 29316 2749
rect 29368 2735 29371 2749
rect 29313 2679 29314 2735
rect 29370 2679 29371 2735
rect 29313 2655 29316 2679
rect 29368 2655 29371 2679
rect 29313 2599 29314 2655
rect 29370 2599 29371 2655
rect 29313 2575 29316 2599
rect 29368 2575 29371 2599
rect 29313 2519 29314 2575
rect 29370 2519 29371 2575
rect 29313 2505 29316 2519
rect 29368 2505 29371 2519
rect 29313 2495 29371 2505
rect 29313 2439 29314 2495
rect 29370 2439 29371 2495
rect 29313 2429 29371 2439
rect 29313 2415 29316 2429
rect 29368 2415 29371 2429
rect 29313 2359 29314 2415
rect 29370 2359 29371 2415
rect 29313 2335 29316 2359
rect 29368 2335 29371 2359
rect 29313 2279 29314 2335
rect 29370 2279 29371 2335
rect 29313 2255 29316 2279
rect 29368 2255 29371 2279
rect 29313 2199 29314 2255
rect 29370 2199 29371 2255
rect 29313 2185 29316 2199
rect 29368 2185 29371 2199
rect 29313 2175 29371 2185
rect 29313 2119 29314 2175
rect 29370 2119 29371 2175
rect 29313 2109 29371 2119
rect 29313 2095 29316 2109
rect 29368 2095 29371 2109
rect 29313 2039 29314 2095
rect 29370 2039 29371 2095
rect 29313 2015 29316 2039
rect 29368 2015 29371 2039
rect 29313 1959 29314 2015
rect 29370 1959 29371 2015
rect 29313 1935 29316 1959
rect 29368 1935 29371 1959
rect 29313 1879 29314 1935
rect 29370 1879 29371 1935
rect 29313 1865 29316 1879
rect 29368 1865 29371 1879
rect 29313 1855 29371 1865
rect 29313 1799 29314 1855
rect 29370 1799 29371 1855
rect 29313 1789 29371 1799
rect 29313 1775 29316 1789
rect 29368 1775 29371 1789
rect 29313 1719 29314 1775
rect 29370 1719 29371 1775
rect 29313 1695 29316 1719
rect 29368 1695 29371 1719
rect 29313 1639 29314 1695
rect 29370 1639 29371 1695
rect 29313 1615 29316 1639
rect 29368 1615 29371 1639
rect 29313 1559 29314 1615
rect 29370 1559 29371 1615
rect 29313 1545 29316 1559
rect 29368 1545 29371 1559
rect 29313 1535 29371 1545
rect 29313 1479 29314 1535
rect 29370 1479 29371 1535
rect 29313 1469 29371 1479
rect 29313 1455 29316 1469
rect 29368 1455 29371 1469
rect 29313 1399 29314 1455
rect 29370 1399 29371 1455
rect 29313 1375 29316 1399
rect 29368 1375 29371 1399
rect 29313 1319 29314 1375
rect 29370 1319 29371 1375
rect 29313 1295 29316 1319
rect 29368 1295 29371 1319
rect 29313 1239 29314 1295
rect 29370 1239 29371 1295
rect 29313 1225 29316 1239
rect 29368 1225 29371 1239
rect 29313 1215 29371 1225
rect 29313 1159 29314 1215
rect 29370 1159 29371 1215
rect 29313 1147 29371 1159
rect 29409 3133 29467 3147
rect 29409 3081 29412 3133
rect 29464 3081 29467 3133
rect 29409 3069 29467 3081
rect 29409 3017 29412 3069
rect 29464 3017 29467 3069
rect 29409 3005 29467 3017
rect 29409 2953 29412 3005
rect 29464 2953 29467 3005
rect 29409 2941 29467 2953
rect 29409 2889 29412 2941
rect 29464 2889 29467 2941
rect 29409 2877 29467 2889
rect 29409 2825 29412 2877
rect 29464 2825 29467 2877
rect 29409 2813 29467 2825
rect 29409 2761 29412 2813
rect 29464 2761 29467 2813
rect 29409 2749 29467 2761
rect 29409 2697 29412 2749
rect 29464 2697 29467 2749
rect 29409 2685 29467 2697
rect 29409 2633 29412 2685
rect 29464 2633 29467 2685
rect 29409 2621 29467 2633
rect 29409 2569 29412 2621
rect 29464 2569 29467 2621
rect 29409 2557 29467 2569
rect 29409 2505 29412 2557
rect 29464 2505 29467 2557
rect 29409 2493 29467 2505
rect 29409 2441 29412 2493
rect 29464 2441 29467 2493
rect 29409 2429 29467 2441
rect 29409 2377 29412 2429
rect 29464 2377 29467 2429
rect 29409 2365 29467 2377
rect 29409 2313 29412 2365
rect 29464 2313 29467 2365
rect 29409 2301 29467 2313
rect 29409 2249 29412 2301
rect 29464 2249 29467 2301
rect 29409 2237 29467 2249
rect 29409 2185 29412 2237
rect 29464 2185 29467 2237
rect 29409 2173 29467 2185
rect 29409 2121 29412 2173
rect 29464 2121 29467 2173
rect 29409 2109 29467 2121
rect 29409 2057 29412 2109
rect 29464 2057 29467 2109
rect 29409 2045 29467 2057
rect 29409 1993 29412 2045
rect 29464 1993 29467 2045
rect 29409 1981 29467 1993
rect 29409 1929 29412 1981
rect 29464 1929 29467 1981
rect 29409 1917 29467 1929
rect 29409 1865 29412 1917
rect 29464 1865 29467 1917
rect 29409 1853 29467 1865
rect 29409 1801 29412 1853
rect 29464 1801 29467 1853
rect 29409 1789 29467 1801
rect 29409 1737 29412 1789
rect 29464 1737 29467 1789
rect 29409 1725 29467 1737
rect 29409 1673 29412 1725
rect 29464 1673 29467 1725
rect 29409 1661 29467 1673
rect 29409 1609 29412 1661
rect 29464 1609 29467 1661
rect 29409 1597 29467 1609
rect 29409 1545 29412 1597
rect 29464 1545 29467 1597
rect 29409 1533 29467 1545
rect 29409 1481 29412 1533
rect 29464 1481 29467 1533
rect 29409 1469 29467 1481
rect 29409 1417 29412 1469
rect 29464 1417 29467 1469
rect 29409 1405 29467 1417
rect 29409 1353 29412 1405
rect 29464 1353 29467 1405
rect 29409 1341 29467 1353
rect 29409 1289 29412 1341
rect 29464 1289 29467 1341
rect 29409 1277 29467 1289
rect 29409 1225 29412 1277
rect 29464 1225 29467 1277
rect 29409 1213 29467 1225
rect 29409 1161 29412 1213
rect 29464 1161 29467 1213
rect 29409 830 29467 1161
rect 29505 3135 29563 3147
rect 29505 3079 29506 3135
rect 29562 3079 29563 3135
rect 29505 3069 29563 3079
rect 29505 3055 29508 3069
rect 29560 3055 29563 3069
rect 29505 2999 29506 3055
rect 29562 2999 29563 3055
rect 29505 2975 29508 2999
rect 29560 2975 29563 2999
rect 29505 2919 29506 2975
rect 29562 2919 29563 2975
rect 29505 2895 29508 2919
rect 29560 2895 29563 2919
rect 29505 2839 29506 2895
rect 29562 2839 29563 2895
rect 29505 2825 29508 2839
rect 29560 2825 29563 2839
rect 29505 2815 29563 2825
rect 29505 2759 29506 2815
rect 29562 2759 29563 2815
rect 29505 2749 29563 2759
rect 29505 2735 29508 2749
rect 29560 2735 29563 2749
rect 29505 2679 29506 2735
rect 29562 2679 29563 2735
rect 29505 2655 29508 2679
rect 29560 2655 29563 2679
rect 29505 2599 29506 2655
rect 29562 2599 29563 2655
rect 29505 2575 29508 2599
rect 29560 2575 29563 2599
rect 29505 2519 29506 2575
rect 29562 2519 29563 2575
rect 29505 2505 29508 2519
rect 29560 2505 29563 2519
rect 29505 2495 29563 2505
rect 29505 2439 29506 2495
rect 29562 2439 29563 2495
rect 29505 2429 29563 2439
rect 29505 2415 29508 2429
rect 29560 2415 29563 2429
rect 29505 2359 29506 2415
rect 29562 2359 29563 2415
rect 29505 2335 29508 2359
rect 29560 2335 29563 2359
rect 29505 2279 29506 2335
rect 29562 2279 29563 2335
rect 29505 2255 29508 2279
rect 29560 2255 29563 2279
rect 29505 2199 29506 2255
rect 29562 2199 29563 2255
rect 29505 2185 29508 2199
rect 29560 2185 29563 2199
rect 29505 2175 29563 2185
rect 29505 2119 29506 2175
rect 29562 2119 29563 2175
rect 29505 2109 29563 2119
rect 29505 2095 29508 2109
rect 29560 2095 29563 2109
rect 29505 2039 29506 2095
rect 29562 2039 29563 2095
rect 29505 2015 29508 2039
rect 29560 2015 29563 2039
rect 29505 1959 29506 2015
rect 29562 1959 29563 2015
rect 29505 1935 29508 1959
rect 29560 1935 29563 1959
rect 29505 1879 29506 1935
rect 29562 1879 29563 1935
rect 29505 1865 29508 1879
rect 29560 1865 29563 1879
rect 29505 1855 29563 1865
rect 29505 1799 29506 1855
rect 29562 1799 29563 1855
rect 29505 1789 29563 1799
rect 29505 1775 29508 1789
rect 29560 1775 29563 1789
rect 29505 1719 29506 1775
rect 29562 1719 29563 1775
rect 29505 1695 29508 1719
rect 29560 1695 29563 1719
rect 29505 1639 29506 1695
rect 29562 1639 29563 1695
rect 29505 1615 29508 1639
rect 29560 1615 29563 1639
rect 29505 1559 29506 1615
rect 29562 1559 29563 1615
rect 29505 1545 29508 1559
rect 29560 1545 29563 1559
rect 29505 1535 29563 1545
rect 29505 1479 29506 1535
rect 29562 1479 29563 1535
rect 29505 1469 29563 1479
rect 29505 1455 29508 1469
rect 29560 1455 29563 1469
rect 29505 1399 29506 1455
rect 29562 1399 29563 1455
rect 29505 1375 29508 1399
rect 29560 1375 29563 1399
rect 29505 1319 29506 1375
rect 29562 1319 29563 1375
rect 29505 1295 29508 1319
rect 29560 1295 29563 1319
rect 29505 1239 29506 1295
rect 29562 1239 29563 1295
rect 29505 1225 29508 1239
rect 29560 1225 29563 1239
rect 29505 1215 29563 1225
rect 29505 1159 29506 1215
rect 29562 1159 29563 1215
rect 29505 1147 29563 1159
rect 29601 3133 29659 3147
rect 29601 3081 29604 3133
rect 29656 3081 29659 3133
rect 29601 3069 29659 3081
rect 29601 3017 29604 3069
rect 29656 3017 29659 3069
rect 29601 3005 29659 3017
rect 29601 2953 29604 3005
rect 29656 2953 29659 3005
rect 29601 2941 29659 2953
rect 29601 2889 29604 2941
rect 29656 2889 29659 2941
rect 29601 2877 29659 2889
rect 29601 2825 29604 2877
rect 29656 2825 29659 2877
rect 29601 2813 29659 2825
rect 29601 2761 29604 2813
rect 29656 2761 29659 2813
rect 29601 2749 29659 2761
rect 29601 2697 29604 2749
rect 29656 2697 29659 2749
rect 29601 2685 29659 2697
rect 29601 2633 29604 2685
rect 29656 2633 29659 2685
rect 29601 2621 29659 2633
rect 29601 2569 29604 2621
rect 29656 2569 29659 2621
rect 29601 2557 29659 2569
rect 29601 2505 29604 2557
rect 29656 2505 29659 2557
rect 29601 2493 29659 2505
rect 29601 2441 29604 2493
rect 29656 2441 29659 2493
rect 29601 2429 29659 2441
rect 29601 2377 29604 2429
rect 29656 2377 29659 2429
rect 29601 2365 29659 2377
rect 29601 2313 29604 2365
rect 29656 2313 29659 2365
rect 29601 2301 29659 2313
rect 29601 2249 29604 2301
rect 29656 2249 29659 2301
rect 29601 2237 29659 2249
rect 29601 2185 29604 2237
rect 29656 2185 29659 2237
rect 29601 2173 29659 2185
rect 29601 2121 29604 2173
rect 29656 2121 29659 2173
rect 29601 2109 29659 2121
rect 29601 2057 29604 2109
rect 29656 2057 29659 2109
rect 29601 2045 29659 2057
rect 29601 1993 29604 2045
rect 29656 1993 29659 2045
rect 29601 1981 29659 1993
rect 29601 1929 29604 1981
rect 29656 1929 29659 1981
rect 29601 1917 29659 1929
rect 29601 1865 29604 1917
rect 29656 1865 29659 1917
rect 29601 1853 29659 1865
rect 29601 1801 29604 1853
rect 29656 1801 29659 1853
rect 29601 1789 29659 1801
rect 29601 1737 29604 1789
rect 29656 1737 29659 1789
rect 29601 1725 29659 1737
rect 29601 1673 29604 1725
rect 29656 1673 29659 1725
rect 29601 1661 29659 1673
rect 29601 1609 29604 1661
rect 29656 1609 29659 1661
rect 29601 1597 29659 1609
rect 29601 1545 29604 1597
rect 29656 1545 29659 1597
rect 29601 1533 29659 1545
rect 29601 1481 29604 1533
rect 29656 1481 29659 1533
rect 29601 1469 29659 1481
rect 29601 1417 29604 1469
rect 29656 1417 29659 1469
rect 29601 1405 29659 1417
rect 29601 1353 29604 1405
rect 29656 1353 29659 1405
rect 29601 1341 29659 1353
rect 29601 1289 29604 1341
rect 29656 1289 29659 1341
rect 29601 1277 29659 1289
rect 29601 1225 29604 1277
rect 29656 1225 29659 1277
rect 29601 1213 29659 1225
rect 29601 1161 29604 1213
rect 29656 1161 29659 1213
rect 29601 830 29659 1161
rect 29697 3135 29755 3147
rect 29697 3079 29698 3135
rect 29754 3079 29755 3135
rect 29697 3069 29755 3079
rect 29697 3055 29700 3069
rect 29752 3055 29755 3069
rect 29697 2999 29698 3055
rect 29754 2999 29755 3055
rect 29697 2975 29700 2999
rect 29752 2975 29755 2999
rect 29697 2919 29698 2975
rect 29754 2919 29755 2975
rect 29697 2895 29700 2919
rect 29752 2895 29755 2919
rect 29697 2839 29698 2895
rect 29754 2839 29755 2895
rect 29697 2825 29700 2839
rect 29752 2825 29755 2839
rect 29697 2815 29755 2825
rect 29697 2759 29698 2815
rect 29754 2759 29755 2815
rect 29697 2749 29755 2759
rect 29697 2735 29700 2749
rect 29752 2735 29755 2749
rect 29697 2679 29698 2735
rect 29754 2679 29755 2735
rect 29697 2655 29700 2679
rect 29752 2655 29755 2679
rect 29697 2599 29698 2655
rect 29754 2599 29755 2655
rect 29697 2575 29700 2599
rect 29752 2575 29755 2599
rect 29697 2519 29698 2575
rect 29754 2519 29755 2575
rect 29697 2505 29700 2519
rect 29752 2505 29755 2519
rect 29697 2495 29755 2505
rect 29697 2439 29698 2495
rect 29754 2439 29755 2495
rect 29697 2429 29755 2439
rect 29697 2415 29700 2429
rect 29752 2415 29755 2429
rect 29697 2359 29698 2415
rect 29754 2359 29755 2415
rect 29697 2335 29700 2359
rect 29752 2335 29755 2359
rect 29697 2279 29698 2335
rect 29754 2279 29755 2335
rect 29697 2255 29700 2279
rect 29752 2255 29755 2279
rect 29697 2199 29698 2255
rect 29754 2199 29755 2255
rect 29697 2185 29700 2199
rect 29752 2185 29755 2199
rect 29697 2175 29755 2185
rect 29697 2119 29698 2175
rect 29754 2119 29755 2175
rect 29697 2109 29755 2119
rect 29697 2095 29700 2109
rect 29752 2095 29755 2109
rect 29697 2039 29698 2095
rect 29754 2039 29755 2095
rect 29697 2015 29700 2039
rect 29752 2015 29755 2039
rect 29697 1959 29698 2015
rect 29754 1959 29755 2015
rect 29697 1935 29700 1959
rect 29752 1935 29755 1959
rect 29697 1879 29698 1935
rect 29754 1879 29755 1935
rect 29697 1865 29700 1879
rect 29752 1865 29755 1879
rect 29697 1855 29755 1865
rect 29697 1799 29698 1855
rect 29754 1799 29755 1855
rect 29697 1789 29755 1799
rect 29697 1775 29700 1789
rect 29752 1775 29755 1789
rect 29697 1719 29698 1775
rect 29754 1719 29755 1775
rect 29697 1695 29700 1719
rect 29752 1695 29755 1719
rect 29697 1639 29698 1695
rect 29754 1639 29755 1695
rect 29697 1615 29700 1639
rect 29752 1615 29755 1639
rect 29697 1559 29698 1615
rect 29754 1559 29755 1615
rect 29697 1545 29700 1559
rect 29752 1545 29755 1559
rect 29697 1535 29755 1545
rect 29697 1479 29698 1535
rect 29754 1479 29755 1535
rect 29697 1469 29755 1479
rect 29697 1455 29700 1469
rect 29752 1455 29755 1469
rect 29697 1399 29698 1455
rect 29754 1399 29755 1455
rect 29697 1375 29700 1399
rect 29752 1375 29755 1399
rect 29697 1319 29698 1375
rect 29754 1319 29755 1375
rect 29697 1295 29700 1319
rect 29752 1295 29755 1319
rect 29697 1239 29698 1295
rect 29754 1239 29755 1295
rect 29697 1225 29700 1239
rect 29752 1225 29755 1239
rect 29697 1215 29755 1225
rect 29697 1159 29698 1215
rect 29754 1159 29755 1215
rect 29697 1147 29755 1159
rect 29793 3133 29851 3147
rect 29793 3081 29796 3133
rect 29848 3081 29851 3133
rect 29793 3069 29851 3081
rect 29793 3017 29796 3069
rect 29848 3017 29851 3069
rect 29793 3005 29851 3017
rect 29793 2953 29796 3005
rect 29848 2953 29851 3005
rect 29793 2941 29851 2953
rect 29793 2889 29796 2941
rect 29848 2889 29851 2941
rect 29793 2877 29851 2889
rect 29793 2825 29796 2877
rect 29848 2825 29851 2877
rect 29793 2813 29851 2825
rect 29793 2761 29796 2813
rect 29848 2761 29851 2813
rect 29793 2749 29851 2761
rect 29793 2697 29796 2749
rect 29848 2697 29851 2749
rect 29793 2685 29851 2697
rect 29793 2633 29796 2685
rect 29848 2633 29851 2685
rect 29793 2621 29851 2633
rect 29793 2569 29796 2621
rect 29848 2569 29851 2621
rect 29793 2557 29851 2569
rect 29793 2505 29796 2557
rect 29848 2505 29851 2557
rect 29793 2493 29851 2505
rect 29793 2441 29796 2493
rect 29848 2441 29851 2493
rect 29793 2429 29851 2441
rect 29793 2377 29796 2429
rect 29848 2377 29851 2429
rect 29793 2365 29851 2377
rect 29793 2313 29796 2365
rect 29848 2313 29851 2365
rect 29793 2301 29851 2313
rect 29793 2249 29796 2301
rect 29848 2249 29851 2301
rect 29793 2237 29851 2249
rect 29793 2185 29796 2237
rect 29848 2185 29851 2237
rect 29793 2173 29851 2185
rect 29793 2121 29796 2173
rect 29848 2121 29851 2173
rect 29793 2109 29851 2121
rect 29793 2057 29796 2109
rect 29848 2057 29851 2109
rect 29793 2045 29851 2057
rect 29793 1993 29796 2045
rect 29848 1993 29851 2045
rect 29793 1981 29851 1993
rect 29793 1929 29796 1981
rect 29848 1929 29851 1981
rect 29793 1917 29851 1929
rect 29793 1865 29796 1917
rect 29848 1865 29851 1917
rect 29793 1853 29851 1865
rect 29793 1801 29796 1853
rect 29848 1801 29851 1853
rect 29793 1789 29851 1801
rect 29793 1737 29796 1789
rect 29848 1737 29851 1789
rect 29793 1725 29851 1737
rect 29793 1673 29796 1725
rect 29848 1673 29851 1725
rect 29793 1661 29851 1673
rect 29793 1609 29796 1661
rect 29848 1609 29851 1661
rect 29793 1597 29851 1609
rect 29793 1545 29796 1597
rect 29848 1545 29851 1597
rect 29793 1533 29851 1545
rect 29793 1481 29796 1533
rect 29848 1481 29851 1533
rect 29793 1469 29851 1481
rect 29793 1417 29796 1469
rect 29848 1417 29851 1469
rect 29793 1405 29851 1417
rect 29793 1353 29796 1405
rect 29848 1353 29851 1405
rect 29793 1341 29851 1353
rect 29793 1289 29796 1341
rect 29848 1289 29851 1341
rect 29793 1277 29851 1289
rect 29793 1225 29796 1277
rect 29848 1225 29851 1277
rect 29793 1213 29851 1225
rect 29793 1161 29796 1213
rect 29848 1161 29851 1213
rect 29793 830 29851 1161
rect 29889 3135 29947 3147
rect 29889 3079 29890 3135
rect 29946 3079 29947 3135
rect 29889 3069 29947 3079
rect 29889 3055 29892 3069
rect 29944 3055 29947 3069
rect 29889 2999 29890 3055
rect 29946 2999 29947 3055
rect 29889 2975 29892 2999
rect 29944 2975 29947 2999
rect 29889 2919 29890 2975
rect 29946 2919 29947 2975
rect 29889 2895 29892 2919
rect 29944 2895 29947 2919
rect 29889 2839 29890 2895
rect 29946 2839 29947 2895
rect 29889 2825 29892 2839
rect 29944 2825 29947 2839
rect 29889 2815 29947 2825
rect 29889 2759 29890 2815
rect 29946 2759 29947 2815
rect 29889 2749 29947 2759
rect 29889 2735 29892 2749
rect 29944 2735 29947 2749
rect 29889 2679 29890 2735
rect 29946 2679 29947 2735
rect 29889 2655 29892 2679
rect 29944 2655 29947 2679
rect 29889 2599 29890 2655
rect 29946 2599 29947 2655
rect 29889 2575 29892 2599
rect 29944 2575 29947 2599
rect 29889 2519 29890 2575
rect 29946 2519 29947 2575
rect 29889 2505 29892 2519
rect 29944 2505 29947 2519
rect 29889 2495 29947 2505
rect 29889 2439 29890 2495
rect 29946 2439 29947 2495
rect 29889 2429 29947 2439
rect 29889 2415 29892 2429
rect 29944 2415 29947 2429
rect 29889 2359 29890 2415
rect 29946 2359 29947 2415
rect 29889 2335 29892 2359
rect 29944 2335 29947 2359
rect 29889 2279 29890 2335
rect 29946 2279 29947 2335
rect 29889 2255 29892 2279
rect 29944 2255 29947 2279
rect 29889 2199 29890 2255
rect 29946 2199 29947 2255
rect 29889 2185 29892 2199
rect 29944 2185 29947 2199
rect 29889 2175 29947 2185
rect 29889 2119 29890 2175
rect 29946 2119 29947 2175
rect 29889 2109 29947 2119
rect 29889 2095 29892 2109
rect 29944 2095 29947 2109
rect 29889 2039 29890 2095
rect 29946 2039 29947 2095
rect 29889 2015 29892 2039
rect 29944 2015 29947 2039
rect 29889 1959 29890 2015
rect 29946 1959 29947 2015
rect 29889 1935 29892 1959
rect 29944 1935 29947 1959
rect 29889 1879 29890 1935
rect 29946 1879 29947 1935
rect 29889 1865 29892 1879
rect 29944 1865 29947 1879
rect 29889 1855 29947 1865
rect 29889 1799 29890 1855
rect 29946 1799 29947 1855
rect 29889 1789 29947 1799
rect 29889 1775 29892 1789
rect 29944 1775 29947 1789
rect 29889 1719 29890 1775
rect 29946 1719 29947 1775
rect 29889 1695 29892 1719
rect 29944 1695 29947 1719
rect 29889 1639 29890 1695
rect 29946 1639 29947 1695
rect 29889 1615 29892 1639
rect 29944 1615 29947 1639
rect 29889 1559 29890 1615
rect 29946 1559 29947 1615
rect 29889 1545 29892 1559
rect 29944 1545 29947 1559
rect 29889 1535 29947 1545
rect 29889 1479 29890 1535
rect 29946 1479 29947 1535
rect 29889 1469 29947 1479
rect 29889 1455 29892 1469
rect 29944 1455 29947 1469
rect 29889 1399 29890 1455
rect 29946 1399 29947 1455
rect 29889 1375 29892 1399
rect 29944 1375 29947 1399
rect 29889 1319 29890 1375
rect 29946 1319 29947 1375
rect 29889 1295 29892 1319
rect 29944 1295 29947 1319
rect 29889 1239 29890 1295
rect 29946 1239 29947 1295
rect 29889 1225 29892 1239
rect 29944 1225 29947 1239
rect 29889 1215 29947 1225
rect 29889 1159 29890 1215
rect 29946 1159 29947 1215
rect 29889 1147 29947 1159
rect 29985 3133 30043 3147
rect 29985 3081 29988 3133
rect 30040 3081 30043 3133
rect 29985 3069 30043 3081
rect 29985 3017 29988 3069
rect 30040 3017 30043 3069
rect 29985 3005 30043 3017
rect 29985 2953 29988 3005
rect 30040 2953 30043 3005
rect 29985 2941 30043 2953
rect 29985 2889 29988 2941
rect 30040 2889 30043 2941
rect 29985 2877 30043 2889
rect 29985 2825 29988 2877
rect 30040 2825 30043 2877
rect 29985 2813 30043 2825
rect 29985 2761 29988 2813
rect 30040 2761 30043 2813
rect 29985 2749 30043 2761
rect 29985 2697 29988 2749
rect 30040 2697 30043 2749
rect 29985 2685 30043 2697
rect 29985 2633 29988 2685
rect 30040 2633 30043 2685
rect 29985 2621 30043 2633
rect 29985 2569 29988 2621
rect 30040 2569 30043 2621
rect 29985 2557 30043 2569
rect 29985 2505 29988 2557
rect 30040 2505 30043 2557
rect 29985 2493 30043 2505
rect 29985 2441 29988 2493
rect 30040 2441 30043 2493
rect 29985 2429 30043 2441
rect 29985 2377 29988 2429
rect 30040 2377 30043 2429
rect 29985 2365 30043 2377
rect 29985 2313 29988 2365
rect 30040 2313 30043 2365
rect 29985 2301 30043 2313
rect 29985 2249 29988 2301
rect 30040 2249 30043 2301
rect 29985 2237 30043 2249
rect 29985 2185 29988 2237
rect 30040 2185 30043 2237
rect 29985 2173 30043 2185
rect 29985 2121 29988 2173
rect 30040 2121 30043 2173
rect 29985 2109 30043 2121
rect 29985 2057 29988 2109
rect 30040 2057 30043 2109
rect 29985 2045 30043 2057
rect 29985 1993 29988 2045
rect 30040 1993 30043 2045
rect 29985 1981 30043 1993
rect 29985 1929 29988 1981
rect 30040 1929 30043 1981
rect 29985 1917 30043 1929
rect 29985 1865 29988 1917
rect 30040 1865 30043 1917
rect 29985 1853 30043 1865
rect 29985 1801 29988 1853
rect 30040 1801 30043 1853
rect 29985 1789 30043 1801
rect 29985 1737 29988 1789
rect 30040 1737 30043 1789
rect 29985 1725 30043 1737
rect 29985 1673 29988 1725
rect 30040 1673 30043 1725
rect 29985 1661 30043 1673
rect 29985 1609 29988 1661
rect 30040 1609 30043 1661
rect 29985 1597 30043 1609
rect 29985 1545 29988 1597
rect 30040 1545 30043 1597
rect 29985 1533 30043 1545
rect 29985 1481 29988 1533
rect 30040 1481 30043 1533
rect 29985 1469 30043 1481
rect 29985 1417 29988 1469
rect 30040 1417 30043 1469
rect 29985 1405 30043 1417
rect 29985 1353 29988 1405
rect 30040 1353 30043 1405
rect 29985 1341 30043 1353
rect 29985 1289 29988 1341
rect 30040 1289 30043 1341
rect 29985 1277 30043 1289
rect 29985 1225 29988 1277
rect 30040 1225 30043 1277
rect 29985 1213 30043 1225
rect 29985 1161 29988 1213
rect 30040 1161 30043 1213
rect 29985 830 30043 1161
rect 30081 3135 30139 3147
rect 30081 3079 30082 3135
rect 30138 3079 30139 3135
rect 30081 3069 30139 3079
rect 30081 3055 30084 3069
rect 30136 3055 30139 3069
rect 30081 2999 30082 3055
rect 30138 2999 30139 3055
rect 30081 2975 30084 2999
rect 30136 2975 30139 2999
rect 30081 2919 30082 2975
rect 30138 2919 30139 2975
rect 30081 2895 30084 2919
rect 30136 2895 30139 2919
rect 30081 2839 30082 2895
rect 30138 2839 30139 2895
rect 30081 2825 30084 2839
rect 30136 2825 30139 2839
rect 30081 2815 30139 2825
rect 30081 2759 30082 2815
rect 30138 2759 30139 2815
rect 30081 2749 30139 2759
rect 30081 2735 30084 2749
rect 30136 2735 30139 2749
rect 30081 2679 30082 2735
rect 30138 2679 30139 2735
rect 30081 2655 30084 2679
rect 30136 2655 30139 2679
rect 30081 2599 30082 2655
rect 30138 2599 30139 2655
rect 30081 2575 30084 2599
rect 30136 2575 30139 2599
rect 30081 2519 30082 2575
rect 30138 2519 30139 2575
rect 30081 2505 30084 2519
rect 30136 2505 30139 2519
rect 30081 2495 30139 2505
rect 30081 2439 30082 2495
rect 30138 2439 30139 2495
rect 30081 2429 30139 2439
rect 30081 2415 30084 2429
rect 30136 2415 30139 2429
rect 30081 2359 30082 2415
rect 30138 2359 30139 2415
rect 30081 2335 30084 2359
rect 30136 2335 30139 2359
rect 30081 2279 30082 2335
rect 30138 2279 30139 2335
rect 30081 2255 30084 2279
rect 30136 2255 30139 2279
rect 30081 2199 30082 2255
rect 30138 2199 30139 2255
rect 30081 2185 30084 2199
rect 30136 2185 30139 2199
rect 30081 2175 30139 2185
rect 30081 2119 30082 2175
rect 30138 2119 30139 2175
rect 30081 2109 30139 2119
rect 30081 2095 30084 2109
rect 30136 2095 30139 2109
rect 30081 2039 30082 2095
rect 30138 2039 30139 2095
rect 30081 2015 30084 2039
rect 30136 2015 30139 2039
rect 30081 1959 30082 2015
rect 30138 1959 30139 2015
rect 30081 1935 30084 1959
rect 30136 1935 30139 1959
rect 30081 1879 30082 1935
rect 30138 1879 30139 1935
rect 30081 1865 30084 1879
rect 30136 1865 30139 1879
rect 30081 1855 30139 1865
rect 30081 1799 30082 1855
rect 30138 1799 30139 1855
rect 30081 1789 30139 1799
rect 30081 1775 30084 1789
rect 30136 1775 30139 1789
rect 30081 1719 30082 1775
rect 30138 1719 30139 1775
rect 30081 1695 30084 1719
rect 30136 1695 30139 1719
rect 30081 1639 30082 1695
rect 30138 1639 30139 1695
rect 30081 1615 30084 1639
rect 30136 1615 30139 1639
rect 30081 1559 30082 1615
rect 30138 1559 30139 1615
rect 30081 1545 30084 1559
rect 30136 1545 30139 1559
rect 30081 1535 30139 1545
rect 30081 1479 30082 1535
rect 30138 1479 30139 1535
rect 30081 1469 30139 1479
rect 30081 1455 30084 1469
rect 30136 1455 30139 1469
rect 30081 1399 30082 1455
rect 30138 1399 30139 1455
rect 30081 1375 30084 1399
rect 30136 1375 30139 1399
rect 30081 1319 30082 1375
rect 30138 1319 30139 1375
rect 30081 1295 30084 1319
rect 30136 1295 30139 1319
rect 30081 1239 30082 1295
rect 30138 1239 30139 1295
rect 30081 1225 30084 1239
rect 30136 1225 30139 1239
rect 30081 1215 30139 1225
rect 30081 1159 30082 1215
rect 30138 1159 30139 1215
rect 30081 1147 30139 1159
rect 30177 3133 30235 3147
rect 30177 3081 30180 3133
rect 30232 3081 30235 3133
rect 30177 3069 30235 3081
rect 30177 3017 30180 3069
rect 30232 3017 30235 3069
rect 30177 3005 30235 3017
rect 30177 2953 30180 3005
rect 30232 2953 30235 3005
rect 30177 2941 30235 2953
rect 30177 2889 30180 2941
rect 30232 2889 30235 2941
rect 30177 2877 30235 2889
rect 30177 2825 30180 2877
rect 30232 2825 30235 2877
rect 30177 2813 30235 2825
rect 30177 2761 30180 2813
rect 30232 2761 30235 2813
rect 30177 2749 30235 2761
rect 30177 2697 30180 2749
rect 30232 2697 30235 2749
rect 30177 2685 30235 2697
rect 30177 2633 30180 2685
rect 30232 2633 30235 2685
rect 30177 2621 30235 2633
rect 30177 2569 30180 2621
rect 30232 2569 30235 2621
rect 30177 2557 30235 2569
rect 30177 2505 30180 2557
rect 30232 2505 30235 2557
rect 30177 2493 30235 2505
rect 30177 2441 30180 2493
rect 30232 2441 30235 2493
rect 30177 2429 30235 2441
rect 30177 2377 30180 2429
rect 30232 2377 30235 2429
rect 30177 2365 30235 2377
rect 30177 2313 30180 2365
rect 30232 2313 30235 2365
rect 30177 2301 30235 2313
rect 30177 2249 30180 2301
rect 30232 2249 30235 2301
rect 30177 2237 30235 2249
rect 30177 2185 30180 2237
rect 30232 2185 30235 2237
rect 30177 2173 30235 2185
rect 30177 2121 30180 2173
rect 30232 2121 30235 2173
rect 30177 2109 30235 2121
rect 30177 2057 30180 2109
rect 30232 2057 30235 2109
rect 30177 2045 30235 2057
rect 30177 1993 30180 2045
rect 30232 1993 30235 2045
rect 30177 1981 30235 1993
rect 30177 1929 30180 1981
rect 30232 1929 30235 1981
rect 30177 1917 30235 1929
rect 30177 1865 30180 1917
rect 30232 1865 30235 1917
rect 30177 1853 30235 1865
rect 30177 1801 30180 1853
rect 30232 1801 30235 1853
rect 30177 1789 30235 1801
rect 30177 1737 30180 1789
rect 30232 1737 30235 1789
rect 30177 1725 30235 1737
rect 30177 1673 30180 1725
rect 30232 1673 30235 1725
rect 30177 1661 30235 1673
rect 30177 1609 30180 1661
rect 30232 1609 30235 1661
rect 30177 1597 30235 1609
rect 30177 1545 30180 1597
rect 30232 1545 30235 1597
rect 30177 1533 30235 1545
rect 30177 1481 30180 1533
rect 30232 1481 30235 1533
rect 30177 1469 30235 1481
rect 30177 1417 30180 1469
rect 30232 1417 30235 1469
rect 30177 1405 30235 1417
rect 30177 1353 30180 1405
rect 30232 1353 30235 1405
rect 30177 1341 30235 1353
rect 30177 1289 30180 1341
rect 30232 1289 30235 1341
rect 30177 1277 30235 1289
rect 30177 1225 30180 1277
rect 30232 1225 30235 1277
rect 30177 1213 30235 1225
rect 30177 1161 30180 1213
rect 30232 1161 30235 1213
rect 30177 830 30235 1161
rect 30273 3135 30331 3147
rect 30273 3079 30274 3135
rect 30330 3079 30331 3135
rect 30273 3069 30331 3079
rect 30273 3055 30276 3069
rect 30328 3055 30331 3069
rect 30273 2999 30274 3055
rect 30330 2999 30331 3055
rect 30273 2975 30276 2999
rect 30328 2975 30331 2999
rect 30273 2919 30274 2975
rect 30330 2919 30331 2975
rect 30273 2895 30276 2919
rect 30328 2895 30331 2919
rect 30273 2839 30274 2895
rect 30330 2839 30331 2895
rect 30273 2825 30276 2839
rect 30328 2825 30331 2839
rect 30273 2815 30331 2825
rect 30273 2759 30274 2815
rect 30330 2759 30331 2815
rect 30273 2749 30331 2759
rect 30273 2735 30276 2749
rect 30328 2735 30331 2749
rect 30273 2679 30274 2735
rect 30330 2679 30331 2735
rect 30273 2655 30276 2679
rect 30328 2655 30331 2679
rect 30273 2599 30274 2655
rect 30330 2599 30331 2655
rect 30273 2575 30276 2599
rect 30328 2575 30331 2599
rect 30273 2519 30274 2575
rect 30330 2519 30331 2575
rect 30273 2505 30276 2519
rect 30328 2505 30331 2519
rect 30273 2495 30331 2505
rect 30273 2439 30274 2495
rect 30330 2439 30331 2495
rect 30273 2429 30331 2439
rect 30273 2415 30276 2429
rect 30328 2415 30331 2429
rect 30273 2359 30274 2415
rect 30330 2359 30331 2415
rect 30273 2335 30276 2359
rect 30328 2335 30331 2359
rect 30273 2279 30274 2335
rect 30330 2279 30331 2335
rect 30273 2255 30276 2279
rect 30328 2255 30331 2279
rect 30273 2199 30274 2255
rect 30330 2199 30331 2255
rect 30273 2185 30276 2199
rect 30328 2185 30331 2199
rect 30273 2175 30331 2185
rect 30273 2119 30274 2175
rect 30330 2119 30331 2175
rect 30273 2109 30331 2119
rect 30273 2095 30276 2109
rect 30328 2095 30331 2109
rect 30273 2039 30274 2095
rect 30330 2039 30331 2095
rect 30273 2015 30276 2039
rect 30328 2015 30331 2039
rect 30273 1959 30274 2015
rect 30330 1959 30331 2015
rect 30273 1935 30276 1959
rect 30328 1935 30331 1959
rect 30273 1879 30274 1935
rect 30330 1879 30331 1935
rect 30273 1865 30276 1879
rect 30328 1865 30331 1879
rect 30273 1855 30331 1865
rect 30273 1799 30274 1855
rect 30330 1799 30331 1855
rect 30273 1789 30331 1799
rect 30273 1775 30276 1789
rect 30328 1775 30331 1789
rect 30273 1719 30274 1775
rect 30330 1719 30331 1775
rect 30273 1695 30276 1719
rect 30328 1695 30331 1719
rect 30273 1639 30274 1695
rect 30330 1639 30331 1695
rect 30273 1615 30276 1639
rect 30328 1615 30331 1639
rect 30273 1559 30274 1615
rect 30330 1559 30331 1615
rect 30273 1545 30276 1559
rect 30328 1545 30331 1559
rect 30273 1535 30331 1545
rect 30273 1479 30274 1535
rect 30330 1479 30331 1535
rect 30273 1469 30331 1479
rect 30273 1455 30276 1469
rect 30328 1455 30331 1469
rect 30273 1399 30274 1455
rect 30330 1399 30331 1455
rect 30273 1375 30276 1399
rect 30328 1375 30331 1399
rect 30273 1319 30274 1375
rect 30330 1319 30331 1375
rect 30273 1295 30276 1319
rect 30328 1295 30331 1319
rect 30273 1239 30274 1295
rect 30330 1239 30331 1295
rect 30273 1225 30276 1239
rect 30328 1225 30331 1239
rect 30273 1215 30331 1225
rect 30273 1159 30274 1215
rect 30330 1159 30331 1215
rect 30273 1147 30331 1159
rect 30369 3133 30427 3147
rect 30369 3081 30372 3133
rect 30424 3081 30427 3133
rect 30369 3069 30427 3081
rect 30369 3017 30372 3069
rect 30424 3017 30427 3069
rect 30369 3005 30427 3017
rect 30369 2953 30372 3005
rect 30424 2953 30427 3005
rect 30369 2941 30427 2953
rect 30369 2889 30372 2941
rect 30424 2889 30427 2941
rect 30369 2877 30427 2889
rect 30369 2825 30372 2877
rect 30424 2825 30427 2877
rect 30369 2813 30427 2825
rect 30369 2761 30372 2813
rect 30424 2761 30427 2813
rect 30369 2749 30427 2761
rect 30369 2697 30372 2749
rect 30424 2697 30427 2749
rect 30369 2685 30427 2697
rect 30369 2633 30372 2685
rect 30424 2633 30427 2685
rect 30369 2621 30427 2633
rect 30369 2569 30372 2621
rect 30424 2569 30427 2621
rect 30369 2557 30427 2569
rect 30369 2505 30372 2557
rect 30424 2505 30427 2557
rect 30369 2493 30427 2505
rect 30369 2441 30372 2493
rect 30424 2441 30427 2493
rect 30369 2429 30427 2441
rect 30369 2377 30372 2429
rect 30424 2377 30427 2429
rect 30369 2365 30427 2377
rect 30369 2313 30372 2365
rect 30424 2313 30427 2365
rect 30369 2301 30427 2313
rect 30369 2249 30372 2301
rect 30424 2249 30427 2301
rect 30369 2237 30427 2249
rect 30369 2185 30372 2237
rect 30424 2185 30427 2237
rect 30369 2173 30427 2185
rect 30369 2121 30372 2173
rect 30424 2121 30427 2173
rect 30369 2109 30427 2121
rect 30369 2057 30372 2109
rect 30424 2057 30427 2109
rect 30369 2045 30427 2057
rect 30369 1993 30372 2045
rect 30424 1993 30427 2045
rect 30369 1981 30427 1993
rect 30369 1929 30372 1981
rect 30424 1929 30427 1981
rect 30369 1917 30427 1929
rect 30369 1865 30372 1917
rect 30424 1865 30427 1917
rect 30369 1853 30427 1865
rect 30369 1801 30372 1853
rect 30424 1801 30427 1853
rect 30369 1789 30427 1801
rect 30369 1737 30372 1789
rect 30424 1737 30427 1789
rect 30369 1725 30427 1737
rect 30369 1673 30372 1725
rect 30424 1673 30427 1725
rect 30369 1661 30427 1673
rect 30369 1609 30372 1661
rect 30424 1609 30427 1661
rect 30369 1597 30427 1609
rect 30369 1545 30372 1597
rect 30424 1545 30427 1597
rect 30369 1533 30427 1545
rect 30369 1481 30372 1533
rect 30424 1481 30427 1533
rect 30369 1469 30427 1481
rect 30369 1417 30372 1469
rect 30424 1417 30427 1469
rect 30369 1405 30427 1417
rect 30369 1353 30372 1405
rect 30424 1353 30427 1405
rect 30369 1341 30427 1353
rect 30369 1289 30372 1341
rect 30424 1289 30427 1341
rect 30369 1277 30427 1289
rect 30369 1225 30372 1277
rect 30424 1225 30427 1277
rect 30369 1213 30427 1225
rect 30369 1161 30372 1213
rect 30424 1161 30427 1213
rect 30369 830 30427 1161
rect 30465 3135 30523 3147
rect 30465 3079 30466 3135
rect 30522 3079 30523 3135
rect 30465 3069 30523 3079
rect 30465 3055 30468 3069
rect 30520 3055 30523 3069
rect 30465 2999 30466 3055
rect 30522 2999 30523 3055
rect 30465 2975 30468 2999
rect 30520 2975 30523 2999
rect 30465 2919 30466 2975
rect 30522 2919 30523 2975
rect 30465 2895 30468 2919
rect 30520 2895 30523 2919
rect 30465 2839 30466 2895
rect 30522 2839 30523 2895
rect 30465 2825 30468 2839
rect 30520 2825 30523 2839
rect 30465 2815 30523 2825
rect 30465 2759 30466 2815
rect 30522 2759 30523 2815
rect 30465 2749 30523 2759
rect 30465 2735 30468 2749
rect 30520 2735 30523 2749
rect 30465 2679 30466 2735
rect 30522 2679 30523 2735
rect 30465 2655 30468 2679
rect 30520 2655 30523 2679
rect 30465 2599 30466 2655
rect 30522 2599 30523 2655
rect 30465 2575 30468 2599
rect 30520 2575 30523 2599
rect 30465 2519 30466 2575
rect 30522 2519 30523 2575
rect 30465 2505 30468 2519
rect 30520 2505 30523 2519
rect 30465 2495 30523 2505
rect 30465 2439 30466 2495
rect 30522 2439 30523 2495
rect 30465 2429 30523 2439
rect 30465 2415 30468 2429
rect 30520 2415 30523 2429
rect 30465 2359 30466 2415
rect 30522 2359 30523 2415
rect 30465 2335 30468 2359
rect 30520 2335 30523 2359
rect 30465 2279 30466 2335
rect 30522 2279 30523 2335
rect 30465 2255 30468 2279
rect 30520 2255 30523 2279
rect 30465 2199 30466 2255
rect 30522 2199 30523 2255
rect 30465 2185 30468 2199
rect 30520 2185 30523 2199
rect 30465 2175 30523 2185
rect 30465 2119 30466 2175
rect 30522 2119 30523 2175
rect 30465 2109 30523 2119
rect 30465 2095 30468 2109
rect 30520 2095 30523 2109
rect 30465 2039 30466 2095
rect 30522 2039 30523 2095
rect 30465 2015 30468 2039
rect 30520 2015 30523 2039
rect 30465 1959 30466 2015
rect 30522 1959 30523 2015
rect 30465 1935 30468 1959
rect 30520 1935 30523 1959
rect 30465 1879 30466 1935
rect 30522 1879 30523 1935
rect 30465 1865 30468 1879
rect 30520 1865 30523 1879
rect 30465 1855 30523 1865
rect 30465 1799 30466 1855
rect 30522 1799 30523 1855
rect 30465 1789 30523 1799
rect 30465 1775 30468 1789
rect 30520 1775 30523 1789
rect 30465 1719 30466 1775
rect 30522 1719 30523 1775
rect 30465 1695 30468 1719
rect 30520 1695 30523 1719
rect 30465 1639 30466 1695
rect 30522 1639 30523 1695
rect 30465 1615 30468 1639
rect 30520 1615 30523 1639
rect 30465 1559 30466 1615
rect 30522 1559 30523 1615
rect 30465 1545 30468 1559
rect 30520 1545 30523 1559
rect 30465 1535 30523 1545
rect 30465 1479 30466 1535
rect 30522 1479 30523 1535
rect 30465 1469 30523 1479
rect 30465 1455 30468 1469
rect 30520 1455 30523 1469
rect 30465 1399 30466 1455
rect 30522 1399 30523 1455
rect 30465 1375 30468 1399
rect 30520 1375 30523 1399
rect 30465 1319 30466 1375
rect 30522 1319 30523 1375
rect 30465 1295 30468 1319
rect 30520 1295 30523 1319
rect 30465 1239 30466 1295
rect 30522 1239 30523 1295
rect 30465 1225 30468 1239
rect 30520 1225 30523 1239
rect 30465 1215 30523 1225
rect 30465 1159 30466 1215
rect 30522 1159 30523 1215
rect 30465 1147 30523 1159
rect 30561 3133 30619 3147
rect 30561 3081 30564 3133
rect 30616 3081 30619 3133
rect 30561 3069 30619 3081
rect 30561 3017 30564 3069
rect 30616 3017 30619 3069
rect 30561 3005 30619 3017
rect 30561 2953 30564 3005
rect 30616 2953 30619 3005
rect 30561 2941 30619 2953
rect 30561 2889 30564 2941
rect 30616 2889 30619 2941
rect 30561 2877 30619 2889
rect 30561 2825 30564 2877
rect 30616 2825 30619 2877
rect 30561 2813 30619 2825
rect 30561 2761 30564 2813
rect 30616 2761 30619 2813
rect 30561 2749 30619 2761
rect 30561 2697 30564 2749
rect 30616 2697 30619 2749
rect 30561 2685 30619 2697
rect 30561 2633 30564 2685
rect 30616 2633 30619 2685
rect 30561 2621 30619 2633
rect 30561 2569 30564 2621
rect 30616 2569 30619 2621
rect 30561 2557 30619 2569
rect 30561 2505 30564 2557
rect 30616 2505 30619 2557
rect 30561 2493 30619 2505
rect 30561 2441 30564 2493
rect 30616 2441 30619 2493
rect 30561 2429 30619 2441
rect 30561 2377 30564 2429
rect 30616 2377 30619 2429
rect 30561 2365 30619 2377
rect 30561 2313 30564 2365
rect 30616 2313 30619 2365
rect 30561 2301 30619 2313
rect 30561 2249 30564 2301
rect 30616 2249 30619 2301
rect 30561 2237 30619 2249
rect 30561 2185 30564 2237
rect 30616 2185 30619 2237
rect 30561 2173 30619 2185
rect 30561 2121 30564 2173
rect 30616 2121 30619 2173
rect 30561 2109 30619 2121
rect 30561 2057 30564 2109
rect 30616 2057 30619 2109
rect 30561 2045 30619 2057
rect 30561 1993 30564 2045
rect 30616 1993 30619 2045
rect 30561 1981 30619 1993
rect 30561 1929 30564 1981
rect 30616 1929 30619 1981
rect 30561 1917 30619 1929
rect 30561 1865 30564 1917
rect 30616 1865 30619 1917
rect 30561 1853 30619 1865
rect 30561 1801 30564 1853
rect 30616 1801 30619 1853
rect 30561 1789 30619 1801
rect 30561 1737 30564 1789
rect 30616 1737 30619 1789
rect 30561 1725 30619 1737
rect 30561 1673 30564 1725
rect 30616 1673 30619 1725
rect 30561 1661 30619 1673
rect 30561 1609 30564 1661
rect 30616 1609 30619 1661
rect 30561 1597 30619 1609
rect 30561 1545 30564 1597
rect 30616 1545 30619 1597
rect 30561 1533 30619 1545
rect 30561 1481 30564 1533
rect 30616 1481 30619 1533
rect 30561 1469 30619 1481
rect 30561 1417 30564 1469
rect 30616 1417 30619 1469
rect 30561 1405 30619 1417
rect 30561 1353 30564 1405
rect 30616 1353 30619 1405
rect 30561 1341 30619 1353
rect 30561 1289 30564 1341
rect 30616 1289 30619 1341
rect 30561 1277 30619 1289
rect 30561 1225 30564 1277
rect 30616 1225 30619 1277
rect 30561 1213 30619 1225
rect 30561 1161 30564 1213
rect 30616 1161 30619 1213
rect 30561 830 30619 1161
rect 30657 3135 30715 3147
rect 30657 3079 30658 3135
rect 30714 3079 30715 3135
rect 30657 3069 30715 3079
rect 30657 3055 30660 3069
rect 30712 3055 30715 3069
rect 30657 2999 30658 3055
rect 30714 2999 30715 3055
rect 30657 2975 30660 2999
rect 30712 2975 30715 2999
rect 30657 2919 30658 2975
rect 30714 2919 30715 2975
rect 30657 2895 30660 2919
rect 30712 2895 30715 2919
rect 30657 2839 30658 2895
rect 30714 2839 30715 2895
rect 30657 2825 30660 2839
rect 30712 2825 30715 2839
rect 30657 2815 30715 2825
rect 30657 2759 30658 2815
rect 30714 2759 30715 2815
rect 30657 2749 30715 2759
rect 30657 2735 30660 2749
rect 30712 2735 30715 2749
rect 30657 2679 30658 2735
rect 30714 2679 30715 2735
rect 30657 2655 30660 2679
rect 30712 2655 30715 2679
rect 30657 2599 30658 2655
rect 30714 2599 30715 2655
rect 30657 2575 30660 2599
rect 30712 2575 30715 2599
rect 30657 2519 30658 2575
rect 30714 2519 30715 2575
rect 30657 2505 30660 2519
rect 30712 2505 30715 2519
rect 30657 2495 30715 2505
rect 30657 2439 30658 2495
rect 30714 2439 30715 2495
rect 30657 2429 30715 2439
rect 30657 2415 30660 2429
rect 30712 2415 30715 2429
rect 30657 2359 30658 2415
rect 30714 2359 30715 2415
rect 30657 2335 30660 2359
rect 30712 2335 30715 2359
rect 30657 2279 30658 2335
rect 30714 2279 30715 2335
rect 30657 2255 30660 2279
rect 30712 2255 30715 2279
rect 30657 2199 30658 2255
rect 30714 2199 30715 2255
rect 30657 2185 30660 2199
rect 30712 2185 30715 2199
rect 30657 2175 30715 2185
rect 30657 2119 30658 2175
rect 30714 2119 30715 2175
rect 30657 2109 30715 2119
rect 30657 2095 30660 2109
rect 30712 2095 30715 2109
rect 30657 2039 30658 2095
rect 30714 2039 30715 2095
rect 30657 2015 30660 2039
rect 30712 2015 30715 2039
rect 30657 1959 30658 2015
rect 30714 1959 30715 2015
rect 30657 1935 30660 1959
rect 30712 1935 30715 1959
rect 30657 1879 30658 1935
rect 30714 1879 30715 1935
rect 30657 1865 30660 1879
rect 30712 1865 30715 1879
rect 30657 1855 30715 1865
rect 30657 1799 30658 1855
rect 30714 1799 30715 1855
rect 30657 1789 30715 1799
rect 30657 1775 30660 1789
rect 30712 1775 30715 1789
rect 30657 1719 30658 1775
rect 30714 1719 30715 1775
rect 30657 1695 30660 1719
rect 30712 1695 30715 1719
rect 30657 1639 30658 1695
rect 30714 1639 30715 1695
rect 30657 1615 30660 1639
rect 30712 1615 30715 1639
rect 30657 1559 30658 1615
rect 30714 1559 30715 1615
rect 30657 1545 30660 1559
rect 30712 1545 30715 1559
rect 30657 1535 30715 1545
rect 30657 1479 30658 1535
rect 30714 1479 30715 1535
rect 30657 1469 30715 1479
rect 30657 1455 30660 1469
rect 30712 1455 30715 1469
rect 30657 1399 30658 1455
rect 30714 1399 30715 1455
rect 30657 1375 30660 1399
rect 30712 1375 30715 1399
rect 30657 1319 30658 1375
rect 30714 1319 30715 1375
rect 30657 1295 30660 1319
rect 30712 1295 30715 1319
rect 30657 1239 30658 1295
rect 30714 1239 30715 1295
rect 30657 1225 30660 1239
rect 30712 1225 30715 1239
rect 30657 1215 30715 1225
rect 30657 1159 30658 1215
rect 30714 1159 30715 1215
rect 30657 1147 30715 1159
rect 30753 3133 30811 3147
rect 30753 3081 30756 3133
rect 30808 3081 30811 3133
rect 30753 3069 30811 3081
rect 30753 3017 30756 3069
rect 30808 3017 30811 3069
rect 30753 3005 30811 3017
rect 30753 2953 30756 3005
rect 30808 2953 30811 3005
rect 30753 2941 30811 2953
rect 30753 2889 30756 2941
rect 30808 2889 30811 2941
rect 30753 2877 30811 2889
rect 30753 2825 30756 2877
rect 30808 2825 30811 2877
rect 30753 2813 30811 2825
rect 30753 2761 30756 2813
rect 30808 2761 30811 2813
rect 30753 2749 30811 2761
rect 30753 2697 30756 2749
rect 30808 2697 30811 2749
rect 30753 2685 30811 2697
rect 30753 2633 30756 2685
rect 30808 2633 30811 2685
rect 30753 2621 30811 2633
rect 30753 2569 30756 2621
rect 30808 2569 30811 2621
rect 30753 2557 30811 2569
rect 30753 2505 30756 2557
rect 30808 2505 30811 2557
rect 30753 2493 30811 2505
rect 30753 2441 30756 2493
rect 30808 2441 30811 2493
rect 30753 2429 30811 2441
rect 30753 2377 30756 2429
rect 30808 2377 30811 2429
rect 30753 2365 30811 2377
rect 30753 2313 30756 2365
rect 30808 2313 30811 2365
rect 30753 2301 30811 2313
rect 30753 2249 30756 2301
rect 30808 2249 30811 2301
rect 30753 2237 30811 2249
rect 30753 2185 30756 2237
rect 30808 2185 30811 2237
rect 30753 2173 30811 2185
rect 30753 2121 30756 2173
rect 30808 2121 30811 2173
rect 30753 2109 30811 2121
rect 30753 2057 30756 2109
rect 30808 2057 30811 2109
rect 30753 2045 30811 2057
rect 30753 1993 30756 2045
rect 30808 1993 30811 2045
rect 30753 1981 30811 1993
rect 30753 1929 30756 1981
rect 30808 1929 30811 1981
rect 30753 1917 30811 1929
rect 30753 1865 30756 1917
rect 30808 1865 30811 1917
rect 30753 1853 30811 1865
rect 30753 1801 30756 1853
rect 30808 1801 30811 1853
rect 30753 1789 30811 1801
rect 30753 1737 30756 1789
rect 30808 1737 30811 1789
rect 30753 1725 30811 1737
rect 30753 1673 30756 1725
rect 30808 1673 30811 1725
rect 30753 1661 30811 1673
rect 30753 1609 30756 1661
rect 30808 1609 30811 1661
rect 30753 1597 30811 1609
rect 30753 1545 30756 1597
rect 30808 1545 30811 1597
rect 30753 1533 30811 1545
rect 30753 1481 30756 1533
rect 30808 1481 30811 1533
rect 30753 1469 30811 1481
rect 30753 1417 30756 1469
rect 30808 1417 30811 1469
rect 30753 1405 30811 1417
rect 30753 1353 30756 1405
rect 30808 1353 30811 1405
rect 30753 1341 30811 1353
rect 30753 1289 30756 1341
rect 30808 1289 30811 1341
rect 30753 1277 30811 1289
rect 30753 1225 30756 1277
rect 30808 1225 30811 1277
rect 30753 1213 30811 1225
rect 30753 1161 30756 1213
rect 30808 1161 30811 1213
rect 30753 830 30811 1161
rect 30849 3135 30907 3147
rect 30849 3079 30850 3135
rect 30906 3079 30907 3135
rect 30849 3069 30907 3079
rect 30849 3055 30852 3069
rect 30904 3055 30907 3069
rect 30849 2999 30850 3055
rect 30906 2999 30907 3055
rect 30849 2975 30852 2999
rect 30904 2975 30907 2999
rect 30849 2919 30850 2975
rect 30906 2919 30907 2975
rect 30849 2895 30852 2919
rect 30904 2895 30907 2919
rect 30849 2839 30850 2895
rect 30906 2839 30907 2895
rect 30849 2825 30852 2839
rect 30904 2825 30907 2839
rect 30849 2815 30907 2825
rect 30849 2759 30850 2815
rect 30906 2759 30907 2815
rect 30849 2749 30907 2759
rect 30849 2735 30852 2749
rect 30904 2735 30907 2749
rect 30849 2679 30850 2735
rect 30906 2679 30907 2735
rect 30849 2655 30852 2679
rect 30904 2655 30907 2679
rect 30849 2599 30850 2655
rect 30906 2599 30907 2655
rect 30849 2575 30852 2599
rect 30904 2575 30907 2599
rect 30849 2519 30850 2575
rect 30906 2519 30907 2575
rect 30849 2505 30852 2519
rect 30904 2505 30907 2519
rect 30849 2495 30907 2505
rect 30849 2439 30850 2495
rect 30906 2439 30907 2495
rect 30849 2429 30907 2439
rect 30849 2415 30852 2429
rect 30904 2415 30907 2429
rect 30849 2359 30850 2415
rect 30906 2359 30907 2415
rect 30849 2335 30852 2359
rect 30904 2335 30907 2359
rect 30849 2279 30850 2335
rect 30906 2279 30907 2335
rect 30849 2255 30852 2279
rect 30904 2255 30907 2279
rect 30849 2199 30850 2255
rect 30906 2199 30907 2255
rect 30849 2185 30852 2199
rect 30904 2185 30907 2199
rect 30849 2175 30907 2185
rect 30849 2119 30850 2175
rect 30906 2119 30907 2175
rect 30849 2109 30907 2119
rect 30849 2095 30852 2109
rect 30904 2095 30907 2109
rect 30849 2039 30850 2095
rect 30906 2039 30907 2095
rect 30849 2015 30852 2039
rect 30904 2015 30907 2039
rect 30849 1959 30850 2015
rect 30906 1959 30907 2015
rect 30849 1935 30852 1959
rect 30904 1935 30907 1959
rect 30849 1879 30850 1935
rect 30906 1879 30907 1935
rect 30849 1865 30852 1879
rect 30904 1865 30907 1879
rect 30849 1855 30907 1865
rect 30849 1799 30850 1855
rect 30906 1799 30907 1855
rect 30849 1789 30907 1799
rect 30849 1775 30852 1789
rect 30904 1775 30907 1789
rect 30849 1719 30850 1775
rect 30906 1719 30907 1775
rect 30849 1695 30852 1719
rect 30904 1695 30907 1719
rect 30849 1639 30850 1695
rect 30906 1639 30907 1695
rect 30849 1615 30852 1639
rect 30904 1615 30907 1639
rect 30849 1559 30850 1615
rect 30906 1559 30907 1615
rect 30849 1545 30852 1559
rect 30904 1545 30907 1559
rect 30849 1535 30907 1545
rect 30849 1479 30850 1535
rect 30906 1479 30907 1535
rect 30849 1469 30907 1479
rect 30849 1455 30852 1469
rect 30904 1455 30907 1469
rect 30849 1399 30850 1455
rect 30906 1399 30907 1455
rect 30849 1375 30852 1399
rect 30904 1375 30907 1399
rect 30849 1319 30850 1375
rect 30906 1319 30907 1375
rect 30849 1295 30852 1319
rect 30904 1295 30907 1319
rect 30849 1239 30850 1295
rect 30906 1239 30907 1295
rect 30849 1225 30852 1239
rect 30904 1225 30907 1239
rect 30849 1215 30907 1225
rect 30849 1159 30850 1215
rect 30906 1159 30907 1215
rect 30849 1147 30907 1159
rect 30945 3133 31003 3147
rect 30945 3081 30948 3133
rect 31000 3081 31003 3133
rect 30945 3069 31003 3081
rect 30945 3017 30948 3069
rect 31000 3017 31003 3069
rect 30945 3005 31003 3017
rect 30945 2953 30948 3005
rect 31000 2953 31003 3005
rect 30945 2941 31003 2953
rect 30945 2889 30948 2941
rect 31000 2889 31003 2941
rect 30945 2877 31003 2889
rect 30945 2825 30948 2877
rect 31000 2825 31003 2877
rect 30945 2813 31003 2825
rect 30945 2761 30948 2813
rect 31000 2761 31003 2813
rect 30945 2749 31003 2761
rect 30945 2697 30948 2749
rect 31000 2697 31003 2749
rect 30945 2685 31003 2697
rect 30945 2633 30948 2685
rect 31000 2633 31003 2685
rect 30945 2621 31003 2633
rect 30945 2569 30948 2621
rect 31000 2569 31003 2621
rect 30945 2557 31003 2569
rect 30945 2505 30948 2557
rect 31000 2505 31003 2557
rect 30945 2493 31003 2505
rect 30945 2441 30948 2493
rect 31000 2441 31003 2493
rect 30945 2429 31003 2441
rect 30945 2377 30948 2429
rect 31000 2377 31003 2429
rect 30945 2365 31003 2377
rect 30945 2313 30948 2365
rect 31000 2313 31003 2365
rect 30945 2301 31003 2313
rect 30945 2249 30948 2301
rect 31000 2249 31003 2301
rect 30945 2237 31003 2249
rect 30945 2185 30948 2237
rect 31000 2185 31003 2237
rect 30945 2173 31003 2185
rect 30945 2121 30948 2173
rect 31000 2121 31003 2173
rect 30945 2109 31003 2121
rect 30945 2057 30948 2109
rect 31000 2057 31003 2109
rect 30945 2045 31003 2057
rect 30945 1993 30948 2045
rect 31000 1993 31003 2045
rect 30945 1981 31003 1993
rect 30945 1929 30948 1981
rect 31000 1929 31003 1981
rect 30945 1917 31003 1929
rect 30945 1865 30948 1917
rect 31000 1865 31003 1917
rect 30945 1853 31003 1865
rect 30945 1801 30948 1853
rect 31000 1801 31003 1853
rect 30945 1789 31003 1801
rect 30945 1737 30948 1789
rect 31000 1737 31003 1789
rect 30945 1725 31003 1737
rect 30945 1673 30948 1725
rect 31000 1673 31003 1725
rect 30945 1661 31003 1673
rect 30945 1609 30948 1661
rect 31000 1609 31003 1661
rect 30945 1597 31003 1609
rect 30945 1545 30948 1597
rect 31000 1545 31003 1597
rect 30945 1533 31003 1545
rect 30945 1481 30948 1533
rect 31000 1481 31003 1533
rect 30945 1469 31003 1481
rect 30945 1417 30948 1469
rect 31000 1417 31003 1469
rect 30945 1405 31003 1417
rect 30945 1353 30948 1405
rect 31000 1353 31003 1405
rect 30945 1341 31003 1353
rect 30945 1289 30948 1341
rect 31000 1289 31003 1341
rect 30945 1277 31003 1289
rect 30945 1225 30948 1277
rect 31000 1225 31003 1277
rect 30945 1213 31003 1225
rect 30945 1161 30948 1213
rect 31000 1161 31003 1213
rect 30945 830 31003 1161
rect 31041 3135 31099 3147
rect 31041 3079 31042 3135
rect 31098 3079 31099 3135
rect 31041 3069 31099 3079
rect 31041 3055 31044 3069
rect 31096 3055 31099 3069
rect 31041 2999 31042 3055
rect 31098 2999 31099 3055
rect 31041 2975 31044 2999
rect 31096 2975 31099 2999
rect 31041 2919 31042 2975
rect 31098 2919 31099 2975
rect 31041 2895 31044 2919
rect 31096 2895 31099 2919
rect 31041 2839 31042 2895
rect 31098 2839 31099 2895
rect 31041 2825 31044 2839
rect 31096 2825 31099 2839
rect 31041 2815 31099 2825
rect 31041 2759 31042 2815
rect 31098 2759 31099 2815
rect 31041 2749 31099 2759
rect 31041 2735 31044 2749
rect 31096 2735 31099 2749
rect 31041 2679 31042 2735
rect 31098 2679 31099 2735
rect 31041 2655 31044 2679
rect 31096 2655 31099 2679
rect 31041 2599 31042 2655
rect 31098 2599 31099 2655
rect 31041 2575 31044 2599
rect 31096 2575 31099 2599
rect 31041 2519 31042 2575
rect 31098 2519 31099 2575
rect 31041 2505 31044 2519
rect 31096 2505 31099 2519
rect 31041 2495 31099 2505
rect 31041 2439 31042 2495
rect 31098 2439 31099 2495
rect 31041 2429 31099 2439
rect 31041 2415 31044 2429
rect 31096 2415 31099 2429
rect 31041 2359 31042 2415
rect 31098 2359 31099 2415
rect 31041 2335 31044 2359
rect 31096 2335 31099 2359
rect 31041 2279 31042 2335
rect 31098 2279 31099 2335
rect 31041 2255 31044 2279
rect 31096 2255 31099 2279
rect 31041 2199 31042 2255
rect 31098 2199 31099 2255
rect 31041 2185 31044 2199
rect 31096 2185 31099 2199
rect 31041 2175 31099 2185
rect 31041 2119 31042 2175
rect 31098 2119 31099 2175
rect 31041 2109 31099 2119
rect 31041 2095 31044 2109
rect 31096 2095 31099 2109
rect 31041 2039 31042 2095
rect 31098 2039 31099 2095
rect 31041 2015 31044 2039
rect 31096 2015 31099 2039
rect 31041 1959 31042 2015
rect 31098 1959 31099 2015
rect 31041 1935 31044 1959
rect 31096 1935 31099 1959
rect 31041 1879 31042 1935
rect 31098 1879 31099 1935
rect 31041 1865 31044 1879
rect 31096 1865 31099 1879
rect 31041 1855 31099 1865
rect 31041 1799 31042 1855
rect 31098 1799 31099 1855
rect 31041 1789 31099 1799
rect 31041 1775 31044 1789
rect 31096 1775 31099 1789
rect 31041 1719 31042 1775
rect 31098 1719 31099 1775
rect 31041 1695 31044 1719
rect 31096 1695 31099 1719
rect 31041 1639 31042 1695
rect 31098 1639 31099 1695
rect 31041 1615 31044 1639
rect 31096 1615 31099 1639
rect 31041 1559 31042 1615
rect 31098 1559 31099 1615
rect 31041 1545 31044 1559
rect 31096 1545 31099 1559
rect 31041 1535 31099 1545
rect 31041 1479 31042 1535
rect 31098 1479 31099 1535
rect 31041 1469 31099 1479
rect 31041 1455 31044 1469
rect 31096 1455 31099 1469
rect 31041 1399 31042 1455
rect 31098 1399 31099 1455
rect 31041 1375 31044 1399
rect 31096 1375 31099 1399
rect 31041 1319 31042 1375
rect 31098 1319 31099 1375
rect 31041 1295 31044 1319
rect 31096 1295 31099 1319
rect 31041 1239 31042 1295
rect 31098 1239 31099 1295
rect 31041 1225 31044 1239
rect 31096 1225 31099 1239
rect 31041 1215 31099 1225
rect 31041 1159 31042 1215
rect 31098 1159 31099 1215
rect 31041 1147 31099 1159
rect 31137 3133 31195 3147
rect 31137 3081 31140 3133
rect 31192 3081 31195 3133
rect 31137 3069 31195 3081
rect 31137 3017 31140 3069
rect 31192 3017 31195 3069
rect 31137 3005 31195 3017
rect 31137 2953 31140 3005
rect 31192 2953 31195 3005
rect 31137 2941 31195 2953
rect 31137 2889 31140 2941
rect 31192 2889 31195 2941
rect 31137 2877 31195 2889
rect 31137 2825 31140 2877
rect 31192 2825 31195 2877
rect 31137 2813 31195 2825
rect 31137 2761 31140 2813
rect 31192 2761 31195 2813
rect 31137 2749 31195 2761
rect 31137 2697 31140 2749
rect 31192 2697 31195 2749
rect 31137 2685 31195 2697
rect 31137 2633 31140 2685
rect 31192 2633 31195 2685
rect 31137 2621 31195 2633
rect 31137 2569 31140 2621
rect 31192 2569 31195 2621
rect 31137 2557 31195 2569
rect 31137 2505 31140 2557
rect 31192 2505 31195 2557
rect 31137 2493 31195 2505
rect 31137 2441 31140 2493
rect 31192 2441 31195 2493
rect 31137 2429 31195 2441
rect 31137 2377 31140 2429
rect 31192 2377 31195 2429
rect 31137 2365 31195 2377
rect 31137 2313 31140 2365
rect 31192 2313 31195 2365
rect 31137 2301 31195 2313
rect 31137 2249 31140 2301
rect 31192 2249 31195 2301
rect 31137 2237 31195 2249
rect 31137 2185 31140 2237
rect 31192 2185 31195 2237
rect 31137 2173 31195 2185
rect 31137 2121 31140 2173
rect 31192 2121 31195 2173
rect 31137 2109 31195 2121
rect 31137 2057 31140 2109
rect 31192 2057 31195 2109
rect 31137 2045 31195 2057
rect 31137 1993 31140 2045
rect 31192 1993 31195 2045
rect 31137 1981 31195 1993
rect 31137 1929 31140 1981
rect 31192 1929 31195 1981
rect 31137 1917 31195 1929
rect 31137 1865 31140 1917
rect 31192 1865 31195 1917
rect 31137 1853 31195 1865
rect 31137 1801 31140 1853
rect 31192 1801 31195 1853
rect 31137 1789 31195 1801
rect 31137 1737 31140 1789
rect 31192 1737 31195 1789
rect 31137 1725 31195 1737
rect 31137 1673 31140 1725
rect 31192 1673 31195 1725
rect 31137 1661 31195 1673
rect 31137 1609 31140 1661
rect 31192 1609 31195 1661
rect 31137 1597 31195 1609
rect 31137 1545 31140 1597
rect 31192 1545 31195 1597
rect 31137 1533 31195 1545
rect 31137 1481 31140 1533
rect 31192 1481 31195 1533
rect 31137 1469 31195 1481
rect 31137 1417 31140 1469
rect 31192 1417 31195 1469
rect 31137 1405 31195 1417
rect 31137 1353 31140 1405
rect 31192 1353 31195 1405
rect 31137 1341 31195 1353
rect 31137 1289 31140 1341
rect 31192 1289 31195 1341
rect 31137 1277 31195 1289
rect 31137 1225 31140 1277
rect 31192 1225 31195 1277
rect 31137 1213 31195 1225
rect 31137 1161 31140 1213
rect 31192 1161 31195 1213
rect 31137 830 31195 1161
rect 31233 3135 31291 3147
rect 31233 3079 31234 3135
rect 31290 3079 31291 3135
rect 31233 3069 31291 3079
rect 31233 3055 31236 3069
rect 31288 3055 31291 3069
rect 31233 2999 31234 3055
rect 31290 2999 31291 3055
rect 31233 2975 31236 2999
rect 31288 2975 31291 2999
rect 31233 2919 31234 2975
rect 31290 2919 31291 2975
rect 31233 2895 31236 2919
rect 31288 2895 31291 2919
rect 31233 2839 31234 2895
rect 31290 2839 31291 2895
rect 31233 2825 31236 2839
rect 31288 2825 31291 2839
rect 31233 2815 31291 2825
rect 31233 2759 31234 2815
rect 31290 2759 31291 2815
rect 31233 2749 31291 2759
rect 31233 2735 31236 2749
rect 31288 2735 31291 2749
rect 31233 2679 31234 2735
rect 31290 2679 31291 2735
rect 31233 2655 31236 2679
rect 31288 2655 31291 2679
rect 31233 2599 31234 2655
rect 31290 2599 31291 2655
rect 31233 2575 31236 2599
rect 31288 2575 31291 2599
rect 31233 2519 31234 2575
rect 31290 2519 31291 2575
rect 31233 2505 31236 2519
rect 31288 2505 31291 2519
rect 31233 2495 31291 2505
rect 31233 2439 31234 2495
rect 31290 2439 31291 2495
rect 31233 2429 31291 2439
rect 31233 2415 31236 2429
rect 31288 2415 31291 2429
rect 31233 2359 31234 2415
rect 31290 2359 31291 2415
rect 31233 2335 31236 2359
rect 31288 2335 31291 2359
rect 31233 2279 31234 2335
rect 31290 2279 31291 2335
rect 31233 2255 31236 2279
rect 31288 2255 31291 2279
rect 31233 2199 31234 2255
rect 31290 2199 31291 2255
rect 31233 2185 31236 2199
rect 31288 2185 31291 2199
rect 31233 2175 31291 2185
rect 31233 2119 31234 2175
rect 31290 2119 31291 2175
rect 31233 2109 31291 2119
rect 31233 2095 31236 2109
rect 31288 2095 31291 2109
rect 31233 2039 31234 2095
rect 31290 2039 31291 2095
rect 31233 2015 31236 2039
rect 31288 2015 31291 2039
rect 31233 1959 31234 2015
rect 31290 1959 31291 2015
rect 31233 1935 31236 1959
rect 31288 1935 31291 1959
rect 31233 1879 31234 1935
rect 31290 1879 31291 1935
rect 31233 1865 31236 1879
rect 31288 1865 31291 1879
rect 31233 1855 31291 1865
rect 31233 1799 31234 1855
rect 31290 1799 31291 1855
rect 31233 1789 31291 1799
rect 31233 1775 31236 1789
rect 31288 1775 31291 1789
rect 31233 1719 31234 1775
rect 31290 1719 31291 1775
rect 31233 1695 31236 1719
rect 31288 1695 31291 1719
rect 31233 1639 31234 1695
rect 31290 1639 31291 1695
rect 31233 1615 31236 1639
rect 31288 1615 31291 1639
rect 31233 1559 31234 1615
rect 31290 1559 31291 1615
rect 31233 1545 31236 1559
rect 31288 1545 31291 1559
rect 31233 1535 31291 1545
rect 31233 1479 31234 1535
rect 31290 1479 31291 1535
rect 31233 1469 31291 1479
rect 31233 1455 31236 1469
rect 31288 1455 31291 1469
rect 31233 1399 31234 1455
rect 31290 1399 31291 1455
rect 31233 1375 31236 1399
rect 31288 1375 31291 1399
rect 31233 1319 31234 1375
rect 31290 1319 31291 1375
rect 31233 1295 31236 1319
rect 31288 1295 31291 1319
rect 31233 1239 31234 1295
rect 31290 1239 31291 1295
rect 31233 1225 31236 1239
rect 31288 1225 31291 1239
rect 31233 1215 31291 1225
rect 31233 1159 31234 1215
rect 31290 1159 31291 1215
rect 31233 1147 31291 1159
rect 31329 3133 31387 3147
rect 31329 3081 31332 3133
rect 31384 3081 31387 3133
rect 31329 3069 31387 3081
rect 31329 3017 31332 3069
rect 31384 3017 31387 3069
rect 31329 3005 31387 3017
rect 31329 2953 31332 3005
rect 31384 2953 31387 3005
rect 31329 2941 31387 2953
rect 31329 2889 31332 2941
rect 31384 2889 31387 2941
rect 31329 2877 31387 2889
rect 31329 2825 31332 2877
rect 31384 2825 31387 2877
rect 31329 2813 31387 2825
rect 31329 2761 31332 2813
rect 31384 2761 31387 2813
rect 31329 2749 31387 2761
rect 31329 2697 31332 2749
rect 31384 2697 31387 2749
rect 31329 2685 31387 2697
rect 31329 2633 31332 2685
rect 31384 2633 31387 2685
rect 31329 2621 31387 2633
rect 31329 2569 31332 2621
rect 31384 2569 31387 2621
rect 31329 2557 31387 2569
rect 31329 2505 31332 2557
rect 31384 2505 31387 2557
rect 31329 2493 31387 2505
rect 31329 2441 31332 2493
rect 31384 2441 31387 2493
rect 31329 2429 31387 2441
rect 31329 2377 31332 2429
rect 31384 2377 31387 2429
rect 31329 2365 31387 2377
rect 31329 2313 31332 2365
rect 31384 2313 31387 2365
rect 31329 2301 31387 2313
rect 31329 2249 31332 2301
rect 31384 2249 31387 2301
rect 31329 2237 31387 2249
rect 31329 2185 31332 2237
rect 31384 2185 31387 2237
rect 31329 2173 31387 2185
rect 31329 2121 31332 2173
rect 31384 2121 31387 2173
rect 31329 2109 31387 2121
rect 31329 2057 31332 2109
rect 31384 2057 31387 2109
rect 31329 2045 31387 2057
rect 31329 1993 31332 2045
rect 31384 1993 31387 2045
rect 31329 1981 31387 1993
rect 31329 1929 31332 1981
rect 31384 1929 31387 1981
rect 31329 1917 31387 1929
rect 31329 1865 31332 1917
rect 31384 1865 31387 1917
rect 31329 1853 31387 1865
rect 31329 1801 31332 1853
rect 31384 1801 31387 1853
rect 31329 1789 31387 1801
rect 31329 1737 31332 1789
rect 31384 1737 31387 1789
rect 31329 1725 31387 1737
rect 31329 1673 31332 1725
rect 31384 1673 31387 1725
rect 31329 1661 31387 1673
rect 31329 1609 31332 1661
rect 31384 1609 31387 1661
rect 31329 1597 31387 1609
rect 31329 1545 31332 1597
rect 31384 1545 31387 1597
rect 31329 1533 31387 1545
rect 31329 1481 31332 1533
rect 31384 1481 31387 1533
rect 31329 1469 31387 1481
rect 31329 1417 31332 1469
rect 31384 1417 31387 1469
rect 31329 1405 31387 1417
rect 31329 1353 31332 1405
rect 31384 1353 31387 1405
rect 31329 1341 31387 1353
rect 31329 1289 31332 1341
rect 31384 1289 31387 1341
rect 31329 1277 31387 1289
rect 31329 1225 31332 1277
rect 31384 1225 31387 1277
rect 31329 1213 31387 1225
rect 31329 1161 31332 1213
rect 31384 1161 31387 1213
rect 31329 830 31387 1161
rect 31425 3135 31483 3147
rect 31425 3079 31426 3135
rect 31482 3079 31483 3135
rect 31425 3069 31483 3079
rect 31425 3055 31428 3069
rect 31480 3055 31483 3069
rect 31425 2999 31426 3055
rect 31482 2999 31483 3055
rect 31425 2975 31428 2999
rect 31480 2975 31483 2999
rect 31425 2919 31426 2975
rect 31482 2919 31483 2975
rect 31425 2895 31428 2919
rect 31480 2895 31483 2919
rect 31425 2839 31426 2895
rect 31482 2839 31483 2895
rect 31425 2825 31428 2839
rect 31480 2825 31483 2839
rect 31425 2815 31483 2825
rect 31425 2759 31426 2815
rect 31482 2759 31483 2815
rect 31425 2749 31483 2759
rect 31425 2735 31428 2749
rect 31480 2735 31483 2749
rect 31425 2679 31426 2735
rect 31482 2679 31483 2735
rect 31425 2655 31428 2679
rect 31480 2655 31483 2679
rect 31425 2599 31426 2655
rect 31482 2599 31483 2655
rect 31425 2575 31428 2599
rect 31480 2575 31483 2599
rect 31425 2519 31426 2575
rect 31482 2519 31483 2575
rect 31425 2505 31428 2519
rect 31480 2505 31483 2519
rect 31425 2495 31483 2505
rect 31425 2439 31426 2495
rect 31482 2439 31483 2495
rect 31425 2429 31483 2439
rect 31425 2415 31428 2429
rect 31480 2415 31483 2429
rect 31425 2359 31426 2415
rect 31482 2359 31483 2415
rect 31425 2335 31428 2359
rect 31480 2335 31483 2359
rect 31425 2279 31426 2335
rect 31482 2279 31483 2335
rect 31425 2255 31428 2279
rect 31480 2255 31483 2279
rect 31425 2199 31426 2255
rect 31482 2199 31483 2255
rect 31425 2185 31428 2199
rect 31480 2185 31483 2199
rect 31425 2175 31483 2185
rect 31425 2119 31426 2175
rect 31482 2119 31483 2175
rect 31425 2109 31483 2119
rect 31425 2095 31428 2109
rect 31480 2095 31483 2109
rect 31425 2039 31426 2095
rect 31482 2039 31483 2095
rect 31425 2015 31428 2039
rect 31480 2015 31483 2039
rect 31425 1959 31426 2015
rect 31482 1959 31483 2015
rect 31425 1935 31428 1959
rect 31480 1935 31483 1959
rect 31425 1879 31426 1935
rect 31482 1879 31483 1935
rect 31425 1865 31428 1879
rect 31480 1865 31483 1879
rect 31425 1855 31483 1865
rect 31425 1799 31426 1855
rect 31482 1799 31483 1855
rect 31425 1789 31483 1799
rect 31425 1775 31428 1789
rect 31480 1775 31483 1789
rect 31425 1719 31426 1775
rect 31482 1719 31483 1775
rect 31425 1695 31428 1719
rect 31480 1695 31483 1719
rect 31425 1639 31426 1695
rect 31482 1639 31483 1695
rect 31425 1615 31428 1639
rect 31480 1615 31483 1639
rect 31425 1559 31426 1615
rect 31482 1559 31483 1615
rect 31425 1545 31428 1559
rect 31480 1545 31483 1559
rect 31425 1535 31483 1545
rect 31425 1479 31426 1535
rect 31482 1479 31483 1535
rect 31425 1469 31483 1479
rect 31425 1455 31428 1469
rect 31480 1455 31483 1469
rect 31425 1399 31426 1455
rect 31482 1399 31483 1455
rect 31425 1375 31428 1399
rect 31480 1375 31483 1399
rect 31425 1319 31426 1375
rect 31482 1319 31483 1375
rect 31425 1295 31428 1319
rect 31480 1295 31483 1319
rect 31425 1239 31426 1295
rect 31482 1239 31483 1295
rect 31425 1225 31428 1239
rect 31480 1225 31483 1239
rect 31425 1215 31483 1225
rect 31425 1159 31426 1215
rect 31482 1159 31483 1215
rect 31425 1147 31483 1159
rect 31521 3133 31579 3147
rect 31521 3081 31524 3133
rect 31576 3081 31579 3133
rect 31521 3069 31579 3081
rect 31521 3017 31524 3069
rect 31576 3017 31579 3069
rect 31521 3005 31579 3017
rect 31521 2953 31524 3005
rect 31576 2953 31579 3005
rect 31521 2941 31579 2953
rect 31521 2889 31524 2941
rect 31576 2889 31579 2941
rect 31521 2877 31579 2889
rect 31521 2825 31524 2877
rect 31576 2825 31579 2877
rect 31521 2813 31579 2825
rect 31521 2761 31524 2813
rect 31576 2761 31579 2813
rect 31521 2749 31579 2761
rect 31521 2697 31524 2749
rect 31576 2697 31579 2749
rect 31521 2685 31579 2697
rect 31521 2633 31524 2685
rect 31576 2633 31579 2685
rect 31521 2621 31579 2633
rect 31521 2569 31524 2621
rect 31576 2569 31579 2621
rect 31521 2557 31579 2569
rect 31521 2505 31524 2557
rect 31576 2505 31579 2557
rect 31521 2493 31579 2505
rect 31521 2441 31524 2493
rect 31576 2441 31579 2493
rect 31521 2429 31579 2441
rect 31521 2377 31524 2429
rect 31576 2377 31579 2429
rect 31521 2365 31579 2377
rect 31521 2313 31524 2365
rect 31576 2313 31579 2365
rect 31521 2301 31579 2313
rect 31521 2249 31524 2301
rect 31576 2249 31579 2301
rect 31521 2237 31579 2249
rect 31521 2185 31524 2237
rect 31576 2185 31579 2237
rect 31521 2173 31579 2185
rect 31521 2121 31524 2173
rect 31576 2121 31579 2173
rect 31521 2109 31579 2121
rect 31521 2057 31524 2109
rect 31576 2057 31579 2109
rect 31521 2045 31579 2057
rect 31521 1993 31524 2045
rect 31576 1993 31579 2045
rect 31521 1981 31579 1993
rect 31521 1929 31524 1981
rect 31576 1929 31579 1981
rect 31521 1917 31579 1929
rect 31521 1865 31524 1917
rect 31576 1865 31579 1917
rect 31521 1853 31579 1865
rect 31521 1801 31524 1853
rect 31576 1801 31579 1853
rect 31521 1789 31579 1801
rect 31521 1737 31524 1789
rect 31576 1737 31579 1789
rect 31521 1725 31579 1737
rect 31521 1673 31524 1725
rect 31576 1673 31579 1725
rect 31521 1661 31579 1673
rect 31521 1609 31524 1661
rect 31576 1609 31579 1661
rect 31521 1597 31579 1609
rect 31521 1545 31524 1597
rect 31576 1545 31579 1597
rect 31521 1533 31579 1545
rect 31521 1481 31524 1533
rect 31576 1481 31579 1533
rect 31521 1469 31579 1481
rect 31521 1417 31524 1469
rect 31576 1417 31579 1469
rect 31521 1405 31579 1417
rect 31521 1353 31524 1405
rect 31576 1353 31579 1405
rect 31521 1341 31579 1353
rect 31521 1289 31524 1341
rect 31576 1289 31579 1341
rect 31521 1277 31579 1289
rect 31521 1225 31524 1277
rect 31576 1225 31579 1277
rect 31521 1213 31579 1225
rect 31521 1161 31524 1213
rect 31576 1161 31579 1213
rect 31521 830 31579 1161
rect 31617 3135 31675 3147
rect 31617 3079 31618 3135
rect 31674 3079 31675 3135
rect 31617 3069 31675 3079
rect 31617 3055 31620 3069
rect 31672 3055 31675 3069
rect 31617 2999 31618 3055
rect 31674 2999 31675 3055
rect 31617 2975 31620 2999
rect 31672 2975 31675 2999
rect 31617 2919 31618 2975
rect 31674 2919 31675 2975
rect 31617 2895 31620 2919
rect 31672 2895 31675 2919
rect 31617 2839 31618 2895
rect 31674 2839 31675 2895
rect 31617 2825 31620 2839
rect 31672 2825 31675 2839
rect 31617 2815 31675 2825
rect 31617 2759 31618 2815
rect 31674 2759 31675 2815
rect 31617 2749 31675 2759
rect 31617 2735 31620 2749
rect 31672 2735 31675 2749
rect 31617 2679 31618 2735
rect 31674 2679 31675 2735
rect 31617 2655 31620 2679
rect 31672 2655 31675 2679
rect 31617 2599 31618 2655
rect 31674 2599 31675 2655
rect 31617 2575 31620 2599
rect 31672 2575 31675 2599
rect 31617 2519 31618 2575
rect 31674 2519 31675 2575
rect 31617 2505 31620 2519
rect 31672 2505 31675 2519
rect 31617 2495 31675 2505
rect 31617 2439 31618 2495
rect 31674 2439 31675 2495
rect 31617 2429 31675 2439
rect 31617 2415 31620 2429
rect 31672 2415 31675 2429
rect 31617 2359 31618 2415
rect 31674 2359 31675 2415
rect 31617 2335 31620 2359
rect 31672 2335 31675 2359
rect 31617 2279 31618 2335
rect 31674 2279 31675 2335
rect 31617 2255 31620 2279
rect 31672 2255 31675 2279
rect 31617 2199 31618 2255
rect 31674 2199 31675 2255
rect 31617 2185 31620 2199
rect 31672 2185 31675 2199
rect 31617 2175 31675 2185
rect 31617 2119 31618 2175
rect 31674 2119 31675 2175
rect 31617 2109 31675 2119
rect 31617 2095 31620 2109
rect 31672 2095 31675 2109
rect 31617 2039 31618 2095
rect 31674 2039 31675 2095
rect 31617 2015 31620 2039
rect 31672 2015 31675 2039
rect 31617 1959 31618 2015
rect 31674 1959 31675 2015
rect 31617 1935 31620 1959
rect 31672 1935 31675 1959
rect 31617 1879 31618 1935
rect 31674 1879 31675 1935
rect 31617 1865 31620 1879
rect 31672 1865 31675 1879
rect 31617 1855 31675 1865
rect 31617 1799 31618 1855
rect 31674 1799 31675 1855
rect 31617 1789 31675 1799
rect 31617 1775 31620 1789
rect 31672 1775 31675 1789
rect 31617 1719 31618 1775
rect 31674 1719 31675 1775
rect 31617 1695 31620 1719
rect 31672 1695 31675 1719
rect 31617 1639 31618 1695
rect 31674 1639 31675 1695
rect 31617 1615 31620 1639
rect 31672 1615 31675 1639
rect 31617 1559 31618 1615
rect 31674 1559 31675 1615
rect 31617 1545 31620 1559
rect 31672 1545 31675 1559
rect 31617 1535 31675 1545
rect 31617 1479 31618 1535
rect 31674 1479 31675 1535
rect 31617 1469 31675 1479
rect 31617 1455 31620 1469
rect 31672 1455 31675 1469
rect 31617 1399 31618 1455
rect 31674 1399 31675 1455
rect 31617 1375 31620 1399
rect 31672 1375 31675 1399
rect 31617 1319 31618 1375
rect 31674 1319 31675 1375
rect 31617 1295 31620 1319
rect 31672 1295 31675 1319
rect 31617 1239 31618 1295
rect 31674 1239 31675 1295
rect 31617 1225 31620 1239
rect 31672 1225 31675 1239
rect 31617 1215 31675 1225
rect 31617 1159 31618 1215
rect 31674 1159 31675 1215
rect 31617 1147 31675 1159
rect 31713 3133 31771 3147
rect 31713 3081 31716 3133
rect 31768 3081 31771 3133
rect 31713 3069 31771 3081
rect 31713 3017 31716 3069
rect 31768 3017 31771 3069
rect 31713 3005 31771 3017
rect 31713 2953 31716 3005
rect 31768 2953 31771 3005
rect 31713 2941 31771 2953
rect 31713 2889 31716 2941
rect 31768 2889 31771 2941
rect 31713 2877 31771 2889
rect 31713 2825 31716 2877
rect 31768 2825 31771 2877
rect 31713 2813 31771 2825
rect 31713 2761 31716 2813
rect 31768 2761 31771 2813
rect 31713 2749 31771 2761
rect 31713 2697 31716 2749
rect 31768 2697 31771 2749
rect 31713 2685 31771 2697
rect 31713 2633 31716 2685
rect 31768 2633 31771 2685
rect 31713 2621 31771 2633
rect 31713 2569 31716 2621
rect 31768 2569 31771 2621
rect 31713 2557 31771 2569
rect 31713 2505 31716 2557
rect 31768 2505 31771 2557
rect 31713 2493 31771 2505
rect 31713 2441 31716 2493
rect 31768 2441 31771 2493
rect 31713 2429 31771 2441
rect 31713 2377 31716 2429
rect 31768 2377 31771 2429
rect 31713 2365 31771 2377
rect 31713 2313 31716 2365
rect 31768 2313 31771 2365
rect 31713 2301 31771 2313
rect 31713 2249 31716 2301
rect 31768 2249 31771 2301
rect 31713 2237 31771 2249
rect 31713 2185 31716 2237
rect 31768 2185 31771 2237
rect 31713 2173 31771 2185
rect 31713 2121 31716 2173
rect 31768 2121 31771 2173
rect 31713 2109 31771 2121
rect 31713 2057 31716 2109
rect 31768 2057 31771 2109
rect 31713 2045 31771 2057
rect 31713 1993 31716 2045
rect 31768 1993 31771 2045
rect 31713 1981 31771 1993
rect 31713 1929 31716 1981
rect 31768 1929 31771 1981
rect 31713 1917 31771 1929
rect 31713 1865 31716 1917
rect 31768 1865 31771 1917
rect 31713 1853 31771 1865
rect 31713 1801 31716 1853
rect 31768 1801 31771 1853
rect 31713 1789 31771 1801
rect 31713 1737 31716 1789
rect 31768 1737 31771 1789
rect 31713 1725 31771 1737
rect 31713 1673 31716 1725
rect 31768 1673 31771 1725
rect 31713 1661 31771 1673
rect 31713 1609 31716 1661
rect 31768 1609 31771 1661
rect 31713 1597 31771 1609
rect 31713 1545 31716 1597
rect 31768 1545 31771 1597
rect 31713 1533 31771 1545
rect 31713 1481 31716 1533
rect 31768 1481 31771 1533
rect 31713 1469 31771 1481
rect 31713 1417 31716 1469
rect 31768 1417 31771 1469
rect 31713 1405 31771 1417
rect 31713 1353 31716 1405
rect 31768 1353 31771 1405
rect 31713 1341 31771 1353
rect 31713 1289 31716 1341
rect 31768 1289 31771 1341
rect 31713 1277 31771 1289
rect 31713 1225 31716 1277
rect 31768 1225 31771 1277
rect 31713 1213 31771 1225
rect 31713 1161 31716 1213
rect 31768 1161 31771 1213
rect 31713 830 31771 1161
rect 31809 3135 31867 3147
rect 31809 3079 31810 3135
rect 31866 3079 31867 3135
rect 31809 3069 31867 3079
rect 31809 3055 31812 3069
rect 31864 3055 31867 3069
rect 31809 2999 31810 3055
rect 31866 2999 31867 3055
rect 31809 2975 31812 2999
rect 31864 2975 31867 2999
rect 31809 2919 31810 2975
rect 31866 2919 31867 2975
rect 31809 2895 31812 2919
rect 31864 2895 31867 2919
rect 31809 2839 31810 2895
rect 31866 2839 31867 2895
rect 31809 2825 31812 2839
rect 31864 2825 31867 2839
rect 31809 2815 31867 2825
rect 31809 2759 31810 2815
rect 31866 2759 31867 2815
rect 31809 2749 31867 2759
rect 31809 2735 31812 2749
rect 31864 2735 31867 2749
rect 31809 2679 31810 2735
rect 31866 2679 31867 2735
rect 31809 2655 31812 2679
rect 31864 2655 31867 2679
rect 31809 2599 31810 2655
rect 31866 2599 31867 2655
rect 31809 2575 31812 2599
rect 31864 2575 31867 2599
rect 31809 2519 31810 2575
rect 31866 2519 31867 2575
rect 31809 2505 31812 2519
rect 31864 2505 31867 2519
rect 31809 2495 31867 2505
rect 31809 2439 31810 2495
rect 31866 2439 31867 2495
rect 31809 2429 31867 2439
rect 31809 2415 31812 2429
rect 31864 2415 31867 2429
rect 31809 2359 31810 2415
rect 31866 2359 31867 2415
rect 31809 2335 31812 2359
rect 31864 2335 31867 2359
rect 31809 2279 31810 2335
rect 31866 2279 31867 2335
rect 31809 2255 31812 2279
rect 31864 2255 31867 2279
rect 31809 2199 31810 2255
rect 31866 2199 31867 2255
rect 31809 2185 31812 2199
rect 31864 2185 31867 2199
rect 31809 2175 31867 2185
rect 31809 2119 31810 2175
rect 31866 2119 31867 2175
rect 31809 2109 31867 2119
rect 31809 2095 31812 2109
rect 31864 2095 31867 2109
rect 31809 2039 31810 2095
rect 31866 2039 31867 2095
rect 31809 2015 31812 2039
rect 31864 2015 31867 2039
rect 31809 1959 31810 2015
rect 31866 1959 31867 2015
rect 31809 1935 31812 1959
rect 31864 1935 31867 1959
rect 31809 1879 31810 1935
rect 31866 1879 31867 1935
rect 31809 1865 31812 1879
rect 31864 1865 31867 1879
rect 31809 1855 31867 1865
rect 31809 1799 31810 1855
rect 31866 1799 31867 1855
rect 31809 1789 31867 1799
rect 31809 1775 31812 1789
rect 31864 1775 31867 1789
rect 31809 1719 31810 1775
rect 31866 1719 31867 1775
rect 31809 1695 31812 1719
rect 31864 1695 31867 1719
rect 31809 1639 31810 1695
rect 31866 1639 31867 1695
rect 31809 1615 31812 1639
rect 31864 1615 31867 1639
rect 31809 1559 31810 1615
rect 31866 1559 31867 1615
rect 31809 1545 31812 1559
rect 31864 1545 31867 1559
rect 31809 1535 31867 1545
rect 31809 1479 31810 1535
rect 31866 1479 31867 1535
rect 31809 1469 31867 1479
rect 31809 1455 31812 1469
rect 31864 1455 31867 1469
rect 31809 1399 31810 1455
rect 31866 1399 31867 1455
rect 31809 1375 31812 1399
rect 31864 1375 31867 1399
rect 31809 1319 31810 1375
rect 31866 1319 31867 1375
rect 31809 1295 31812 1319
rect 31864 1295 31867 1319
rect 31809 1239 31810 1295
rect 31866 1239 31867 1295
rect 31809 1225 31812 1239
rect 31864 1225 31867 1239
rect 31809 1215 31867 1225
rect 31809 1159 31810 1215
rect 31866 1159 31867 1215
rect 31809 1147 31867 1159
rect 31905 3133 31963 3147
rect 31905 3081 31908 3133
rect 31960 3081 31963 3133
rect 31905 3069 31963 3081
rect 31905 3017 31908 3069
rect 31960 3017 31963 3069
rect 31905 3005 31963 3017
rect 31905 2953 31908 3005
rect 31960 2953 31963 3005
rect 31905 2941 31963 2953
rect 31905 2889 31908 2941
rect 31960 2889 31963 2941
rect 31905 2877 31963 2889
rect 31905 2825 31908 2877
rect 31960 2825 31963 2877
rect 31905 2813 31963 2825
rect 31905 2761 31908 2813
rect 31960 2761 31963 2813
rect 31905 2749 31963 2761
rect 31905 2697 31908 2749
rect 31960 2697 31963 2749
rect 31905 2685 31963 2697
rect 31905 2633 31908 2685
rect 31960 2633 31963 2685
rect 31905 2621 31963 2633
rect 31905 2569 31908 2621
rect 31960 2569 31963 2621
rect 31905 2557 31963 2569
rect 31905 2505 31908 2557
rect 31960 2505 31963 2557
rect 31905 2493 31963 2505
rect 31905 2441 31908 2493
rect 31960 2441 31963 2493
rect 31905 2429 31963 2441
rect 31905 2377 31908 2429
rect 31960 2377 31963 2429
rect 31905 2365 31963 2377
rect 31905 2313 31908 2365
rect 31960 2313 31963 2365
rect 31905 2301 31963 2313
rect 31905 2249 31908 2301
rect 31960 2249 31963 2301
rect 31905 2237 31963 2249
rect 31905 2185 31908 2237
rect 31960 2185 31963 2237
rect 31905 2173 31963 2185
rect 31905 2121 31908 2173
rect 31960 2121 31963 2173
rect 31905 2109 31963 2121
rect 31905 2057 31908 2109
rect 31960 2057 31963 2109
rect 31905 2045 31963 2057
rect 31905 1993 31908 2045
rect 31960 1993 31963 2045
rect 31905 1981 31963 1993
rect 31905 1929 31908 1981
rect 31960 1929 31963 1981
rect 31905 1917 31963 1929
rect 31905 1865 31908 1917
rect 31960 1865 31963 1917
rect 31905 1853 31963 1865
rect 31905 1801 31908 1853
rect 31960 1801 31963 1853
rect 31905 1789 31963 1801
rect 31905 1737 31908 1789
rect 31960 1737 31963 1789
rect 31905 1725 31963 1737
rect 31905 1673 31908 1725
rect 31960 1673 31963 1725
rect 31905 1661 31963 1673
rect 31905 1609 31908 1661
rect 31960 1609 31963 1661
rect 31905 1597 31963 1609
rect 31905 1545 31908 1597
rect 31960 1545 31963 1597
rect 31905 1533 31963 1545
rect 31905 1481 31908 1533
rect 31960 1481 31963 1533
rect 31905 1469 31963 1481
rect 31905 1417 31908 1469
rect 31960 1417 31963 1469
rect 31905 1405 31963 1417
rect 31905 1353 31908 1405
rect 31960 1353 31963 1405
rect 31905 1341 31963 1353
rect 31905 1289 31908 1341
rect 31960 1289 31963 1341
rect 31905 1277 31963 1289
rect 31905 1225 31908 1277
rect 31960 1225 31963 1277
rect 31905 1213 31963 1225
rect 31905 1161 31908 1213
rect 31960 1161 31963 1213
rect 31905 830 31963 1161
rect 32001 3135 32059 3147
rect 32001 3079 32002 3135
rect 32058 3079 32059 3135
rect 32001 3069 32059 3079
rect 32001 3055 32004 3069
rect 32056 3055 32059 3069
rect 32001 2999 32002 3055
rect 32058 2999 32059 3055
rect 32001 2975 32004 2999
rect 32056 2975 32059 2999
rect 32001 2919 32002 2975
rect 32058 2919 32059 2975
rect 32001 2895 32004 2919
rect 32056 2895 32059 2919
rect 32001 2839 32002 2895
rect 32058 2839 32059 2895
rect 32001 2825 32004 2839
rect 32056 2825 32059 2839
rect 32001 2815 32059 2825
rect 32001 2759 32002 2815
rect 32058 2759 32059 2815
rect 32001 2749 32059 2759
rect 32001 2735 32004 2749
rect 32056 2735 32059 2749
rect 32001 2679 32002 2735
rect 32058 2679 32059 2735
rect 32001 2655 32004 2679
rect 32056 2655 32059 2679
rect 32001 2599 32002 2655
rect 32058 2599 32059 2655
rect 32001 2575 32004 2599
rect 32056 2575 32059 2599
rect 32001 2519 32002 2575
rect 32058 2519 32059 2575
rect 32001 2505 32004 2519
rect 32056 2505 32059 2519
rect 32001 2495 32059 2505
rect 32001 2439 32002 2495
rect 32058 2439 32059 2495
rect 32001 2429 32059 2439
rect 32001 2415 32004 2429
rect 32056 2415 32059 2429
rect 32001 2359 32002 2415
rect 32058 2359 32059 2415
rect 32001 2335 32004 2359
rect 32056 2335 32059 2359
rect 32001 2279 32002 2335
rect 32058 2279 32059 2335
rect 32001 2255 32004 2279
rect 32056 2255 32059 2279
rect 32001 2199 32002 2255
rect 32058 2199 32059 2255
rect 32001 2185 32004 2199
rect 32056 2185 32059 2199
rect 32001 2175 32059 2185
rect 32001 2119 32002 2175
rect 32058 2119 32059 2175
rect 32001 2109 32059 2119
rect 32001 2095 32004 2109
rect 32056 2095 32059 2109
rect 32001 2039 32002 2095
rect 32058 2039 32059 2095
rect 32001 2015 32004 2039
rect 32056 2015 32059 2039
rect 32001 1959 32002 2015
rect 32058 1959 32059 2015
rect 32001 1935 32004 1959
rect 32056 1935 32059 1959
rect 32001 1879 32002 1935
rect 32058 1879 32059 1935
rect 32001 1865 32004 1879
rect 32056 1865 32059 1879
rect 32001 1855 32059 1865
rect 32001 1799 32002 1855
rect 32058 1799 32059 1855
rect 32001 1789 32059 1799
rect 32001 1775 32004 1789
rect 32056 1775 32059 1789
rect 32001 1719 32002 1775
rect 32058 1719 32059 1775
rect 32001 1695 32004 1719
rect 32056 1695 32059 1719
rect 32001 1639 32002 1695
rect 32058 1639 32059 1695
rect 32001 1615 32004 1639
rect 32056 1615 32059 1639
rect 32001 1559 32002 1615
rect 32058 1559 32059 1615
rect 32001 1545 32004 1559
rect 32056 1545 32059 1559
rect 32001 1535 32059 1545
rect 32001 1479 32002 1535
rect 32058 1479 32059 1535
rect 32001 1469 32059 1479
rect 32001 1455 32004 1469
rect 32056 1455 32059 1469
rect 32001 1399 32002 1455
rect 32058 1399 32059 1455
rect 32001 1375 32004 1399
rect 32056 1375 32059 1399
rect 32001 1319 32002 1375
rect 32058 1319 32059 1375
rect 32001 1295 32004 1319
rect 32056 1295 32059 1319
rect 32001 1239 32002 1295
rect 32058 1239 32059 1295
rect 32001 1225 32004 1239
rect 32056 1225 32059 1239
rect 32001 1215 32059 1225
rect 32001 1159 32002 1215
rect 32058 1159 32059 1215
rect 32001 1147 32059 1159
rect 32097 3133 32155 3147
rect 32097 3081 32100 3133
rect 32152 3081 32155 3133
rect 32097 3069 32155 3081
rect 32097 3017 32100 3069
rect 32152 3017 32155 3069
rect 32097 3005 32155 3017
rect 32097 2953 32100 3005
rect 32152 2953 32155 3005
rect 32097 2941 32155 2953
rect 32097 2889 32100 2941
rect 32152 2889 32155 2941
rect 32097 2877 32155 2889
rect 32097 2825 32100 2877
rect 32152 2825 32155 2877
rect 32097 2813 32155 2825
rect 32097 2761 32100 2813
rect 32152 2761 32155 2813
rect 32097 2749 32155 2761
rect 32097 2697 32100 2749
rect 32152 2697 32155 2749
rect 32097 2685 32155 2697
rect 32097 2633 32100 2685
rect 32152 2633 32155 2685
rect 32097 2621 32155 2633
rect 32097 2569 32100 2621
rect 32152 2569 32155 2621
rect 32097 2557 32155 2569
rect 32097 2505 32100 2557
rect 32152 2505 32155 2557
rect 32097 2493 32155 2505
rect 32097 2441 32100 2493
rect 32152 2441 32155 2493
rect 32097 2429 32155 2441
rect 32097 2377 32100 2429
rect 32152 2377 32155 2429
rect 32097 2365 32155 2377
rect 32097 2313 32100 2365
rect 32152 2313 32155 2365
rect 32097 2301 32155 2313
rect 32097 2249 32100 2301
rect 32152 2249 32155 2301
rect 32097 2237 32155 2249
rect 32097 2185 32100 2237
rect 32152 2185 32155 2237
rect 32097 2173 32155 2185
rect 32097 2121 32100 2173
rect 32152 2121 32155 2173
rect 32097 2109 32155 2121
rect 32097 2057 32100 2109
rect 32152 2057 32155 2109
rect 32097 2045 32155 2057
rect 32097 1993 32100 2045
rect 32152 1993 32155 2045
rect 32097 1981 32155 1993
rect 32097 1929 32100 1981
rect 32152 1929 32155 1981
rect 32097 1917 32155 1929
rect 32097 1865 32100 1917
rect 32152 1865 32155 1917
rect 32097 1853 32155 1865
rect 32097 1801 32100 1853
rect 32152 1801 32155 1853
rect 32097 1789 32155 1801
rect 32097 1737 32100 1789
rect 32152 1737 32155 1789
rect 32097 1725 32155 1737
rect 32097 1673 32100 1725
rect 32152 1673 32155 1725
rect 32097 1661 32155 1673
rect 32097 1609 32100 1661
rect 32152 1609 32155 1661
rect 32097 1597 32155 1609
rect 32097 1545 32100 1597
rect 32152 1545 32155 1597
rect 32097 1533 32155 1545
rect 32097 1481 32100 1533
rect 32152 1481 32155 1533
rect 32097 1469 32155 1481
rect 32097 1417 32100 1469
rect 32152 1417 32155 1469
rect 32097 1405 32155 1417
rect 32097 1353 32100 1405
rect 32152 1353 32155 1405
rect 32097 1341 32155 1353
rect 32097 1289 32100 1341
rect 32152 1289 32155 1341
rect 32097 1277 32155 1289
rect 32097 1225 32100 1277
rect 32152 1225 32155 1277
rect 32097 1213 32155 1225
rect 32097 1161 32100 1213
rect 32152 1161 32155 1213
rect 32097 830 32155 1161
rect 32193 3135 32251 3147
rect 32193 3079 32194 3135
rect 32250 3079 32251 3135
rect 32193 3069 32251 3079
rect 32193 3055 32196 3069
rect 32248 3055 32251 3069
rect 32193 2999 32194 3055
rect 32250 2999 32251 3055
rect 32193 2975 32196 2999
rect 32248 2975 32251 2999
rect 32193 2919 32194 2975
rect 32250 2919 32251 2975
rect 32193 2895 32196 2919
rect 32248 2895 32251 2919
rect 32193 2839 32194 2895
rect 32250 2839 32251 2895
rect 32193 2825 32196 2839
rect 32248 2825 32251 2839
rect 32193 2815 32251 2825
rect 32193 2759 32194 2815
rect 32250 2759 32251 2815
rect 32193 2749 32251 2759
rect 32193 2735 32196 2749
rect 32248 2735 32251 2749
rect 32193 2679 32194 2735
rect 32250 2679 32251 2735
rect 32193 2655 32196 2679
rect 32248 2655 32251 2679
rect 32193 2599 32194 2655
rect 32250 2599 32251 2655
rect 32193 2575 32196 2599
rect 32248 2575 32251 2599
rect 32193 2519 32194 2575
rect 32250 2519 32251 2575
rect 32193 2505 32196 2519
rect 32248 2505 32251 2519
rect 32193 2495 32251 2505
rect 32193 2439 32194 2495
rect 32250 2439 32251 2495
rect 32193 2429 32251 2439
rect 32193 2415 32196 2429
rect 32248 2415 32251 2429
rect 32193 2359 32194 2415
rect 32250 2359 32251 2415
rect 32193 2335 32196 2359
rect 32248 2335 32251 2359
rect 32193 2279 32194 2335
rect 32250 2279 32251 2335
rect 32193 2255 32196 2279
rect 32248 2255 32251 2279
rect 32193 2199 32194 2255
rect 32250 2199 32251 2255
rect 32193 2185 32196 2199
rect 32248 2185 32251 2199
rect 32193 2175 32251 2185
rect 32193 2119 32194 2175
rect 32250 2119 32251 2175
rect 32193 2109 32251 2119
rect 32193 2095 32196 2109
rect 32248 2095 32251 2109
rect 32193 2039 32194 2095
rect 32250 2039 32251 2095
rect 32193 2015 32196 2039
rect 32248 2015 32251 2039
rect 32193 1959 32194 2015
rect 32250 1959 32251 2015
rect 32193 1935 32196 1959
rect 32248 1935 32251 1959
rect 32193 1879 32194 1935
rect 32250 1879 32251 1935
rect 32193 1865 32196 1879
rect 32248 1865 32251 1879
rect 32193 1855 32251 1865
rect 32193 1799 32194 1855
rect 32250 1799 32251 1855
rect 32193 1789 32251 1799
rect 32193 1775 32196 1789
rect 32248 1775 32251 1789
rect 32193 1719 32194 1775
rect 32250 1719 32251 1775
rect 32193 1695 32196 1719
rect 32248 1695 32251 1719
rect 32193 1639 32194 1695
rect 32250 1639 32251 1695
rect 32193 1615 32196 1639
rect 32248 1615 32251 1639
rect 32193 1559 32194 1615
rect 32250 1559 32251 1615
rect 32193 1545 32196 1559
rect 32248 1545 32251 1559
rect 32193 1535 32251 1545
rect 32193 1479 32194 1535
rect 32250 1479 32251 1535
rect 32193 1469 32251 1479
rect 32193 1455 32196 1469
rect 32248 1455 32251 1469
rect 32193 1399 32194 1455
rect 32250 1399 32251 1455
rect 32193 1375 32196 1399
rect 32248 1375 32251 1399
rect 32193 1319 32194 1375
rect 32250 1319 32251 1375
rect 32193 1295 32196 1319
rect 32248 1295 32251 1319
rect 32193 1239 32194 1295
rect 32250 1239 32251 1295
rect 32193 1225 32196 1239
rect 32248 1225 32251 1239
rect 32193 1215 32251 1225
rect 32193 1159 32194 1215
rect 32250 1159 32251 1215
rect 32193 1147 32251 1159
rect 32289 3133 32347 3147
rect 32289 3081 32292 3133
rect 32344 3081 32347 3133
rect 32289 3069 32347 3081
rect 32289 3017 32292 3069
rect 32344 3017 32347 3069
rect 32289 3005 32347 3017
rect 32289 2953 32292 3005
rect 32344 2953 32347 3005
rect 32289 2941 32347 2953
rect 32289 2889 32292 2941
rect 32344 2889 32347 2941
rect 32289 2877 32347 2889
rect 32289 2825 32292 2877
rect 32344 2825 32347 2877
rect 32289 2813 32347 2825
rect 32289 2761 32292 2813
rect 32344 2761 32347 2813
rect 32289 2749 32347 2761
rect 32289 2697 32292 2749
rect 32344 2697 32347 2749
rect 32289 2685 32347 2697
rect 32289 2633 32292 2685
rect 32344 2633 32347 2685
rect 32289 2621 32347 2633
rect 32289 2569 32292 2621
rect 32344 2569 32347 2621
rect 32289 2557 32347 2569
rect 32289 2505 32292 2557
rect 32344 2505 32347 2557
rect 32289 2493 32347 2505
rect 32289 2441 32292 2493
rect 32344 2441 32347 2493
rect 32289 2429 32347 2441
rect 32289 2377 32292 2429
rect 32344 2377 32347 2429
rect 32289 2365 32347 2377
rect 32289 2313 32292 2365
rect 32344 2313 32347 2365
rect 32289 2301 32347 2313
rect 32289 2249 32292 2301
rect 32344 2249 32347 2301
rect 32289 2237 32347 2249
rect 32289 2185 32292 2237
rect 32344 2185 32347 2237
rect 32289 2173 32347 2185
rect 32289 2121 32292 2173
rect 32344 2121 32347 2173
rect 32289 2109 32347 2121
rect 32289 2057 32292 2109
rect 32344 2057 32347 2109
rect 32289 2045 32347 2057
rect 32289 1993 32292 2045
rect 32344 1993 32347 2045
rect 32289 1981 32347 1993
rect 32289 1929 32292 1981
rect 32344 1929 32347 1981
rect 32289 1917 32347 1929
rect 32289 1865 32292 1917
rect 32344 1865 32347 1917
rect 32289 1853 32347 1865
rect 32289 1801 32292 1853
rect 32344 1801 32347 1853
rect 32289 1789 32347 1801
rect 32289 1737 32292 1789
rect 32344 1737 32347 1789
rect 32289 1725 32347 1737
rect 32289 1673 32292 1725
rect 32344 1673 32347 1725
rect 32289 1661 32347 1673
rect 32289 1609 32292 1661
rect 32344 1609 32347 1661
rect 32289 1597 32347 1609
rect 32289 1545 32292 1597
rect 32344 1545 32347 1597
rect 32289 1533 32347 1545
rect 32289 1481 32292 1533
rect 32344 1481 32347 1533
rect 32289 1469 32347 1481
rect 32289 1417 32292 1469
rect 32344 1417 32347 1469
rect 32289 1405 32347 1417
rect 32289 1353 32292 1405
rect 32344 1353 32347 1405
rect 32289 1341 32347 1353
rect 32289 1289 32292 1341
rect 32344 1289 32347 1341
rect 32289 1277 32347 1289
rect 32289 1225 32292 1277
rect 32344 1225 32347 1277
rect 32289 1213 32347 1225
rect 32289 1161 32292 1213
rect 32344 1161 32347 1213
rect 32289 830 32347 1161
rect 32385 3135 32443 3147
rect 32385 3079 32386 3135
rect 32442 3079 32443 3135
rect 32385 3069 32443 3079
rect 32385 3055 32388 3069
rect 32440 3055 32443 3069
rect 32385 2999 32386 3055
rect 32442 2999 32443 3055
rect 32385 2975 32388 2999
rect 32440 2975 32443 2999
rect 32385 2919 32386 2975
rect 32442 2919 32443 2975
rect 32385 2895 32388 2919
rect 32440 2895 32443 2919
rect 32385 2839 32386 2895
rect 32442 2839 32443 2895
rect 32385 2825 32388 2839
rect 32440 2825 32443 2839
rect 32385 2815 32443 2825
rect 32385 2759 32386 2815
rect 32442 2759 32443 2815
rect 32385 2749 32443 2759
rect 32385 2735 32388 2749
rect 32440 2735 32443 2749
rect 32385 2679 32386 2735
rect 32442 2679 32443 2735
rect 32385 2655 32388 2679
rect 32440 2655 32443 2679
rect 32385 2599 32386 2655
rect 32442 2599 32443 2655
rect 32385 2575 32388 2599
rect 32440 2575 32443 2599
rect 32385 2519 32386 2575
rect 32442 2519 32443 2575
rect 32385 2505 32388 2519
rect 32440 2505 32443 2519
rect 32385 2495 32443 2505
rect 32385 2439 32386 2495
rect 32442 2439 32443 2495
rect 32385 2429 32443 2439
rect 32385 2415 32388 2429
rect 32440 2415 32443 2429
rect 32385 2359 32386 2415
rect 32442 2359 32443 2415
rect 32385 2335 32388 2359
rect 32440 2335 32443 2359
rect 32385 2279 32386 2335
rect 32442 2279 32443 2335
rect 32385 2255 32388 2279
rect 32440 2255 32443 2279
rect 32385 2199 32386 2255
rect 32442 2199 32443 2255
rect 32385 2185 32388 2199
rect 32440 2185 32443 2199
rect 32385 2175 32443 2185
rect 32385 2119 32386 2175
rect 32442 2119 32443 2175
rect 32385 2109 32443 2119
rect 32385 2095 32388 2109
rect 32440 2095 32443 2109
rect 32385 2039 32386 2095
rect 32442 2039 32443 2095
rect 32385 2015 32388 2039
rect 32440 2015 32443 2039
rect 32385 1959 32386 2015
rect 32442 1959 32443 2015
rect 32385 1935 32388 1959
rect 32440 1935 32443 1959
rect 32385 1879 32386 1935
rect 32442 1879 32443 1935
rect 32385 1865 32388 1879
rect 32440 1865 32443 1879
rect 32385 1855 32443 1865
rect 32385 1799 32386 1855
rect 32442 1799 32443 1855
rect 32385 1789 32443 1799
rect 32385 1775 32388 1789
rect 32440 1775 32443 1789
rect 32385 1719 32386 1775
rect 32442 1719 32443 1775
rect 32385 1695 32388 1719
rect 32440 1695 32443 1719
rect 32385 1639 32386 1695
rect 32442 1639 32443 1695
rect 32385 1615 32388 1639
rect 32440 1615 32443 1639
rect 32385 1559 32386 1615
rect 32442 1559 32443 1615
rect 32385 1545 32388 1559
rect 32440 1545 32443 1559
rect 32385 1535 32443 1545
rect 32385 1479 32386 1535
rect 32442 1479 32443 1535
rect 32385 1469 32443 1479
rect 32385 1455 32388 1469
rect 32440 1455 32443 1469
rect 32385 1399 32386 1455
rect 32442 1399 32443 1455
rect 32385 1375 32388 1399
rect 32440 1375 32443 1399
rect 32385 1319 32386 1375
rect 32442 1319 32443 1375
rect 32385 1295 32388 1319
rect 32440 1295 32443 1319
rect 32385 1239 32386 1295
rect 32442 1239 32443 1295
rect 32385 1225 32388 1239
rect 32440 1225 32443 1239
rect 32385 1215 32443 1225
rect 32385 1159 32386 1215
rect 32442 1159 32443 1215
rect 32385 1147 32443 1159
rect 32481 3133 32539 3147
rect 32481 3081 32484 3133
rect 32536 3081 32539 3133
rect 32481 3069 32539 3081
rect 32481 3017 32484 3069
rect 32536 3017 32539 3069
rect 32481 3005 32539 3017
rect 32481 2953 32484 3005
rect 32536 2953 32539 3005
rect 32481 2941 32539 2953
rect 32481 2889 32484 2941
rect 32536 2889 32539 2941
rect 32481 2877 32539 2889
rect 32481 2825 32484 2877
rect 32536 2825 32539 2877
rect 32481 2813 32539 2825
rect 32481 2761 32484 2813
rect 32536 2761 32539 2813
rect 32481 2749 32539 2761
rect 32481 2697 32484 2749
rect 32536 2697 32539 2749
rect 32481 2685 32539 2697
rect 32481 2633 32484 2685
rect 32536 2633 32539 2685
rect 32481 2621 32539 2633
rect 32481 2569 32484 2621
rect 32536 2569 32539 2621
rect 32481 2557 32539 2569
rect 32481 2505 32484 2557
rect 32536 2505 32539 2557
rect 32481 2493 32539 2505
rect 32481 2441 32484 2493
rect 32536 2441 32539 2493
rect 32481 2429 32539 2441
rect 32481 2377 32484 2429
rect 32536 2377 32539 2429
rect 32481 2365 32539 2377
rect 32481 2313 32484 2365
rect 32536 2313 32539 2365
rect 32481 2301 32539 2313
rect 32481 2249 32484 2301
rect 32536 2249 32539 2301
rect 32481 2237 32539 2249
rect 32481 2185 32484 2237
rect 32536 2185 32539 2237
rect 32481 2173 32539 2185
rect 32481 2121 32484 2173
rect 32536 2121 32539 2173
rect 32481 2109 32539 2121
rect 32481 2057 32484 2109
rect 32536 2057 32539 2109
rect 32481 2045 32539 2057
rect 32481 1993 32484 2045
rect 32536 1993 32539 2045
rect 32481 1981 32539 1993
rect 32481 1929 32484 1981
rect 32536 1929 32539 1981
rect 32481 1917 32539 1929
rect 32481 1865 32484 1917
rect 32536 1865 32539 1917
rect 32481 1853 32539 1865
rect 32481 1801 32484 1853
rect 32536 1801 32539 1853
rect 32481 1789 32539 1801
rect 32481 1737 32484 1789
rect 32536 1737 32539 1789
rect 32481 1725 32539 1737
rect 32481 1673 32484 1725
rect 32536 1673 32539 1725
rect 32481 1661 32539 1673
rect 32481 1609 32484 1661
rect 32536 1609 32539 1661
rect 32481 1597 32539 1609
rect 32481 1545 32484 1597
rect 32536 1545 32539 1597
rect 32481 1533 32539 1545
rect 32481 1481 32484 1533
rect 32536 1481 32539 1533
rect 32481 1469 32539 1481
rect 32481 1417 32484 1469
rect 32536 1417 32539 1469
rect 32481 1405 32539 1417
rect 32481 1353 32484 1405
rect 32536 1353 32539 1405
rect 32481 1341 32539 1353
rect 32481 1289 32484 1341
rect 32536 1289 32539 1341
rect 32481 1277 32539 1289
rect 32481 1225 32484 1277
rect 32536 1225 32539 1277
rect 32481 1213 32539 1225
rect 32481 1161 32484 1213
rect 32536 1161 32539 1213
rect 32481 830 32539 1161
rect 32577 3135 32635 3147
rect 32577 3079 32578 3135
rect 32634 3079 32635 3135
rect 32577 3069 32635 3079
rect 32577 3055 32580 3069
rect 32632 3055 32635 3069
rect 32577 2999 32578 3055
rect 32634 2999 32635 3055
rect 32577 2975 32580 2999
rect 32632 2975 32635 2999
rect 32577 2919 32578 2975
rect 32634 2919 32635 2975
rect 32577 2895 32580 2919
rect 32632 2895 32635 2919
rect 32577 2839 32578 2895
rect 32634 2839 32635 2895
rect 32577 2825 32580 2839
rect 32632 2825 32635 2839
rect 32577 2815 32635 2825
rect 32577 2759 32578 2815
rect 32634 2759 32635 2815
rect 32577 2749 32635 2759
rect 32577 2735 32580 2749
rect 32632 2735 32635 2749
rect 32577 2679 32578 2735
rect 32634 2679 32635 2735
rect 32577 2655 32580 2679
rect 32632 2655 32635 2679
rect 32577 2599 32578 2655
rect 32634 2599 32635 2655
rect 32577 2575 32580 2599
rect 32632 2575 32635 2599
rect 32577 2519 32578 2575
rect 32634 2519 32635 2575
rect 32577 2505 32580 2519
rect 32632 2505 32635 2519
rect 32577 2495 32635 2505
rect 32577 2439 32578 2495
rect 32634 2439 32635 2495
rect 32577 2429 32635 2439
rect 32577 2415 32580 2429
rect 32632 2415 32635 2429
rect 32577 2359 32578 2415
rect 32634 2359 32635 2415
rect 32577 2335 32580 2359
rect 32632 2335 32635 2359
rect 32577 2279 32578 2335
rect 32634 2279 32635 2335
rect 32577 2255 32580 2279
rect 32632 2255 32635 2279
rect 32577 2199 32578 2255
rect 32634 2199 32635 2255
rect 32577 2185 32580 2199
rect 32632 2185 32635 2199
rect 32577 2175 32635 2185
rect 32577 2119 32578 2175
rect 32634 2119 32635 2175
rect 32577 2109 32635 2119
rect 32577 2095 32580 2109
rect 32632 2095 32635 2109
rect 32577 2039 32578 2095
rect 32634 2039 32635 2095
rect 32577 2015 32580 2039
rect 32632 2015 32635 2039
rect 32577 1959 32578 2015
rect 32634 1959 32635 2015
rect 32577 1935 32580 1959
rect 32632 1935 32635 1959
rect 32577 1879 32578 1935
rect 32634 1879 32635 1935
rect 32577 1865 32580 1879
rect 32632 1865 32635 1879
rect 32577 1855 32635 1865
rect 32577 1799 32578 1855
rect 32634 1799 32635 1855
rect 32577 1789 32635 1799
rect 32577 1775 32580 1789
rect 32632 1775 32635 1789
rect 32577 1719 32578 1775
rect 32634 1719 32635 1775
rect 32577 1695 32580 1719
rect 32632 1695 32635 1719
rect 32577 1639 32578 1695
rect 32634 1639 32635 1695
rect 32577 1615 32580 1639
rect 32632 1615 32635 1639
rect 32577 1559 32578 1615
rect 32634 1559 32635 1615
rect 32577 1545 32580 1559
rect 32632 1545 32635 1559
rect 32577 1535 32635 1545
rect 32577 1479 32578 1535
rect 32634 1479 32635 1535
rect 32577 1469 32635 1479
rect 32577 1455 32580 1469
rect 32632 1455 32635 1469
rect 32577 1399 32578 1455
rect 32634 1399 32635 1455
rect 32577 1375 32580 1399
rect 32632 1375 32635 1399
rect 32577 1319 32578 1375
rect 32634 1319 32635 1375
rect 32577 1295 32580 1319
rect 32632 1295 32635 1319
rect 32577 1239 32578 1295
rect 32634 1239 32635 1295
rect 32577 1225 32580 1239
rect 32632 1225 32635 1239
rect 32577 1215 32635 1225
rect 32577 1159 32578 1215
rect 32634 1159 32635 1215
rect 32577 1147 32635 1159
rect 32673 3133 32731 3147
rect 32673 3081 32676 3133
rect 32728 3081 32731 3133
rect 32673 3069 32731 3081
rect 32673 3017 32676 3069
rect 32728 3017 32731 3069
rect 32673 3005 32731 3017
rect 32673 2953 32676 3005
rect 32728 2953 32731 3005
rect 32673 2941 32731 2953
rect 32673 2889 32676 2941
rect 32728 2889 32731 2941
rect 32673 2877 32731 2889
rect 32673 2825 32676 2877
rect 32728 2825 32731 2877
rect 32673 2813 32731 2825
rect 32673 2761 32676 2813
rect 32728 2761 32731 2813
rect 32673 2749 32731 2761
rect 32673 2697 32676 2749
rect 32728 2697 32731 2749
rect 32673 2685 32731 2697
rect 32673 2633 32676 2685
rect 32728 2633 32731 2685
rect 32673 2621 32731 2633
rect 32673 2569 32676 2621
rect 32728 2569 32731 2621
rect 32673 2557 32731 2569
rect 32673 2505 32676 2557
rect 32728 2505 32731 2557
rect 32673 2493 32731 2505
rect 32673 2441 32676 2493
rect 32728 2441 32731 2493
rect 32673 2429 32731 2441
rect 32673 2377 32676 2429
rect 32728 2377 32731 2429
rect 32673 2365 32731 2377
rect 32673 2313 32676 2365
rect 32728 2313 32731 2365
rect 32673 2301 32731 2313
rect 32673 2249 32676 2301
rect 32728 2249 32731 2301
rect 32673 2237 32731 2249
rect 32673 2185 32676 2237
rect 32728 2185 32731 2237
rect 32673 2173 32731 2185
rect 32673 2121 32676 2173
rect 32728 2121 32731 2173
rect 32673 2109 32731 2121
rect 32673 2057 32676 2109
rect 32728 2057 32731 2109
rect 32673 2045 32731 2057
rect 32673 1993 32676 2045
rect 32728 1993 32731 2045
rect 32673 1981 32731 1993
rect 32673 1929 32676 1981
rect 32728 1929 32731 1981
rect 32673 1917 32731 1929
rect 32673 1865 32676 1917
rect 32728 1865 32731 1917
rect 32673 1853 32731 1865
rect 32673 1801 32676 1853
rect 32728 1801 32731 1853
rect 32673 1789 32731 1801
rect 32673 1737 32676 1789
rect 32728 1737 32731 1789
rect 32673 1725 32731 1737
rect 32673 1673 32676 1725
rect 32728 1673 32731 1725
rect 32673 1661 32731 1673
rect 32673 1609 32676 1661
rect 32728 1609 32731 1661
rect 32673 1597 32731 1609
rect 32673 1545 32676 1597
rect 32728 1545 32731 1597
rect 32673 1533 32731 1545
rect 32673 1481 32676 1533
rect 32728 1481 32731 1533
rect 32673 1469 32731 1481
rect 32673 1417 32676 1469
rect 32728 1417 32731 1469
rect 32673 1405 32731 1417
rect 32673 1353 32676 1405
rect 32728 1353 32731 1405
rect 32673 1341 32731 1353
rect 32673 1289 32676 1341
rect 32728 1289 32731 1341
rect 32673 1277 32731 1289
rect 32673 1225 32676 1277
rect 32728 1225 32731 1277
rect 32673 1213 32731 1225
rect 32673 1161 32676 1213
rect 32728 1161 32731 1213
rect 32673 830 32731 1161
rect 32769 3135 32827 3147
rect 32769 3079 32770 3135
rect 32826 3079 32827 3135
rect 32769 3069 32827 3079
rect 32769 3055 32772 3069
rect 32824 3055 32827 3069
rect 32769 2999 32770 3055
rect 32826 2999 32827 3055
rect 32769 2975 32772 2999
rect 32824 2975 32827 2999
rect 32769 2919 32770 2975
rect 32826 2919 32827 2975
rect 32769 2895 32772 2919
rect 32824 2895 32827 2919
rect 32769 2839 32770 2895
rect 32826 2839 32827 2895
rect 32769 2825 32772 2839
rect 32824 2825 32827 2839
rect 32769 2815 32827 2825
rect 32769 2759 32770 2815
rect 32826 2759 32827 2815
rect 32769 2749 32827 2759
rect 32769 2735 32772 2749
rect 32824 2735 32827 2749
rect 32769 2679 32770 2735
rect 32826 2679 32827 2735
rect 32769 2655 32772 2679
rect 32824 2655 32827 2679
rect 32769 2599 32770 2655
rect 32826 2599 32827 2655
rect 32769 2575 32772 2599
rect 32824 2575 32827 2599
rect 32769 2519 32770 2575
rect 32826 2519 32827 2575
rect 32769 2505 32772 2519
rect 32824 2505 32827 2519
rect 32769 2495 32827 2505
rect 32769 2439 32770 2495
rect 32826 2439 32827 2495
rect 32769 2429 32827 2439
rect 32769 2415 32772 2429
rect 32824 2415 32827 2429
rect 32769 2359 32770 2415
rect 32826 2359 32827 2415
rect 32769 2335 32772 2359
rect 32824 2335 32827 2359
rect 32769 2279 32770 2335
rect 32826 2279 32827 2335
rect 32769 2255 32772 2279
rect 32824 2255 32827 2279
rect 32769 2199 32770 2255
rect 32826 2199 32827 2255
rect 32769 2185 32772 2199
rect 32824 2185 32827 2199
rect 32769 2175 32827 2185
rect 32769 2119 32770 2175
rect 32826 2119 32827 2175
rect 32769 2109 32827 2119
rect 32769 2095 32772 2109
rect 32824 2095 32827 2109
rect 32769 2039 32770 2095
rect 32826 2039 32827 2095
rect 32769 2015 32772 2039
rect 32824 2015 32827 2039
rect 32769 1959 32770 2015
rect 32826 1959 32827 2015
rect 32769 1935 32772 1959
rect 32824 1935 32827 1959
rect 32769 1879 32770 1935
rect 32826 1879 32827 1935
rect 32769 1865 32772 1879
rect 32824 1865 32827 1879
rect 32769 1855 32827 1865
rect 32769 1799 32770 1855
rect 32826 1799 32827 1855
rect 32769 1789 32827 1799
rect 32769 1775 32772 1789
rect 32824 1775 32827 1789
rect 32769 1719 32770 1775
rect 32826 1719 32827 1775
rect 32769 1695 32772 1719
rect 32824 1695 32827 1719
rect 32769 1639 32770 1695
rect 32826 1639 32827 1695
rect 32769 1615 32772 1639
rect 32824 1615 32827 1639
rect 32769 1559 32770 1615
rect 32826 1559 32827 1615
rect 32769 1545 32772 1559
rect 32824 1545 32827 1559
rect 32769 1535 32827 1545
rect 32769 1479 32770 1535
rect 32826 1479 32827 1535
rect 32769 1469 32827 1479
rect 32769 1455 32772 1469
rect 32824 1455 32827 1469
rect 32769 1399 32770 1455
rect 32826 1399 32827 1455
rect 32769 1375 32772 1399
rect 32824 1375 32827 1399
rect 32769 1319 32770 1375
rect 32826 1319 32827 1375
rect 32769 1295 32772 1319
rect 32824 1295 32827 1319
rect 32769 1239 32770 1295
rect 32826 1239 32827 1295
rect 32769 1225 32772 1239
rect 32824 1225 32827 1239
rect 32769 1215 32827 1225
rect 32769 1159 32770 1215
rect 32826 1159 32827 1215
rect 32769 1147 32827 1159
rect 32865 3133 32923 3147
rect 32865 3081 32868 3133
rect 32920 3081 32923 3133
rect 32865 3069 32923 3081
rect 32865 3017 32868 3069
rect 32920 3017 32923 3069
rect 32865 3005 32923 3017
rect 32865 2953 32868 3005
rect 32920 2953 32923 3005
rect 32865 2941 32923 2953
rect 32865 2889 32868 2941
rect 32920 2889 32923 2941
rect 32865 2877 32923 2889
rect 32865 2825 32868 2877
rect 32920 2825 32923 2877
rect 32865 2813 32923 2825
rect 32865 2761 32868 2813
rect 32920 2761 32923 2813
rect 32865 2749 32923 2761
rect 32865 2697 32868 2749
rect 32920 2697 32923 2749
rect 32865 2685 32923 2697
rect 32865 2633 32868 2685
rect 32920 2633 32923 2685
rect 32865 2621 32923 2633
rect 32865 2569 32868 2621
rect 32920 2569 32923 2621
rect 32865 2557 32923 2569
rect 32865 2505 32868 2557
rect 32920 2505 32923 2557
rect 32865 2493 32923 2505
rect 32865 2441 32868 2493
rect 32920 2441 32923 2493
rect 32865 2429 32923 2441
rect 32865 2377 32868 2429
rect 32920 2377 32923 2429
rect 32865 2365 32923 2377
rect 32865 2313 32868 2365
rect 32920 2313 32923 2365
rect 32865 2301 32923 2313
rect 32865 2249 32868 2301
rect 32920 2249 32923 2301
rect 32865 2237 32923 2249
rect 32865 2185 32868 2237
rect 32920 2185 32923 2237
rect 32865 2173 32923 2185
rect 32865 2121 32868 2173
rect 32920 2121 32923 2173
rect 32865 2109 32923 2121
rect 32865 2057 32868 2109
rect 32920 2057 32923 2109
rect 32865 2045 32923 2057
rect 32865 1993 32868 2045
rect 32920 1993 32923 2045
rect 32865 1981 32923 1993
rect 32865 1929 32868 1981
rect 32920 1929 32923 1981
rect 32865 1917 32923 1929
rect 32865 1865 32868 1917
rect 32920 1865 32923 1917
rect 32865 1853 32923 1865
rect 32865 1801 32868 1853
rect 32920 1801 32923 1853
rect 32865 1789 32923 1801
rect 32865 1737 32868 1789
rect 32920 1737 32923 1789
rect 32865 1725 32923 1737
rect 32865 1673 32868 1725
rect 32920 1673 32923 1725
rect 32865 1661 32923 1673
rect 32865 1609 32868 1661
rect 32920 1609 32923 1661
rect 32865 1597 32923 1609
rect 32865 1545 32868 1597
rect 32920 1545 32923 1597
rect 32865 1533 32923 1545
rect 32865 1481 32868 1533
rect 32920 1481 32923 1533
rect 32865 1469 32923 1481
rect 32865 1417 32868 1469
rect 32920 1417 32923 1469
rect 32865 1405 32923 1417
rect 32865 1353 32868 1405
rect 32920 1353 32923 1405
rect 32865 1341 32923 1353
rect 32865 1289 32868 1341
rect 32920 1289 32923 1341
rect 32865 1277 32923 1289
rect 32865 1225 32868 1277
rect 32920 1225 32923 1277
rect 32865 1213 32923 1225
rect 32865 1161 32868 1213
rect 32920 1161 32923 1213
rect 32865 830 32923 1161
rect 32961 3135 33019 3147
rect 32961 3079 32962 3135
rect 33018 3079 33019 3135
rect 32961 3069 33019 3079
rect 32961 3055 32964 3069
rect 33016 3055 33019 3069
rect 32961 2999 32962 3055
rect 33018 2999 33019 3055
rect 32961 2975 32964 2999
rect 33016 2975 33019 2999
rect 32961 2919 32962 2975
rect 33018 2919 33019 2975
rect 32961 2895 32964 2919
rect 33016 2895 33019 2919
rect 32961 2839 32962 2895
rect 33018 2839 33019 2895
rect 32961 2825 32964 2839
rect 33016 2825 33019 2839
rect 32961 2815 33019 2825
rect 32961 2759 32962 2815
rect 33018 2759 33019 2815
rect 32961 2749 33019 2759
rect 32961 2735 32964 2749
rect 33016 2735 33019 2749
rect 32961 2679 32962 2735
rect 33018 2679 33019 2735
rect 32961 2655 32964 2679
rect 33016 2655 33019 2679
rect 32961 2599 32962 2655
rect 33018 2599 33019 2655
rect 32961 2575 32964 2599
rect 33016 2575 33019 2599
rect 32961 2519 32962 2575
rect 33018 2519 33019 2575
rect 32961 2505 32964 2519
rect 33016 2505 33019 2519
rect 32961 2495 33019 2505
rect 32961 2439 32962 2495
rect 33018 2439 33019 2495
rect 32961 2429 33019 2439
rect 32961 2415 32964 2429
rect 33016 2415 33019 2429
rect 32961 2359 32962 2415
rect 33018 2359 33019 2415
rect 32961 2335 32964 2359
rect 33016 2335 33019 2359
rect 32961 2279 32962 2335
rect 33018 2279 33019 2335
rect 32961 2255 32964 2279
rect 33016 2255 33019 2279
rect 32961 2199 32962 2255
rect 33018 2199 33019 2255
rect 32961 2185 32964 2199
rect 33016 2185 33019 2199
rect 32961 2175 33019 2185
rect 32961 2119 32962 2175
rect 33018 2119 33019 2175
rect 32961 2109 33019 2119
rect 32961 2095 32964 2109
rect 33016 2095 33019 2109
rect 32961 2039 32962 2095
rect 33018 2039 33019 2095
rect 32961 2015 32964 2039
rect 33016 2015 33019 2039
rect 32961 1959 32962 2015
rect 33018 1959 33019 2015
rect 32961 1935 32964 1959
rect 33016 1935 33019 1959
rect 32961 1879 32962 1935
rect 33018 1879 33019 1935
rect 32961 1865 32964 1879
rect 33016 1865 33019 1879
rect 32961 1855 33019 1865
rect 32961 1799 32962 1855
rect 33018 1799 33019 1855
rect 32961 1789 33019 1799
rect 32961 1775 32964 1789
rect 33016 1775 33019 1789
rect 32961 1719 32962 1775
rect 33018 1719 33019 1775
rect 32961 1695 32964 1719
rect 33016 1695 33019 1719
rect 32961 1639 32962 1695
rect 33018 1639 33019 1695
rect 32961 1615 32964 1639
rect 33016 1615 33019 1639
rect 32961 1559 32962 1615
rect 33018 1559 33019 1615
rect 32961 1545 32964 1559
rect 33016 1545 33019 1559
rect 32961 1535 33019 1545
rect 32961 1479 32962 1535
rect 33018 1479 33019 1535
rect 32961 1469 33019 1479
rect 32961 1455 32964 1469
rect 33016 1455 33019 1469
rect 32961 1399 32962 1455
rect 33018 1399 33019 1455
rect 32961 1375 32964 1399
rect 33016 1375 33019 1399
rect 32961 1319 32962 1375
rect 33018 1319 33019 1375
rect 32961 1295 32964 1319
rect 33016 1295 33019 1319
rect 32961 1239 32962 1295
rect 33018 1239 33019 1295
rect 32961 1225 32964 1239
rect 33016 1225 33019 1239
rect 32961 1215 33019 1225
rect 32961 1159 32962 1215
rect 33018 1159 33019 1215
rect 32961 1147 33019 1159
rect 33057 3133 33115 3147
rect 33057 3081 33060 3133
rect 33112 3081 33115 3133
rect 33057 3069 33115 3081
rect 33057 3017 33060 3069
rect 33112 3017 33115 3069
rect 33057 3005 33115 3017
rect 33057 2953 33060 3005
rect 33112 2953 33115 3005
rect 33057 2941 33115 2953
rect 33057 2889 33060 2941
rect 33112 2889 33115 2941
rect 33057 2877 33115 2889
rect 33057 2825 33060 2877
rect 33112 2825 33115 2877
rect 33057 2813 33115 2825
rect 33057 2761 33060 2813
rect 33112 2761 33115 2813
rect 33057 2749 33115 2761
rect 33057 2697 33060 2749
rect 33112 2697 33115 2749
rect 33057 2685 33115 2697
rect 33057 2633 33060 2685
rect 33112 2633 33115 2685
rect 33057 2621 33115 2633
rect 33057 2569 33060 2621
rect 33112 2569 33115 2621
rect 33057 2557 33115 2569
rect 33057 2505 33060 2557
rect 33112 2505 33115 2557
rect 33057 2493 33115 2505
rect 33057 2441 33060 2493
rect 33112 2441 33115 2493
rect 33057 2429 33115 2441
rect 33057 2377 33060 2429
rect 33112 2377 33115 2429
rect 33057 2365 33115 2377
rect 33057 2313 33060 2365
rect 33112 2313 33115 2365
rect 33057 2301 33115 2313
rect 33057 2249 33060 2301
rect 33112 2249 33115 2301
rect 33057 2237 33115 2249
rect 33057 2185 33060 2237
rect 33112 2185 33115 2237
rect 33057 2173 33115 2185
rect 33057 2121 33060 2173
rect 33112 2121 33115 2173
rect 33057 2109 33115 2121
rect 33057 2057 33060 2109
rect 33112 2057 33115 2109
rect 33057 2045 33115 2057
rect 33057 1993 33060 2045
rect 33112 1993 33115 2045
rect 33057 1981 33115 1993
rect 33057 1929 33060 1981
rect 33112 1929 33115 1981
rect 33057 1917 33115 1929
rect 33057 1865 33060 1917
rect 33112 1865 33115 1917
rect 33057 1853 33115 1865
rect 33057 1801 33060 1853
rect 33112 1801 33115 1853
rect 33057 1789 33115 1801
rect 33057 1737 33060 1789
rect 33112 1737 33115 1789
rect 33057 1725 33115 1737
rect 33057 1673 33060 1725
rect 33112 1673 33115 1725
rect 33057 1661 33115 1673
rect 33057 1609 33060 1661
rect 33112 1609 33115 1661
rect 33057 1597 33115 1609
rect 33057 1545 33060 1597
rect 33112 1545 33115 1597
rect 33057 1533 33115 1545
rect 33057 1481 33060 1533
rect 33112 1481 33115 1533
rect 33057 1469 33115 1481
rect 33057 1417 33060 1469
rect 33112 1417 33115 1469
rect 33057 1405 33115 1417
rect 33057 1353 33060 1405
rect 33112 1353 33115 1405
rect 33057 1341 33115 1353
rect 33057 1289 33060 1341
rect 33112 1289 33115 1341
rect 33057 1277 33115 1289
rect 33057 1225 33060 1277
rect 33112 1225 33115 1277
rect 33057 1213 33115 1225
rect 33057 1161 33060 1213
rect 33112 1161 33115 1213
rect 33057 830 33115 1161
rect 33153 3135 33211 3147
rect 33153 3079 33154 3135
rect 33210 3079 33211 3135
rect 33153 3069 33211 3079
rect 33153 3055 33156 3069
rect 33208 3055 33211 3069
rect 33153 2999 33154 3055
rect 33210 2999 33211 3055
rect 33153 2975 33156 2999
rect 33208 2975 33211 2999
rect 33153 2919 33154 2975
rect 33210 2919 33211 2975
rect 33153 2895 33156 2919
rect 33208 2895 33211 2919
rect 33153 2839 33154 2895
rect 33210 2839 33211 2895
rect 33153 2825 33156 2839
rect 33208 2825 33211 2839
rect 33153 2815 33211 2825
rect 33153 2759 33154 2815
rect 33210 2759 33211 2815
rect 33153 2749 33211 2759
rect 33153 2735 33156 2749
rect 33208 2735 33211 2749
rect 33153 2679 33154 2735
rect 33210 2679 33211 2735
rect 33153 2655 33156 2679
rect 33208 2655 33211 2679
rect 33153 2599 33154 2655
rect 33210 2599 33211 2655
rect 33153 2575 33156 2599
rect 33208 2575 33211 2599
rect 33153 2519 33154 2575
rect 33210 2519 33211 2575
rect 33153 2505 33156 2519
rect 33208 2505 33211 2519
rect 33153 2495 33211 2505
rect 33153 2439 33154 2495
rect 33210 2439 33211 2495
rect 33153 2429 33211 2439
rect 33153 2415 33156 2429
rect 33208 2415 33211 2429
rect 33153 2359 33154 2415
rect 33210 2359 33211 2415
rect 33153 2335 33156 2359
rect 33208 2335 33211 2359
rect 33153 2279 33154 2335
rect 33210 2279 33211 2335
rect 33153 2255 33156 2279
rect 33208 2255 33211 2279
rect 33153 2199 33154 2255
rect 33210 2199 33211 2255
rect 33153 2185 33156 2199
rect 33208 2185 33211 2199
rect 33153 2175 33211 2185
rect 33153 2119 33154 2175
rect 33210 2119 33211 2175
rect 33153 2109 33211 2119
rect 33153 2095 33156 2109
rect 33208 2095 33211 2109
rect 33153 2039 33154 2095
rect 33210 2039 33211 2095
rect 33153 2015 33156 2039
rect 33208 2015 33211 2039
rect 33153 1959 33154 2015
rect 33210 1959 33211 2015
rect 33153 1935 33156 1959
rect 33208 1935 33211 1959
rect 33153 1879 33154 1935
rect 33210 1879 33211 1935
rect 33153 1865 33156 1879
rect 33208 1865 33211 1879
rect 33153 1855 33211 1865
rect 33153 1799 33154 1855
rect 33210 1799 33211 1855
rect 33153 1789 33211 1799
rect 33153 1775 33156 1789
rect 33208 1775 33211 1789
rect 33153 1719 33154 1775
rect 33210 1719 33211 1775
rect 33153 1695 33156 1719
rect 33208 1695 33211 1719
rect 33153 1639 33154 1695
rect 33210 1639 33211 1695
rect 33153 1615 33156 1639
rect 33208 1615 33211 1639
rect 33153 1559 33154 1615
rect 33210 1559 33211 1615
rect 33153 1545 33156 1559
rect 33208 1545 33211 1559
rect 33153 1535 33211 1545
rect 33153 1479 33154 1535
rect 33210 1479 33211 1535
rect 33153 1469 33211 1479
rect 33153 1455 33156 1469
rect 33208 1455 33211 1469
rect 33153 1399 33154 1455
rect 33210 1399 33211 1455
rect 33153 1375 33156 1399
rect 33208 1375 33211 1399
rect 33153 1319 33154 1375
rect 33210 1319 33211 1375
rect 33153 1295 33156 1319
rect 33208 1295 33211 1319
rect 33153 1239 33154 1295
rect 33210 1239 33211 1295
rect 33153 1225 33156 1239
rect 33208 1225 33211 1239
rect 33153 1215 33211 1225
rect 33153 1159 33154 1215
rect 33210 1159 33211 1215
rect 33153 1147 33211 1159
rect 33249 3133 33307 3147
rect 33249 3081 33252 3133
rect 33304 3081 33307 3133
rect 33249 3069 33307 3081
rect 33249 3017 33252 3069
rect 33304 3017 33307 3069
rect 33249 3005 33307 3017
rect 33249 2953 33252 3005
rect 33304 2953 33307 3005
rect 33249 2941 33307 2953
rect 33249 2889 33252 2941
rect 33304 2889 33307 2941
rect 33249 2877 33307 2889
rect 33249 2825 33252 2877
rect 33304 2825 33307 2877
rect 33249 2813 33307 2825
rect 33249 2761 33252 2813
rect 33304 2761 33307 2813
rect 33249 2749 33307 2761
rect 33249 2697 33252 2749
rect 33304 2697 33307 2749
rect 33249 2685 33307 2697
rect 33249 2633 33252 2685
rect 33304 2633 33307 2685
rect 33249 2621 33307 2633
rect 33249 2569 33252 2621
rect 33304 2569 33307 2621
rect 33249 2557 33307 2569
rect 33249 2505 33252 2557
rect 33304 2505 33307 2557
rect 33249 2493 33307 2505
rect 33249 2441 33252 2493
rect 33304 2441 33307 2493
rect 33249 2429 33307 2441
rect 33249 2377 33252 2429
rect 33304 2377 33307 2429
rect 33249 2365 33307 2377
rect 33249 2313 33252 2365
rect 33304 2313 33307 2365
rect 33249 2301 33307 2313
rect 33249 2249 33252 2301
rect 33304 2249 33307 2301
rect 33249 2237 33307 2249
rect 33249 2185 33252 2237
rect 33304 2185 33307 2237
rect 33249 2173 33307 2185
rect 33249 2121 33252 2173
rect 33304 2121 33307 2173
rect 33249 2109 33307 2121
rect 33249 2057 33252 2109
rect 33304 2057 33307 2109
rect 33249 2045 33307 2057
rect 33249 1993 33252 2045
rect 33304 1993 33307 2045
rect 33249 1981 33307 1993
rect 33249 1929 33252 1981
rect 33304 1929 33307 1981
rect 33249 1917 33307 1929
rect 33249 1865 33252 1917
rect 33304 1865 33307 1917
rect 33249 1853 33307 1865
rect 33249 1801 33252 1853
rect 33304 1801 33307 1853
rect 33249 1789 33307 1801
rect 33249 1737 33252 1789
rect 33304 1737 33307 1789
rect 33249 1725 33307 1737
rect 33249 1673 33252 1725
rect 33304 1673 33307 1725
rect 33249 1661 33307 1673
rect 33249 1609 33252 1661
rect 33304 1609 33307 1661
rect 33249 1597 33307 1609
rect 33249 1545 33252 1597
rect 33304 1545 33307 1597
rect 33249 1533 33307 1545
rect 33249 1481 33252 1533
rect 33304 1481 33307 1533
rect 33249 1469 33307 1481
rect 33249 1417 33252 1469
rect 33304 1417 33307 1469
rect 33249 1405 33307 1417
rect 33249 1353 33252 1405
rect 33304 1353 33307 1405
rect 33249 1341 33307 1353
rect 33249 1289 33252 1341
rect 33304 1289 33307 1341
rect 33249 1277 33307 1289
rect 33249 1225 33252 1277
rect 33304 1225 33307 1277
rect 33249 1213 33307 1225
rect 33249 1161 33252 1213
rect 33304 1161 33307 1213
rect 33249 830 33307 1161
rect 33345 3135 33403 3147
rect 33345 3079 33346 3135
rect 33402 3079 33403 3135
rect 33345 3069 33403 3079
rect 33345 3055 33348 3069
rect 33400 3055 33403 3069
rect 33345 2999 33346 3055
rect 33402 2999 33403 3055
rect 33345 2975 33348 2999
rect 33400 2975 33403 2999
rect 33345 2919 33346 2975
rect 33402 2919 33403 2975
rect 33345 2895 33348 2919
rect 33400 2895 33403 2919
rect 33345 2839 33346 2895
rect 33402 2839 33403 2895
rect 33345 2825 33348 2839
rect 33400 2825 33403 2839
rect 33345 2815 33403 2825
rect 33345 2759 33346 2815
rect 33402 2759 33403 2815
rect 33345 2749 33403 2759
rect 33345 2735 33348 2749
rect 33400 2735 33403 2749
rect 33345 2679 33346 2735
rect 33402 2679 33403 2735
rect 33345 2655 33348 2679
rect 33400 2655 33403 2679
rect 33345 2599 33346 2655
rect 33402 2599 33403 2655
rect 33345 2575 33348 2599
rect 33400 2575 33403 2599
rect 33345 2519 33346 2575
rect 33402 2519 33403 2575
rect 33345 2505 33348 2519
rect 33400 2505 33403 2519
rect 33345 2495 33403 2505
rect 33345 2439 33346 2495
rect 33402 2439 33403 2495
rect 33345 2429 33403 2439
rect 33345 2415 33348 2429
rect 33400 2415 33403 2429
rect 33345 2359 33346 2415
rect 33402 2359 33403 2415
rect 33345 2335 33348 2359
rect 33400 2335 33403 2359
rect 33345 2279 33346 2335
rect 33402 2279 33403 2335
rect 33345 2255 33348 2279
rect 33400 2255 33403 2279
rect 33345 2199 33346 2255
rect 33402 2199 33403 2255
rect 33345 2185 33348 2199
rect 33400 2185 33403 2199
rect 33345 2175 33403 2185
rect 33345 2119 33346 2175
rect 33402 2119 33403 2175
rect 33345 2109 33403 2119
rect 33345 2095 33348 2109
rect 33400 2095 33403 2109
rect 33345 2039 33346 2095
rect 33402 2039 33403 2095
rect 33345 2015 33348 2039
rect 33400 2015 33403 2039
rect 33345 1959 33346 2015
rect 33402 1959 33403 2015
rect 33345 1935 33348 1959
rect 33400 1935 33403 1959
rect 33345 1879 33346 1935
rect 33402 1879 33403 1935
rect 33345 1865 33348 1879
rect 33400 1865 33403 1879
rect 33345 1855 33403 1865
rect 33345 1799 33346 1855
rect 33402 1799 33403 1855
rect 33345 1789 33403 1799
rect 33345 1775 33348 1789
rect 33400 1775 33403 1789
rect 33345 1719 33346 1775
rect 33402 1719 33403 1775
rect 33345 1695 33348 1719
rect 33400 1695 33403 1719
rect 33345 1639 33346 1695
rect 33402 1639 33403 1695
rect 33345 1615 33348 1639
rect 33400 1615 33403 1639
rect 33345 1559 33346 1615
rect 33402 1559 33403 1615
rect 33345 1545 33348 1559
rect 33400 1545 33403 1559
rect 33345 1535 33403 1545
rect 33345 1479 33346 1535
rect 33402 1479 33403 1535
rect 33345 1469 33403 1479
rect 33345 1455 33348 1469
rect 33400 1455 33403 1469
rect 33345 1399 33346 1455
rect 33402 1399 33403 1455
rect 33345 1375 33348 1399
rect 33400 1375 33403 1399
rect 33345 1319 33346 1375
rect 33402 1319 33403 1375
rect 33345 1295 33348 1319
rect 33400 1295 33403 1319
rect 33345 1239 33346 1295
rect 33402 1239 33403 1295
rect 33345 1225 33348 1239
rect 33400 1225 33403 1239
rect 33345 1215 33403 1225
rect 33345 1159 33346 1215
rect 33402 1159 33403 1215
rect 33345 1147 33403 1159
rect 33441 3133 33499 3147
rect 33441 3081 33444 3133
rect 33496 3081 33499 3133
rect 33441 3069 33499 3081
rect 33441 3017 33444 3069
rect 33496 3017 33499 3069
rect 33441 3005 33499 3017
rect 33441 2953 33444 3005
rect 33496 2953 33499 3005
rect 33441 2941 33499 2953
rect 33441 2889 33444 2941
rect 33496 2889 33499 2941
rect 33441 2877 33499 2889
rect 33441 2825 33444 2877
rect 33496 2825 33499 2877
rect 33441 2813 33499 2825
rect 33441 2761 33444 2813
rect 33496 2761 33499 2813
rect 33441 2749 33499 2761
rect 33441 2697 33444 2749
rect 33496 2697 33499 2749
rect 33441 2685 33499 2697
rect 33441 2633 33444 2685
rect 33496 2633 33499 2685
rect 33441 2621 33499 2633
rect 33441 2569 33444 2621
rect 33496 2569 33499 2621
rect 33441 2557 33499 2569
rect 33441 2505 33444 2557
rect 33496 2505 33499 2557
rect 33441 2493 33499 2505
rect 33441 2441 33444 2493
rect 33496 2441 33499 2493
rect 33441 2429 33499 2441
rect 33441 2377 33444 2429
rect 33496 2377 33499 2429
rect 33441 2365 33499 2377
rect 33441 2313 33444 2365
rect 33496 2313 33499 2365
rect 33441 2301 33499 2313
rect 33441 2249 33444 2301
rect 33496 2249 33499 2301
rect 33441 2237 33499 2249
rect 33441 2185 33444 2237
rect 33496 2185 33499 2237
rect 33441 2173 33499 2185
rect 33441 2121 33444 2173
rect 33496 2121 33499 2173
rect 33441 2109 33499 2121
rect 33441 2057 33444 2109
rect 33496 2057 33499 2109
rect 33441 2045 33499 2057
rect 33441 1993 33444 2045
rect 33496 1993 33499 2045
rect 33441 1981 33499 1993
rect 33441 1929 33444 1981
rect 33496 1929 33499 1981
rect 33441 1917 33499 1929
rect 33441 1865 33444 1917
rect 33496 1865 33499 1917
rect 33441 1853 33499 1865
rect 33441 1801 33444 1853
rect 33496 1801 33499 1853
rect 33441 1789 33499 1801
rect 33441 1737 33444 1789
rect 33496 1737 33499 1789
rect 33441 1725 33499 1737
rect 33441 1673 33444 1725
rect 33496 1673 33499 1725
rect 33441 1661 33499 1673
rect 33441 1609 33444 1661
rect 33496 1609 33499 1661
rect 33441 1597 33499 1609
rect 33441 1545 33444 1597
rect 33496 1545 33499 1597
rect 33441 1533 33499 1545
rect 33441 1481 33444 1533
rect 33496 1481 33499 1533
rect 33441 1469 33499 1481
rect 33441 1417 33444 1469
rect 33496 1417 33499 1469
rect 33441 1405 33499 1417
rect 33441 1353 33444 1405
rect 33496 1353 33499 1405
rect 33441 1341 33499 1353
rect 33441 1289 33444 1341
rect 33496 1289 33499 1341
rect 33441 1277 33499 1289
rect 33441 1225 33444 1277
rect 33496 1225 33499 1277
rect 33441 1213 33499 1225
rect 33441 1161 33444 1213
rect 33496 1161 33499 1213
rect 33441 830 33499 1161
rect 33537 3135 33595 3147
rect 33537 3079 33538 3135
rect 33594 3079 33595 3135
rect 33537 3069 33595 3079
rect 33537 3055 33540 3069
rect 33592 3055 33595 3069
rect 33537 2999 33538 3055
rect 33594 2999 33595 3055
rect 33537 2975 33540 2999
rect 33592 2975 33595 2999
rect 33537 2919 33538 2975
rect 33594 2919 33595 2975
rect 33537 2895 33540 2919
rect 33592 2895 33595 2919
rect 33537 2839 33538 2895
rect 33594 2839 33595 2895
rect 33537 2825 33540 2839
rect 33592 2825 33595 2839
rect 33537 2815 33595 2825
rect 33537 2759 33538 2815
rect 33594 2759 33595 2815
rect 33537 2749 33595 2759
rect 33537 2735 33540 2749
rect 33592 2735 33595 2749
rect 33537 2679 33538 2735
rect 33594 2679 33595 2735
rect 33537 2655 33540 2679
rect 33592 2655 33595 2679
rect 33537 2599 33538 2655
rect 33594 2599 33595 2655
rect 33537 2575 33540 2599
rect 33592 2575 33595 2599
rect 33537 2519 33538 2575
rect 33594 2519 33595 2575
rect 33537 2505 33540 2519
rect 33592 2505 33595 2519
rect 33537 2495 33595 2505
rect 33537 2439 33538 2495
rect 33594 2439 33595 2495
rect 33537 2429 33595 2439
rect 33537 2415 33540 2429
rect 33592 2415 33595 2429
rect 33537 2359 33538 2415
rect 33594 2359 33595 2415
rect 33537 2335 33540 2359
rect 33592 2335 33595 2359
rect 33537 2279 33538 2335
rect 33594 2279 33595 2335
rect 33537 2255 33540 2279
rect 33592 2255 33595 2279
rect 33537 2199 33538 2255
rect 33594 2199 33595 2255
rect 33537 2185 33540 2199
rect 33592 2185 33595 2199
rect 33537 2175 33595 2185
rect 33537 2119 33538 2175
rect 33594 2119 33595 2175
rect 33537 2109 33595 2119
rect 33537 2095 33540 2109
rect 33592 2095 33595 2109
rect 33537 2039 33538 2095
rect 33594 2039 33595 2095
rect 33537 2015 33540 2039
rect 33592 2015 33595 2039
rect 33537 1959 33538 2015
rect 33594 1959 33595 2015
rect 33537 1935 33540 1959
rect 33592 1935 33595 1959
rect 33537 1879 33538 1935
rect 33594 1879 33595 1935
rect 33537 1865 33540 1879
rect 33592 1865 33595 1879
rect 33537 1855 33595 1865
rect 33537 1799 33538 1855
rect 33594 1799 33595 1855
rect 33537 1789 33595 1799
rect 33537 1775 33540 1789
rect 33592 1775 33595 1789
rect 33537 1719 33538 1775
rect 33594 1719 33595 1775
rect 33537 1695 33540 1719
rect 33592 1695 33595 1719
rect 33537 1639 33538 1695
rect 33594 1639 33595 1695
rect 33537 1615 33540 1639
rect 33592 1615 33595 1639
rect 33537 1559 33538 1615
rect 33594 1559 33595 1615
rect 33537 1545 33540 1559
rect 33592 1545 33595 1559
rect 33537 1535 33595 1545
rect 33537 1479 33538 1535
rect 33594 1479 33595 1535
rect 33537 1469 33595 1479
rect 33537 1455 33540 1469
rect 33592 1455 33595 1469
rect 33537 1399 33538 1455
rect 33594 1399 33595 1455
rect 33537 1375 33540 1399
rect 33592 1375 33595 1399
rect 33537 1319 33538 1375
rect 33594 1319 33595 1375
rect 33537 1295 33540 1319
rect 33592 1295 33595 1319
rect 33537 1239 33538 1295
rect 33594 1239 33595 1295
rect 33537 1225 33540 1239
rect 33592 1225 33595 1239
rect 33537 1215 33595 1225
rect 33537 1159 33538 1215
rect 33594 1159 33595 1215
rect 33537 1147 33595 1159
rect 33633 3133 33691 3147
rect 33633 3081 33636 3133
rect 33688 3081 33691 3133
rect 33633 3069 33691 3081
rect 33633 3017 33636 3069
rect 33688 3017 33691 3069
rect 33633 3005 33691 3017
rect 33633 2953 33636 3005
rect 33688 2953 33691 3005
rect 33633 2941 33691 2953
rect 33633 2889 33636 2941
rect 33688 2889 33691 2941
rect 33633 2877 33691 2889
rect 33633 2825 33636 2877
rect 33688 2825 33691 2877
rect 33633 2813 33691 2825
rect 33633 2761 33636 2813
rect 33688 2761 33691 2813
rect 33633 2749 33691 2761
rect 33633 2697 33636 2749
rect 33688 2697 33691 2749
rect 33633 2685 33691 2697
rect 33633 2633 33636 2685
rect 33688 2633 33691 2685
rect 33633 2621 33691 2633
rect 33633 2569 33636 2621
rect 33688 2569 33691 2621
rect 33633 2557 33691 2569
rect 33633 2505 33636 2557
rect 33688 2505 33691 2557
rect 33633 2493 33691 2505
rect 33633 2441 33636 2493
rect 33688 2441 33691 2493
rect 33633 2429 33691 2441
rect 33633 2377 33636 2429
rect 33688 2377 33691 2429
rect 33633 2365 33691 2377
rect 33633 2313 33636 2365
rect 33688 2313 33691 2365
rect 33633 2301 33691 2313
rect 33633 2249 33636 2301
rect 33688 2249 33691 2301
rect 33633 2237 33691 2249
rect 33633 2185 33636 2237
rect 33688 2185 33691 2237
rect 33633 2173 33691 2185
rect 33633 2121 33636 2173
rect 33688 2121 33691 2173
rect 33633 2109 33691 2121
rect 33633 2057 33636 2109
rect 33688 2057 33691 2109
rect 33633 2045 33691 2057
rect 33633 1993 33636 2045
rect 33688 1993 33691 2045
rect 33633 1981 33691 1993
rect 33633 1929 33636 1981
rect 33688 1929 33691 1981
rect 33633 1917 33691 1929
rect 33633 1865 33636 1917
rect 33688 1865 33691 1917
rect 33633 1853 33691 1865
rect 33633 1801 33636 1853
rect 33688 1801 33691 1853
rect 33633 1789 33691 1801
rect 33633 1737 33636 1789
rect 33688 1737 33691 1789
rect 33633 1725 33691 1737
rect 33633 1673 33636 1725
rect 33688 1673 33691 1725
rect 33633 1661 33691 1673
rect 33633 1609 33636 1661
rect 33688 1609 33691 1661
rect 33633 1597 33691 1609
rect 33633 1545 33636 1597
rect 33688 1545 33691 1597
rect 33633 1533 33691 1545
rect 33633 1481 33636 1533
rect 33688 1481 33691 1533
rect 33633 1469 33691 1481
rect 33633 1417 33636 1469
rect 33688 1417 33691 1469
rect 33633 1405 33691 1417
rect 33633 1353 33636 1405
rect 33688 1353 33691 1405
rect 33633 1341 33691 1353
rect 33633 1289 33636 1341
rect 33688 1289 33691 1341
rect 33633 1277 33691 1289
rect 33633 1225 33636 1277
rect 33688 1225 33691 1277
rect 33633 1213 33691 1225
rect 33633 1161 33636 1213
rect 33688 1161 33691 1213
rect 33633 830 33691 1161
rect 33729 3135 33787 3147
rect 33729 3079 33730 3135
rect 33786 3079 33787 3135
rect 33729 3069 33787 3079
rect 33729 3055 33732 3069
rect 33784 3055 33787 3069
rect 33729 2999 33730 3055
rect 33786 2999 33787 3055
rect 33729 2975 33732 2999
rect 33784 2975 33787 2999
rect 33729 2919 33730 2975
rect 33786 2919 33787 2975
rect 33729 2895 33732 2919
rect 33784 2895 33787 2919
rect 33729 2839 33730 2895
rect 33786 2839 33787 2895
rect 33729 2825 33732 2839
rect 33784 2825 33787 2839
rect 33729 2815 33787 2825
rect 33729 2759 33730 2815
rect 33786 2759 33787 2815
rect 33729 2749 33787 2759
rect 33729 2735 33732 2749
rect 33784 2735 33787 2749
rect 33729 2679 33730 2735
rect 33786 2679 33787 2735
rect 33729 2655 33732 2679
rect 33784 2655 33787 2679
rect 33729 2599 33730 2655
rect 33786 2599 33787 2655
rect 33729 2575 33732 2599
rect 33784 2575 33787 2599
rect 33729 2519 33730 2575
rect 33786 2519 33787 2575
rect 33729 2505 33732 2519
rect 33784 2505 33787 2519
rect 33729 2495 33787 2505
rect 33729 2439 33730 2495
rect 33786 2439 33787 2495
rect 33729 2429 33787 2439
rect 33729 2415 33732 2429
rect 33784 2415 33787 2429
rect 33729 2359 33730 2415
rect 33786 2359 33787 2415
rect 33729 2335 33732 2359
rect 33784 2335 33787 2359
rect 33729 2279 33730 2335
rect 33786 2279 33787 2335
rect 33729 2255 33732 2279
rect 33784 2255 33787 2279
rect 33729 2199 33730 2255
rect 33786 2199 33787 2255
rect 33729 2185 33732 2199
rect 33784 2185 33787 2199
rect 33729 2175 33787 2185
rect 33729 2119 33730 2175
rect 33786 2119 33787 2175
rect 33729 2109 33787 2119
rect 33729 2095 33732 2109
rect 33784 2095 33787 2109
rect 33729 2039 33730 2095
rect 33786 2039 33787 2095
rect 33729 2015 33732 2039
rect 33784 2015 33787 2039
rect 33729 1959 33730 2015
rect 33786 1959 33787 2015
rect 33729 1935 33732 1959
rect 33784 1935 33787 1959
rect 33729 1879 33730 1935
rect 33786 1879 33787 1935
rect 33729 1865 33732 1879
rect 33784 1865 33787 1879
rect 33729 1855 33787 1865
rect 33729 1799 33730 1855
rect 33786 1799 33787 1855
rect 33729 1789 33787 1799
rect 33729 1775 33732 1789
rect 33784 1775 33787 1789
rect 33729 1719 33730 1775
rect 33786 1719 33787 1775
rect 33729 1695 33732 1719
rect 33784 1695 33787 1719
rect 33729 1639 33730 1695
rect 33786 1639 33787 1695
rect 33729 1615 33732 1639
rect 33784 1615 33787 1639
rect 33729 1559 33730 1615
rect 33786 1559 33787 1615
rect 33729 1545 33732 1559
rect 33784 1545 33787 1559
rect 33729 1535 33787 1545
rect 33729 1479 33730 1535
rect 33786 1479 33787 1535
rect 33729 1469 33787 1479
rect 33729 1455 33732 1469
rect 33784 1455 33787 1469
rect 33729 1399 33730 1455
rect 33786 1399 33787 1455
rect 33729 1375 33732 1399
rect 33784 1375 33787 1399
rect 33729 1319 33730 1375
rect 33786 1319 33787 1375
rect 33729 1295 33732 1319
rect 33784 1295 33787 1319
rect 33729 1239 33730 1295
rect 33786 1239 33787 1295
rect 33729 1225 33732 1239
rect 33784 1225 33787 1239
rect 33729 1215 33787 1225
rect 33729 1159 33730 1215
rect 33786 1159 33787 1215
rect 33729 1147 33787 1159
rect 33825 3133 33883 3147
rect 33825 3081 33828 3133
rect 33880 3081 33883 3133
rect 33825 3069 33883 3081
rect 33825 3017 33828 3069
rect 33880 3017 33883 3069
rect 33825 3005 33883 3017
rect 33825 2953 33828 3005
rect 33880 2953 33883 3005
rect 33825 2941 33883 2953
rect 33825 2889 33828 2941
rect 33880 2889 33883 2941
rect 33825 2877 33883 2889
rect 33825 2825 33828 2877
rect 33880 2825 33883 2877
rect 33825 2813 33883 2825
rect 33825 2761 33828 2813
rect 33880 2761 33883 2813
rect 33825 2749 33883 2761
rect 33825 2697 33828 2749
rect 33880 2697 33883 2749
rect 33825 2685 33883 2697
rect 33825 2633 33828 2685
rect 33880 2633 33883 2685
rect 33825 2621 33883 2633
rect 33825 2569 33828 2621
rect 33880 2569 33883 2621
rect 33825 2557 33883 2569
rect 33825 2505 33828 2557
rect 33880 2505 33883 2557
rect 33825 2493 33883 2505
rect 33825 2441 33828 2493
rect 33880 2441 33883 2493
rect 33825 2429 33883 2441
rect 33825 2377 33828 2429
rect 33880 2377 33883 2429
rect 33825 2365 33883 2377
rect 33825 2313 33828 2365
rect 33880 2313 33883 2365
rect 33825 2301 33883 2313
rect 33825 2249 33828 2301
rect 33880 2249 33883 2301
rect 33825 2237 33883 2249
rect 33825 2185 33828 2237
rect 33880 2185 33883 2237
rect 33825 2173 33883 2185
rect 33825 2121 33828 2173
rect 33880 2121 33883 2173
rect 33825 2109 33883 2121
rect 33825 2057 33828 2109
rect 33880 2057 33883 2109
rect 33825 2045 33883 2057
rect 33825 1993 33828 2045
rect 33880 1993 33883 2045
rect 33825 1981 33883 1993
rect 33825 1929 33828 1981
rect 33880 1929 33883 1981
rect 33825 1917 33883 1929
rect 33825 1865 33828 1917
rect 33880 1865 33883 1917
rect 33825 1853 33883 1865
rect 33825 1801 33828 1853
rect 33880 1801 33883 1853
rect 33825 1789 33883 1801
rect 33825 1737 33828 1789
rect 33880 1737 33883 1789
rect 33825 1725 33883 1737
rect 33825 1673 33828 1725
rect 33880 1673 33883 1725
rect 33825 1661 33883 1673
rect 33825 1609 33828 1661
rect 33880 1609 33883 1661
rect 33825 1597 33883 1609
rect 33825 1545 33828 1597
rect 33880 1545 33883 1597
rect 33825 1533 33883 1545
rect 33825 1481 33828 1533
rect 33880 1481 33883 1533
rect 33825 1469 33883 1481
rect 33825 1417 33828 1469
rect 33880 1417 33883 1469
rect 33825 1405 33883 1417
rect 33825 1353 33828 1405
rect 33880 1353 33883 1405
rect 33825 1341 33883 1353
rect 33825 1289 33828 1341
rect 33880 1289 33883 1341
rect 33825 1277 33883 1289
rect 33825 1225 33828 1277
rect 33880 1225 33883 1277
rect 33825 1213 33883 1225
rect 33825 1161 33828 1213
rect 33880 1161 33883 1213
rect 33825 830 33883 1161
rect 33921 3135 33979 3147
rect 33921 3079 33922 3135
rect 33978 3079 33979 3135
rect 33921 3069 33979 3079
rect 33921 3055 33924 3069
rect 33976 3055 33979 3069
rect 33921 2999 33922 3055
rect 33978 2999 33979 3055
rect 33921 2975 33924 2999
rect 33976 2975 33979 2999
rect 33921 2919 33922 2975
rect 33978 2919 33979 2975
rect 33921 2895 33924 2919
rect 33976 2895 33979 2919
rect 33921 2839 33922 2895
rect 33978 2839 33979 2895
rect 33921 2825 33924 2839
rect 33976 2825 33979 2839
rect 33921 2815 33979 2825
rect 33921 2759 33922 2815
rect 33978 2759 33979 2815
rect 33921 2749 33979 2759
rect 33921 2735 33924 2749
rect 33976 2735 33979 2749
rect 33921 2679 33922 2735
rect 33978 2679 33979 2735
rect 33921 2655 33924 2679
rect 33976 2655 33979 2679
rect 33921 2599 33922 2655
rect 33978 2599 33979 2655
rect 33921 2575 33924 2599
rect 33976 2575 33979 2599
rect 33921 2519 33922 2575
rect 33978 2519 33979 2575
rect 33921 2505 33924 2519
rect 33976 2505 33979 2519
rect 33921 2495 33979 2505
rect 33921 2439 33922 2495
rect 33978 2439 33979 2495
rect 33921 2429 33979 2439
rect 33921 2415 33924 2429
rect 33976 2415 33979 2429
rect 33921 2359 33922 2415
rect 33978 2359 33979 2415
rect 33921 2335 33924 2359
rect 33976 2335 33979 2359
rect 33921 2279 33922 2335
rect 33978 2279 33979 2335
rect 33921 2255 33924 2279
rect 33976 2255 33979 2279
rect 33921 2199 33922 2255
rect 33978 2199 33979 2255
rect 33921 2185 33924 2199
rect 33976 2185 33979 2199
rect 33921 2175 33979 2185
rect 33921 2119 33922 2175
rect 33978 2119 33979 2175
rect 33921 2109 33979 2119
rect 33921 2095 33924 2109
rect 33976 2095 33979 2109
rect 33921 2039 33922 2095
rect 33978 2039 33979 2095
rect 33921 2015 33924 2039
rect 33976 2015 33979 2039
rect 33921 1959 33922 2015
rect 33978 1959 33979 2015
rect 33921 1935 33924 1959
rect 33976 1935 33979 1959
rect 33921 1879 33922 1935
rect 33978 1879 33979 1935
rect 33921 1865 33924 1879
rect 33976 1865 33979 1879
rect 33921 1855 33979 1865
rect 33921 1799 33922 1855
rect 33978 1799 33979 1855
rect 33921 1789 33979 1799
rect 33921 1775 33924 1789
rect 33976 1775 33979 1789
rect 33921 1719 33922 1775
rect 33978 1719 33979 1775
rect 33921 1695 33924 1719
rect 33976 1695 33979 1719
rect 33921 1639 33922 1695
rect 33978 1639 33979 1695
rect 33921 1615 33924 1639
rect 33976 1615 33979 1639
rect 33921 1559 33922 1615
rect 33978 1559 33979 1615
rect 33921 1545 33924 1559
rect 33976 1545 33979 1559
rect 33921 1535 33979 1545
rect 33921 1479 33922 1535
rect 33978 1479 33979 1535
rect 33921 1469 33979 1479
rect 33921 1455 33924 1469
rect 33976 1455 33979 1469
rect 33921 1399 33922 1455
rect 33978 1399 33979 1455
rect 33921 1375 33924 1399
rect 33976 1375 33979 1399
rect 33921 1319 33922 1375
rect 33978 1319 33979 1375
rect 33921 1295 33924 1319
rect 33976 1295 33979 1319
rect 33921 1239 33922 1295
rect 33978 1239 33979 1295
rect 33921 1225 33924 1239
rect 33976 1225 33979 1239
rect 33921 1215 33979 1225
rect 33921 1159 33922 1215
rect 33978 1159 33979 1215
rect 33921 1147 33979 1159
rect 34017 3133 34075 3147
rect 34017 3081 34020 3133
rect 34072 3081 34075 3133
rect 34017 3069 34075 3081
rect 34017 3017 34020 3069
rect 34072 3017 34075 3069
rect 34017 3005 34075 3017
rect 34017 2953 34020 3005
rect 34072 2953 34075 3005
rect 34017 2941 34075 2953
rect 34017 2889 34020 2941
rect 34072 2889 34075 2941
rect 34017 2877 34075 2889
rect 34017 2825 34020 2877
rect 34072 2825 34075 2877
rect 34017 2813 34075 2825
rect 34017 2761 34020 2813
rect 34072 2761 34075 2813
rect 34017 2749 34075 2761
rect 34017 2697 34020 2749
rect 34072 2697 34075 2749
rect 34017 2685 34075 2697
rect 34017 2633 34020 2685
rect 34072 2633 34075 2685
rect 34017 2621 34075 2633
rect 34017 2569 34020 2621
rect 34072 2569 34075 2621
rect 34017 2557 34075 2569
rect 34017 2505 34020 2557
rect 34072 2505 34075 2557
rect 34017 2493 34075 2505
rect 34017 2441 34020 2493
rect 34072 2441 34075 2493
rect 34017 2429 34075 2441
rect 34017 2377 34020 2429
rect 34072 2377 34075 2429
rect 34017 2365 34075 2377
rect 34017 2313 34020 2365
rect 34072 2313 34075 2365
rect 34017 2301 34075 2313
rect 34017 2249 34020 2301
rect 34072 2249 34075 2301
rect 34017 2237 34075 2249
rect 34017 2185 34020 2237
rect 34072 2185 34075 2237
rect 34017 2173 34075 2185
rect 34017 2121 34020 2173
rect 34072 2121 34075 2173
rect 34017 2109 34075 2121
rect 34017 2057 34020 2109
rect 34072 2057 34075 2109
rect 34017 2045 34075 2057
rect 34017 1993 34020 2045
rect 34072 1993 34075 2045
rect 34017 1981 34075 1993
rect 34017 1929 34020 1981
rect 34072 1929 34075 1981
rect 34017 1917 34075 1929
rect 34017 1865 34020 1917
rect 34072 1865 34075 1917
rect 34017 1853 34075 1865
rect 34017 1801 34020 1853
rect 34072 1801 34075 1853
rect 34017 1789 34075 1801
rect 34017 1737 34020 1789
rect 34072 1737 34075 1789
rect 34017 1725 34075 1737
rect 34017 1673 34020 1725
rect 34072 1673 34075 1725
rect 34017 1661 34075 1673
rect 34017 1609 34020 1661
rect 34072 1609 34075 1661
rect 34017 1597 34075 1609
rect 34017 1545 34020 1597
rect 34072 1545 34075 1597
rect 34017 1533 34075 1545
rect 34017 1481 34020 1533
rect 34072 1481 34075 1533
rect 34017 1469 34075 1481
rect 34017 1417 34020 1469
rect 34072 1417 34075 1469
rect 34017 1405 34075 1417
rect 34017 1353 34020 1405
rect 34072 1353 34075 1405
rect 34017 1341 34075 1353
rect 34017 1289 34020 1341
rect 34072 1289 34075 1341
rect 34017 1277 34075 1289
rect 34017 1225 34020 1277
rect 34072 1225 34075 1277
rect 34017 1213 34075 1225
rect 34017 1161 34020 1213
rect 34072 1161 34075 1213
rect 34017 830 34075 1161
rect 34113 3135 34171 3147
rect 34113 3079 34114 3135
rect 34170 3079 34171 3135
rect 34113 3069 34171 3079
rect 34113 3055 34116 3069
rect 34168 3055 34171 3069
rect 34113 2999 34114 3055
rect 34170 2999 34171 3055
rect 34113 2975 34116 2999
rect 34168 2975 34171 2999
rect 34113 2919 34114 2975
rect 34170 2919 34171 2975
rect 34113 2895 34116 2919
rect 34168 2895 34171 2919
rect 34113 2839 34114 2895
rect 34170 2839 34171 2895
rect 34113 2825 34116 2839
rect 34168 2825 34171 2839
rect 34113 2815 34171 2825
rect 34113 2759 34114 2815
rect 34170 2759 34171 2815
rect 34113 2749 34171 2759
rect 34113 2735 34116 2749
rect 34168 2735 34171 2749
rect 34113 2679 34114 2735
rect 34170 2679 34171 2735
rect 34113 2655 34116 2679
rect 34168 2655 34171 2679
rect 34113 2599 34114 2655
rect 34170 2599 34171 2655
rect 34113 2575 34116 2599
rect 34168 2575 34171 2599
rect 34113 2519 34114 2575
rect 34170 2519 34171 2575
rect 34113 2505 34116 2519
rect 34168 2505 34171 2519
rect 34113 2495 34171 2505
rect 34113 2439 34114 2495
rect 34170 2439 34171 2495
rect 34113 2429 34171 2439
rect 34113 2415 34116 2429
rect 34168 2415 34171 2429
rect 34113 2359 34114 2415
rect 34170 2359 34171 2415
rect 34113 2335 34116 2359
rect 34168 2335 34171 2359
rect 34113 2279 34114 2335
rect 34170 2279 34171 2335
rect 34113 2255 34116 2279
rect 34168 2255 34171 2279
rect 34113 2199 34114 2255
rect 34170 2199 34171 2255
rect 34113 2185 34116 2199
rect 34168 2185 34171 2199
rect 34113 2175 34171 2185
rect 34113 2119 34114 2175
rect 34170 2119 34171 2175
rect 34113 2109 34171 2119
rect 34113 2095 34116 2109
rect 34168 2095 34171 2109
rect 34113 2039 34114 2095
rect 34170 2039 34171 2095
rect 34113 2015 34116 2039
rect 34168 2015 34171 2039
rect 34113 1959 34114 2015
rect 34170 1959 34171 2015
rect 34113 1935 34116 1959
rect 34168 1935 34171 1959
rect 34113 1879 34114 1935
rect 34170 1879 34171 1935
rect 34113 1865 34116 1879
rect 34168 1865 34171 1879
rect 34113 1855 34171 1865
rect 34113 1799 34114 1855
rect 34170 1799 34171 1855
rect 34113 1789 34171 1799
rect 34113 1775 34116 1789
rect 34168 1775 34171 1789
rect 34113 1719 34114 1775
rect 34170 1719 34171 1775
rect 34113 1695 34116 1719
rect 34168 1695 34171 1719
rect 34113 1639 34114 1695
rect 34170 1639 34171 1695
rect 34113 1615 34116 1639
rect 34168 1615 34171 1639
rect 34113 1559 34114 1615
rect 34170 1559 34171 1615
rect 34113 1545 34116 1559
rect 34168 1545 34171 1559
rect 34113 1535 34171 1545
rect 34113 1479 34114 1535
rect 34170 1479 34171 1535
rect 34113 1469 34171 1479
rect 34113 1455 34116 1469
rect 34168 1455 34171 1469
rect 34113 1399 34114 1455
rect 34170 1399 34171 1455
rect 34113 1375 34116 1399
rect 34168 1375 34171 1399
rect 34113 1319 34114 1375
rect 34170 1319 34171 1375
rect 34113 1295 34116 1319
rect 34168 1295 34171 1319
rect 34113 1239 34114 1295
rect 34170 1239 34171 1295
rect 34113 1225 34116 1239
rect 34168 1225 34171 1239
rect 34113 1215 34171 1225
rect 34113 1159 34114 1215
rect 34170 1159 34171 1215
rect 34113 1147 34171 1159
rect 34209 3133 34267 3147
rect 34209 3081 34212 3133
rect 34264 3081 34267 3133
rect 34209 3069 34267 3081
rect 34209 3017 34212 3069
rect 34264 3017 34267 3069
rect 34209 3005 34267 3017
rect 34209 2953 34212 3005
rect 34264 2953 34267 3005
rect 34209 2941 34267 2953
rect 34209 2889 34212 2941
rect 34264 2889 34267 2941
rect 34209 2877 34267 2889
rect 34209 2825 34212 2877
rect 34264 2825 34267 2877
rect 34209 2813 34267 2825
rect 34209 2761 34212 2813
rect 34264 2761 34267 2813
rect 34209 2749 34267 2761
rect 34209 2697 34212 2749
rect 34264 2697 34267 2749
rect 34209 2685 34267 2697
rect 34209 2633 34212 2685
rect 34264 2633 34267 2685
rect 34209 2621 34267 2633
rect 34209 2569 34212 2621
rect 34264 2569 34267 2621
rect 34209 2557 34267 2569
rect 34209 2505 34212 2557
rect 34264 2505 34267 2557
rect 34209 2493 34267 2505
rect 34209 2441 34212 2493
rect 34264 2441 34267 2493
rect 34209 2429 34267 2441
rect 34209 2377 34212 2429
rect 34264 2377 34267 2429
rect 34209 2365 34267 2377
rect 34209 2313 34212 2365
rect 34264 2313 34267 2365
rect 34209 2301 34267 2313
rect 34209 2249 34212 2301
rect 34264 2249 34267 2301
rect 34209 2237 34267 2249
rect 34209 2185 34212 2237
rect 34264 2185 34267 2237
rect 34209 2173 34267 2185
rect 34209 2121 34212 2173
rect 34264 2121 34267 2173
rect 34209 2109 34267 2121
rect 34209 2057 34212 2109
rect 34264 2057 34267 2109
rect 34209 2045 34267 2057
rect 34209 1993 34212 2045
rect 34264 1993 34267 2045
rect 34209 1981 34267 1993
rect 34209 1929 34212 1981
rect 34264 1929 34267 1981
rect 34209 1917 34267 1929
rect 34209 1865 34212 1917
rect 34264 1865 34267 1917
rect 34209 1853 34267 1865
rect 34209 1801 34212 1853
rect 34264 1801 34267 1853
rect 34209 1789 34267 1801
rect 34209 1737 34212 1789
rect 34264 1737 34267 1789
rect 34209 1725 34267 1737
rect 34209 1673 34212 1725
rect 34264 1673 34267 1725
rect 34209 1661 34267 1673
rect 34209 1609 34212 1661
rect 34264 1609 34267 1661
rect 34209 1597 34267 1609
rect 34209 1545 34212 1597
rect 34264 1545 34267 1597
rect 34209 1533 34267 1545
rect 34209 1481 34212 1533
rect 34264 1481 34267 1533
rect 34209 1469 34267 1481
rect 34209 1417 34212 1469
rect 34264 1417 34267 1469
rect 34209 1405 34267 1417
rect 34209 1353 34212 1405
rect 34264 1353 34267 1405
rect 34209 1341 34267 1353
rect 34209 1289 34212 1341
rect 34264 1289 34267 1341
rect 34209 1277 34267 1289
rect 34209 1225 34212 1277
rect 34264 1225 34267 1277
rect 34209 1213 34267 1225
rect 34209 1161 34212 1213
rect 34264 1161 34267 1213
rect 34209 830 34267 1161
rect 34305 3135 34363 3147
rect 34305 3079 34306 3135
rect 34362 3079 34363 3135
rect 34305 3069 34363 3079
rect 34305 3055 34308 3069
rect 34360 3055 34363 3069
rect 34305 2999 34306 3055
rect 34362 2999 34363 3055
rect 34305 2975 34308 2999
rect 34360 2975 34363 2999
rect 34305 2919 34306 2975
rect 34362 2919 34363 2975
rect 34305 2895 34308 2919
rect 34360 2895 34363 2919
rect 34305 2839 34306 2895
rect 34362 2839 34363 2895
rect 34305 2825 34308 2839
rect 34360 2825 34363 2839
rect 34305 2815 34363 2825
rect 34305 2759 34306 2815
rect 34362 2759 34363 2815
rect 34305 2749 34363 2759
rect 34305 2735 34308 2749
rect 34360 2735 34363 2749
rect 34305 2679 34306 2735
rect 34362 2679 34363 2735
rect 34305 2655 34308 2679
rect 34360 2655 34363 2679
rect 34305 2599 34306 2655
rect 34362 2599 34363 2655
rect 34305 2575 34308 2599
rect 34360 2575 34363 2599
rect 34305 2519 34306 2575
rect 34362 2519 34363 2575
rect 34305 2505 34308 2519
rect 34360 2505 34363 2519
rect 34305 2495 34363 2505
rect 34305 2439 34306 2495
rect 34362 2439 34363 2495
rect 34305 2429 34363 2439
rect 34305 2415 34308 2429
rect 34360 2415 34363 2429
rect 34305 2359 34306 2415
rect 34362 2359 34363 2415
rect 34305 2335 34308 2359
rect 34360 2335 34363 2359
rect 34305 2279 34306 2335
rect 34362 2279 34363 2335
rect 34305 2255 34308 2279
rect 34360 2255 34363 2279
rect 34305 2199 34306 2255
rect 34362 2199 34363 2255
rect 34305 2185 34308 2199
rect 34360 2185 34363 2199
rect 34305 2175 34363 2185
rect 34305 2119 34306 2175
rect 34362 2119 34363 2175
rect 34305 2109 34363 2119
rect 34305 2095 34308 2109
rect 34360 2095 34363 2109
rect 34305 2039 34306 2095
rect 34362 2039 34363 2095
rect 34305 2015 34308 2039
rect 34360 2015 34363 2039
rect 34305 1959 34306 2015
rect 34362 1959 34363 2015
rect 34305 1935 34308 1959
rect 34360 1935 34363 1959
rect 34305 1879 34306 1935
rect 34362 1879 34363 1935
rect 34305 1865 34308 1879
rect 34360 1865 34363 1879
rect 34305 1855 34363 1865
rect 34305 1799 34306 1855
rect 34362 1799 34363 1855
rect 34305 1789 34363 1799
rect 34305 1775 34308 1789
rect 34360 1775 34363 1789
rect 34305 1719 34306 1775
rect 34362 1719 34363 1775
rect 34305 1695 34308 1719
rect 34360 1695 34363 1719
rect 34305 1639 34306 1695
rect 34362 1639 34363 1695
rect 34305 1615 34308 1639
rect 34360 1615 34363 1639
rect 34305 1559 34306 1615
rect 34362 1559 34363 1615
rect 34305 1545 34308 1559
rect 34360 1545 34363 1559
rect 34305 1535 34363 1545
rect 34305 1479 34306 1535
rect 34362 1479 34363 1535
rect 34305 1469 34363 1479
rect 34305 1455 34308 1469
rect 34360 1455 34363 1469
rect 34305 1399 34306 1455
rect 34362 1399 34363 1455
rect 34305 1375 34308 1399
rect 34360 1375 34363 1399
rect 34305 1319 34306 1375
rect 34362 1319 34363 1375
rect 34305 1295 34308 1319
rect 34360 1295 34363 1319
rect 34305 1239 34306 1295
rect 34362 1239 34363 1295
rect 34305 1225 34308 1239
rect 34360 1225 34363 1239
rect 34305 1215 34363 1225
rect 34305 1159 34306 1215
rect 34362 1159 34363 1215
rect 34305 1147 34363 1159
rect 34401 3133 34459 3147
rect 34401 3081 34404 3133
rect 34456 3081 34459 3133
rect 34401 3069 34459 3081
rect 34401 3017 34404 3069
rect 34456 3017 34459 3069
rect 34401 3005 34459 3017
rect 34401 2953 34404 3005
rect 34456 2953 34459 3005
rect 34401 2941 34459 2953
rect 34401 2889 34404 2941
rect 34456 2889 34459 2941
rect 34401 2877 34459 2889
rect 34401 2825 34404 2877
rect 34456 2825 34459 2877
rect 34401 2813 34459 2825
rect 34401 2761 34404 2813
rect 34456 2761 34459 2813
rect 34401 2749 34459 2761
rect 34401 2697 34404 2749
rect 34456 2697 34459 2749
rect 34401 2685 34459 2697
rect 34401 2633 34404 2685
rect 34456 2633 34459 2685
rect 34401 2621 34459 2633
rect 34401 2569 34404 2621
rect 34456 2569 34459 2621
rect 34401 2557 34459 2569
rect 34401 2505 34404 2557
rect 34456 2505 34459 2557
rect 34401 2493 34459 2505
rect 34401 2441 34404 2493
rect 34456 2441 34459 2493
rect 34401 2429 34459 2441
rect 34401 2377 34404 2429
rect 34456 2377 34459 2429
rect 34401 2365 34459 2377
rect 34401 2313 34404 2365
rect 34456 2313 34459 2365
rect 34401 2301 34459 2313
rect 34401 2249 34404 2301
rect 34456 2249 34459 2301
rect 34401 2237 34459 2249
rect 34401 2185 34404 2237
rect 34456 2185 34459 2237
rect 34401 2173 34459 2185
rect 34401 2121 34404 2173
rect 34456 2121 34459 2173
rect 34401 2109 34459 2121
rect 34401 2057 34404 2109
rect 34456 2057 34459 2109
rect 34401 2045 34459 2057
rect 34401 1993 34404 2045
rect 34456 1993 34459 2045
rect 34401 1981 34459 1993
rect 34401 1929 34404 1981
rect 34456 1929 34459 1981
rect 34401 1917 34459 1929
rect 34401 1865 34404 1917
rect 34456 1865 34459 1917
rect 34401 1853 34459 1865
rect 34401 1801 34404 1853
rect 34456 1801 34459 1853
rect 34401 1789 34459 1801
rect 34401 1737 34404 1789
rect 34456 1737 34459 1789
rect 34401 1725 34459 1737
rect 34401 1673 34404 1725
rect 34456 1673 34459 1725
rect 34401 1661 34459 1673
rect 34401 1609 34404 1661
rect 34456 1609 34459 1661
rect 34401 1597 34459 1609
rect 34401 1545 34404 1597
rect 34456 1545 34459 1597
rect 34401 1533 34459 1545
rect 34401 1481 34404 1533
rect 34456 1481 34459 1533
rect 34401 1469 34459 1481
rect 34401 1417 34404 1469
rect 34456 1417 34459 1469
rect 34401 1405 34459 1417
rect 34401 1353 34404 1405
rect 34456 1353 34459 1405
rect 34401 1341 34459 1353
rect 34401 1289 34404 1341
rect 34456 1289 34459 1341
rect 34401 1277 34459 1289
rect 34401 1225 34404 1277
rect 34456 1225 34459 1277
rect 34401 1213 34459 1225
rect 34401 1161 34404 1213
rect 34456 1161 34459 1213
rect 34401 830 34459 1161
rect 34497 3135 34555 3147
rect 34497 3079 34498 3135
rect 34554 3079 34555 3135
rect 34497 3069 34555 3079
rect 34497 3055 34500 3069
rect 34552 3055 34555 3069
rect 34497 2999 34498 3055
rect 34554 2999 34555 3055
rect 34497 2975 34500 2999
rect 34552 2975 34555 2999
rect 34497 2919 34498 2975
rect 34554 2919 34555 2975
rect 34497 2895 34500 2919
rect 34552 2895 34555 2919
rect 34497 2839 34498 2895
rect 34554 2839 34555 2895
rect 34497 2825 34500 2839
rect 34552 2825 34555 2839
rect 34497 2815 34555 2825
rect 34497 2759 34498 2815
rect 34554 2759 34555 2815
rect 34497 2749 34555 2759
rect 34497 2735 34500 2749
rect 34552 2735 34555 2749
rect 34497 2679 34498 2735
rect 34554 2679 34555 2735
rect 34497 2655 34500 2679
rect 34552 2655 34555 2679
rect 34497 2599 34498 2655
rect 34554 2599 34555 2655
rect 34497 2575 34500 2599
rect 34552 2575 34555 2599
rect 34497 2519 34498 2575
rect 34554 2519 34555 2575
rect 34497 2505 34500 2519
rect 34552 2505 34555 2519
rect 34497 2495 34555 2505
rect 34497 2439 34498 2495
rect 34554 2439 34555 2495
rect 34497 2429 34555 2439
rect 34497 2415 34500 2429
rect 34552 2415 34555 2429
rect 34497 2359 34498 2415
rect 34554 2359 34555 2415
rect 34497 2335 34500 2359
rect 34552 2335 34555 2359
rect 34497 2279 34498 2335
rect 34554 2279 34555 2335
rect 34497 2255 34500 2279
rect 34552 2255 34555 2279
rect 34497 2199 34498 2255
rect 34554 2199 34555 2255
rect 34497 2185 34500 2199
rect 34552 2185 34555 2199
rect 34497 2175 34555 2185
rect 34497 2119 34498 2175
rect 34554 2119 34555 2175
rect 34497 2109 34555 2119
rect 34497 2095 34500 2109
rect 34552 2095 34555 2109
rect 34497 2039 34498 2095
rect 34554 2039 34555 2095
rect 34497 2015 34500 2039
rect 34552 2015 34555 2039
rect 34497 1959 34498 2015
rect 34554 1959 34555 2015
rect 34497 1935 34500 1959
rect 34552 1935 34555 1959
rect 34497 1879 34498 1935
rect 34554 1879 34555 1935
rect 34497 1865 34500 1879
rect 34552 1865 34555 1879
rect 34497 1855 34555 1865
rect 34497 1799 34498 1855
rect 34554 1799 34555 1855
rect 34497 1789 34555 1799
rect 34497 1775 34500 1789
rect 34552 1775 34555 1789
rect 34497 1719 34498 1775
rect 34554 1719 34555 1775
rect 34497 1695 34500 1719
rect 34552 1695 34555 1719
rect 34497 1639 34498 1695
rect 34554 1639 34555 1695
rect 34497 1615 34500 1639
rect 34552 1615 34555 1639
rect 34497 1559 34498 1615
rect 34554 1559 34555 1615
rect 34497 1545 34500 1559
rect 34552 1545 34555 1559
rect 34497 1535 34555 1545
rect 34497 1479 34498 1535
rect 34554 1479 34555 1535
rect 34497 1469 34555 1479
rect 34497 1455 34500 1469
rect 34552 1455 34555 1469
rect 34497 1399 34498 1455
rect 34554 1399 34555 1455
rect 34497 1375 34500 1399
rect 34552 1375 34555 1399
rect 34497 1319 34498 1375
rect 34554 1319 34555 1375
rect 34497 1295 34500 1319
rect 34552 1295 34555 1319
rect 34497 1239 34498 1295
rect 34554 1239 34555 1295
rect 34497 1225 34500 1239
rect 34552 1225 34555 1239
rect 34497 1215 34555 1225
rect 34497 1159 34498 1215
rect 34554 1159 34555 1215
rect 34497 1147 34555 1159
rect 34593 3133 34651 3147
rect 34593 3081 34596 3133
rect 34648 3081 34651 3133
rect 34593 3069 34651 3081
rect 34593 3017 34596 3069
rect 34648 3017 34651 3069
rect 34593 3005 34651 3017
rect 34593 2953 34596 3005
rect 34648 2953 34651 3005
rect 34593 2941 34651 2953
rect 34593 2889 34596 2941
rect 34648 2889 34651 2941
rect 34593 2877 34651 2889
rect 34593 2825 34596 2877
rect 34648 2825 34651 2877
rect 34593 2813 34651 2825
rect 34593 2761 34596 2813
rect 34648 2761 34651 2813
rect 34593 2749 34651 2761
rect 34593 2697 34596 2749
rect 34648 2697 34651 2749
rect 34593 2685 34651 2697
rect 34593 2633 34596 2685
rect 34648 2633 34651 2685
rect 34593 2621 34651 2633
rect 34593 2569 34596 2621
rect 34648 2569 34651 2621
rect 34593 2557 34651 2569
rect 34593 2505 34596 2557
rect 34648 2505 34651 2557
rect 34593 2493 34651 2505
rect 34593 2441 34596 2493
rect 34648 2441 34651 2493
rect 34593 2429 34651 2441
rect 34593 2377 34596 2429
rect 34648 2377 34651 2429
rect 34593 2365 34651 2377
rect 34593 2313 34596 2365
rect 34648 2313 34651 2365
rect 34593 2301 34651 2313
rect 34593 2249 34596 2301
rect 34648 2249 34651 2301
rect 34593 2237 34651 2249
rect 34593 2185 34596 2237
rect 34648 2185 34651 2237
rect 34593 2173 34651 2185
rect 34593 2121 34596 2173
rect 34648 2121 34651 2173
rect 34593 2109 34651 2121
rect 34593 2057 34596 2109
rect 34648 2057 34651 2109
rect 34593 2045 34651 2057
rect 34593 1993 34596 2045
rect 34648 1993 34651 2045
rect 34593 1981 34651 1993
rect 34593 1929 34596 1981
rect 34648 1929 34651 1981
rect 34593 1917 34651 1929
rect 34593 1865 34596 1917
rect 34648 1865 34651 1917
rect 34593 1853 34651 1865
rect 34593 1801 34596 1853
rect 34648 1801 34651 1853
rect 34593 1789 34651 1801
rect 34593 1737 34596 1789
rect 34648 1737 34651 1789
rect 34593 1725 34651 1737
rect 34593 1673 34596 1725
rect 34648 1673 34651 1725
rect 34593 1661 34651 1673
rect 34593 1609 34596 1661
rect 34648 1609 34651 1661
rect 34593 1597 34651 1609
rect 34593 1545 34596 1597
rect 34648 1545 34651 1597
rect 34593 1533 34651 1545
rect 34593 1481 34596 1533
rect 34648 1481 34651 1533
rect 34593 1469 34651 1481
rect 34593 1417 34596 1469
rect 34648 1417 34651 1469
rect 34593 1405 34651 1417
rect 34593 1353 34596 1405
rect 34648 1353 34651 1405
rect 34593 1341 34651 1353
rect 34593 1289 34596 1341
rect 34648 1289 34651 1341
rect 34593 1277 34651 1289
rect 34593 1225 34596 1277
rect 34648 1225 34651 1277
rect 34593 1213 34651 1225
rect 34593 1161 34596 1213
rect 34648 1161 34651 1213
rect 34593 830 34651 1161
rect 34689 3135 34747 3147
rect 34689 3079 34690 3135
rect 34746 3079 34747 3135
rect 34689 3069 34747 3079
rect 34689 3055 34692 3069
rect 34744 3055 34747 3069
rect 34689 2999 34690 3055
rect 34746 2999 34747 3055
rect 34689 2975 34692 2999
rect 34744 2975 34747 2999
rect 34689 2919 34690 2975
rect 34746 2919 34747 2975
rect 34689 2895 34692 2919
rect 34744 2895 34747 2919
rect 34689 2839 34690 2895
rect 34746 2839 34747 2895
rect 34689 2825 34692 2839
rect 34744 2825 34747 2839
rect 34689 2815 34747 2825
rect 34689 2759 34690 2815
rect 34746 2759 34747 2815
rect 34689 2749 34747 2759
rect 34689 2735 34692 2749
rect 34744 2735 34747 2749
rect 34689 2679 34690 2735
rect 34746 2679 34747 2735
rect 34689 2655 34692 2679
rect 34744 2655 34747 2679
rect 34689 2599 34690 2655
rect 34746 2599 34747 2655
rect 34689 2575 34692 2599
rect 34744 2575 34747 2599
rect 34689 2519 34690 2575
rect 34746 2519 34747 2575
rect 34689 2505 34692 2519
rect 34744 2505 34747 2519
rect 34689 2495 34747 2505
rect 34689 2439 34690 2495
rect 34746 2439 34747 2495
rect 34689 2429 34747 2439
rect 34689 2415 34692 2429
rect 34744 2415 34747 2429
rect 34689 2359 34690 2415
rect 34746 2359 34747 2415
rect 34689 2335 34692 2359
rect 34744 2335 34747 2359
rect 34689 2279 34690 2335
rect 34746 2279 34747 2335
rect 34689 2255 34692 2279
rect 34744 2255 34747 2279
rect 34689 2199 34690 2255
rect 34746 2199 34747 2255
rect 34689 2185 34692 2199
rect 34744 2185 34747 2199
rect 34689 2175 34747 2185
rect 34689 2119 34690 2175
rect 34746 2119 34747 2175
rect 34689 2109 34747 2119
rect 34689 2095 34692 2109
rect 34744 2095 34747 2109
rect 34689 2039 34690 2095
rect 34746 2039 34747 2095
rect 34689 2015 34692 2039
rect 34744 2015 34747 2039
rect 34689 1959 34690 2015
rect 34746 1959 34747 2015
rect 34689 1935 34692 1959
rect 34744 1935 34747 1959
rect 34689 1879 34690 1935
rect 34746 1879 34747 1935
rect 34689 1865 34692 1879
rect 34744 1865 34747 1879
rect 34689 1855 34747 1865
rect 34689 1799 34690 1855
rect 34746 1799 34747 1855
rect 34689 1789 34747 1799
rect 34689 1775 34692 1789
rect 34744 1775 34747 1789
rect 34689 1719 34690 1775
rect 34746 1719 34747 1775
rect 34689 1695 34692 1719
rect 34744 1695 34747 1719
rect 34689 1639 34690 1695
rect 34746 1639 34747 1695
rect 34689 1615 34692 1639
rect 34744 1615 34747 1639
rect 34689 1559 34690 1615
rect 34746 1559 34747 1615
rect 34689 1545 34692 1559
rect 34744 1545 34747 1559
rect 34689 1535 34747 1545
rect 34689 1479 34690 1535
rect 34746 1479 34747 1535
rect 34689 1469 34747 1479
rect 34689 1455 34692 1469
rect 34744 1455 34747 1469
rect 34689 1399 34690 1455
rect 34746 1399 34747 1455
rect 34689 1375 34692 1399
rect 34744 1375 34747 1399
rect 34689 1319 34690 1375
rect 34746 1319 34747 1375
rect 34689 1295 34692 1319
rect 34744 1295 34747 1319
rect 34689 1239 34690 1295
rect 34746 1239 34747 1295
rect 34689 1225 34692 1239
rect 34744 1225 34747 1239
rect 34689 1215 34747 1225
rect 34689 1159 34690 1215
rect 34746 1159 34747 1215
rect 34689 1147 34747 1159
rect 34785 3133 34843 3147
rect 34785 3081 34788 3133
rect 34840 3081 34843 3133
rect 34785 3069 34843 3081
rect 34785 3017 34788 3069
rect 34840 3017 34843 3069
rect 34785 3005 34843 3017
rect 34785 2953 34788 3005
rect 34840 2953 34843 3005
rect 34785 2941 34843 2953
rect 34785 2889 34788 2941
rect 34840 2889 34843 2941
rect 34785 2877 34843 2889
rect 34785 2825 34788 2877
rect 34840 2825 34843 2877
rect 34785 2813 34843 2825
rect 34785 2761 34788 2813
rect 34840 2761 34843 2813
rect 34785 2749 34843 2761
rect 34785 2697 34788 2749
rect 34840 2697 34843 2749
rect 34785 2685 34843 2697
rect 34785 2633 34788 2685
rect 34840 2633 34843 2685
rect 34785 2621 34843 2633
rect 34785 2569 34788 2621
rect 34840 2569 34843 2621
rect 34785 2557 34843 2569
rect 34785 2505 34788 2557
rect 34840 2505 34843 2557
rect 34785 2493 34843 2505
rect 34785 2441 34788 2493
rect 34840 2441 34843 2493
rect 34785 2429 34843 2441
rect 34785 2377 34788 2429
rect 34840 2377 34843 2429
rect 34785 2365 34843 2377
rect 34785 2313 34788 2365
rect 34840 2313 34843 2365
rect 34785 2301 34843 2313
rect 34785 2249 34788 2301
rect 34840 2249 34843 2301
rect 34785 2237 34843 2249
rect 34785 2185 34788 2237
rect 34840 2185 34843 2237
rect 34785 2173 34843 2185
rect 34785 2121 34788 2173
rect 34840 2121 34843 2173
rect 34785 2109 34843 2121
rect 34785 2057 34788 2109
rect 34840 2057 34843 2109
rect 34785 2045 34843 2057
rect 34785 1993 34788 2045
rect 34840 1993 34843 2045
rect 34785 1981 34843 1993
rect 34785 1929 34788 1981
rect 34840 1929 34843 1981
rect 34785 1917 34843 1929
rect 34785 1865 34788 1917
rect 34840 1865 34843 1917
rect 34785 1853 34843 1865
rect 34785 1801 34788 1853
rect 34840 1801 34843 1853
rect 34785 1789 34843 1801
rect 34785 1737 34788 1789
rect 34840 1737 34843 1789
rect 34785 1725 34843 1737
rect 34785 1673 34788 1725
rect 34840 1673 34843 1725
rect 34785 1661 34843 1673
rect 34785 1609 34788 1661
rect 34840 1609 34843 1661
rect 34785 1597 34843 1609
rect 34785 1545 34788 1597
rect 34840 1545 34843 1597
rect 34785 1533 34843 1545
rect 34785 1481 34788 1533
rect 34840 1481 34843 1533
rect 34785 1469 34843 1481
rect 34785 1417 34788 1469
rect 34840 1417 34843 1469
rect 34785 1405 34843 1417
rect 34785 1353 34788 1405
rect 34840 1353 34843 1405
rect 34785 1341 34843 1353
rect 34785 1289 34788 1341
rect 34840 1289 34843 1341
rect 34785 1277 34843 1289
rect 34785 1225 34788 1277
rect 34840 1225 34843 1277
rect 34785 1213 34843 1225
rect 34785 1161 34788 1213
rect 34840 1161 34843 1213
rect 34785 830 34843 1161
rect 34881 3135 34939 3147
rect 34881 3079 34882 3135
rect 34938 3079 34939 3135
rect 34881 3069 34939 3079
rect 34881 3055 34884 3069
rect 34936 3055 34939 3069
rect 34881 2999 34882 3055
rect 34938 2999 34939 3055
rect 34881 2975 34884 2999
rect 34936 2975 34939 2999
rect 34881 2919 34882 2975
rect 34938 2919 34939 2975
rect 34881 2895 34884 2919
rect 34936 2895 34939 2919
rect 34881 2839 34882 2895
rect 34938 2839 34939 2895
rect 34881 2825 34884 2839
rect 34936 2825 34939 2839
rect 34881 2815 34939 2825
rect 34881 2759 34882 2815
rect 34938 2759 34939 2815
rect 34881 2749 34939 2759
rect 34881 2735 34884 2749
rect 34936 2735 34939 2749
rect 34881 2679 34882 2735
rect 34938 2679 34939 2735
rect 34881 2655 34884 2679
rect 34936 2655 34939 2679
rect 34881 2599 34882 2655
rect 34938 2599 34939 2655
rect 34881 2575 34884 2599
rect 34936 2575 34939 2599
rect 34881 2519 34882 2575
rect 34938 2519 34939 2575
rect 34881 2505 34884 2519
rect 34936 2505 34939 2519
rect 34881 2495 34939 2505
rect 34881 2439 34882 2495
rect 34938 2439 34939 2495
rect 34881 2429 34939 2439
rect 34881 2415 34884 2429
rect 34936 2415 34939 2429
rect 34881 2359 34882 2415
rect 34938 2359 34939 2415
rect 34881 2335 34884 2359
rect 34936 2335 34939 2359
rect 34881 2279 34882 2335
rect 34938 2279 34939 2335
rect 34881 2255 34884 2279
rect 34936 2255 34939 2279
rect 34881 2199 34882 2255
rect 34938 2199 34939 2255
rect 34881 2185 34884 2199
rect 34936 2185 34939 2199
rect 34881 2175 34939 2185
rect 34881 2119 34882 2175
rect 34938 2119 34939 2175
rect 34881 2109 34939 2119
rect 34881 2095 34884 2109
rect 34936 2095 34939 2109
rect 34881 2039 34882 2095
rect 34938 2039 34939 2095
rect 34881 2015 34884 2039
rect 34936 2015 34939 2039
rect 34881 1959 34882 2015
rect 34938 1959 34939 2015
rect 34881 1935 34884 1959
rect 34936 1935 34939 1959
rect 34881 1879 34882 1935
rect 34938 1879 34939 1935
rect 34881 1865 34884 1879
rect 34936 1865 34939 1879
rect 34881 1855 34939 1865
rect 34881 1799 34882 1855
rect 34938 1799 34939 1855
rect 34881 1789 34939 1799
rect 34881 1775 34884 1789
rect 34936 1775 34939 1789
rect 34881 1719 34882 1775
rect 34938 1719 34939 1775
rect 34881 1695 34884 1719
rect 34936 1695 34939 1719
rect 34881 1639 34882 1695
rect 34938 1639 34939 1695
rect 34881 1615 34884 1639
rect 34936 1615 34939 1639
rect 34881 1559 34882 1615
rect 34938 1559 34939 1615
rect 34881 1545 34884 1559
rect 34936 1545 34939 1559
rect 34881 1535 34939 1545
rect 34881 1479 34882 1535
rect 34938 1479 34939 1535
rect 34881 1469 34939 1479
rect 34881 1455 34884 1469
rect 34936 1455 34939 1469
rect 34881 1399 34882 1455
rect 34938 1399 34939 1455
rect 34881 1375 34884 1399
rect 34936 1375 34939 1399
rect 34881 1319 34882 1375
rect 34938 1319 34939 1375
rect 34881 1295 34884 1319
rect 34936 1295 34939 1319
rect 34881 1239 34882 1295
rect 34938 1239 34939 1295
rect 34881 1225 34884 1239
rect 34936 1225 34939 1239
rect 34881 1215 34939 1225
rect 34881 1159 34882 1215
rect 34938 1159 34939 1215
rect 34881 1147 34939 1159
rect 34977 3133 35035 3147
rect 34977 3081 34980 3133
rect 35032 3081 35035 3133
rect 34977 3069 35035 3081
rect 34977 3017 34980 3069
rect 35032 3017 35035 3069
rect 34977 3005 35035 3017
rect 34977 2953 34980 3005
rect 35032 2953 35035 3005
rect 34977 2941 35035 2953
rect 34977 2889 34980 2941
rect 35032 2889 35035 2941
rect 34977 2877 35035 2889
rect 34977 2825 34980 2877
rect 35032 2825 35035 2877
rect 34977 2813 35035 2825
rect 34977 2761 34980 2813
rect 35032 2761 35035 2813
rect 34977 2749 35035 2761
rect 34977 2697 34980 2749
rect 35032 2697 35035 2749
rect 34977 2685 35035 2697
rect 34977 2633 34980 2685
rect 35032 2633 35035 2685
rect 34977 2621 35035 2633
rect 34977 2569 34980 2621
rect 35032 2569 35035 2621
rect 34977 2557 35035 2569
rect 34977 2505 34980 2557
rect 35032 2505 35035 2557
rect 34977 2493 35035 2505
rect 34977 2441 34980 2493
rect 35032 2441 35035 2493
rect 34977 2429 35035 2441
rect 34977 2377 34980 2429
rect 35032 2377 35035 2429
rect 34977 2365 35035 2377
rect 34977 2313 34980 2365
rect 35032 2313 35035 2365
rect 34977 2301 35035 2313
rect 34977 2249 34980 2301
rect 35032 2249 35035 2301
rect 34977 2237 35035 2249
rect 34977 2185 34980 2237
rect 35032 2185 35035 2237
rect 34977 2173 35035 2185
rect 34977 2121 34980 2173
rect 35032 2121 35035 2173
rect 34977 2109 35035 2121
rect 34977 2057 34980 2109
rect 35032 2057 35035 2109
rect 34977 2045 35035 2057
rect 34977 1993 34980 2045
rect 35032 1993 35035 2045
rect 34977 1981 35035 1993
rect 34977 1929 34980 1981
rect 35032 1929 35035 1981
rect 34977 1917 35035 1929
rect 34977 1865 34980 1917
rect 35032 1865 35035 1917
rect 34977 1853 35035 1865
rect 34977 1801 34980 1853
rect 35032 1801 35035 1853
rect 34977 1789 35035 1801
rect 34977 1737 34980 1789
rect 35032 1737 35035 1789
rect 34977 1725 35035 1737
rect 34977 1673 34980 1725
rect 35032 1673 35035 1725
rect 34977 1661 35035 1673
rect 34977 1609 34980 1661
rect 35032 1609 35035 1661
rect 34977 1597 35035 1609
rect 34977 1545 34980 1597
rect 35032 1545 35035 1597
rect 34977 1533 35035 1545
rect 34977 1481 34980 1533
rect 35032 1481 35035 1533
rect 34977 1469 35035 1481
rect 34977 1417 34980 1469
rect 35032 1417 35035 1469
rect 34977 1405 35035 1417
rect 34977 1353 34980 1405
rect 35032 1353 35035 1405
rect 34977 1341 35035 1353
rect 34977 1289 34980 1341
rect 35032 1289 35035 1341
rect 34977 1277 35035 1289
rect 34977 1225 34980 1277
rect 35032 1225 35035 1277
rect 34977 1213 35035 1225
rect 34977 1161 34980 1213
rect 35032 1161 35035 1213
rect 34977 830 35035 1161
rect 35073 3135 35131 3147
rect 35073 3079 35074 3135
rect 35130 3079 35131 3135
rect 35073 3069 35131 3079
rect 35073 3055 35076 3069
rect 35128 3055 35131 3069
rect 35073 2999 35074 3055
rect 35130 2999 35131 3055
rect 35073 2975 35076 2999
rect 35128 2975 35131 2999
rect 35073 2919 35074 2975
rect 35130 2919 35131 2975
rect 35073 2895 35076 2919
rect 35128 2895 35131 2919
rect 35073 2839 35074 2895
rect 35130 2839 35131 2895
rect 35073 2825 35076 2839
rect 35128 2825 35131 2839
rect 35073 2815 35131 2825
rect 35073 2759 35074 2815
rect 35130 2759 35131 2815
rect 35073 2749 35131 2759
rect 35073 2735 35076 2749
rect 35128 2735 35131 2749
rect 35073 2679 35074 2735
rect 35130 2679 35131 2735
rect 35073 2655 35076 2679
rect 35128 2655 35131 2679
rect 35073 2599 35074 2655
rect 35130 2599 35131 2655
rect 35073 2575 35076 2599
rect 35128 2575 35131 2599
rect 35073 2519 35074 2575
rect 35130 2519 35131 2575
rect 35073 2505 35076 2519
rect 35128 2505 35131 2519
rect 35073 2495 35131 2505
rect 35073 2439 35074 2495
rect 35130 2439 35131 2495
rect 35073 2429 35131 2439
rect 35073 2415 35076 2429
rect 35128 2415 35131 2429
rect 35073 2359 35074 2415
rect 35130 2359 35131 2415
rect 35073 2335 35076 2359
rect 35128 2335 35131 2359
rect 35073 2279 35074 2335
rect 35130 2279 35131 2335
rect 35073 2255 35076 2279
rect 35128 2255 35131 2279
rect 35073 2199 35074 2255
rect 35130 2199 35131 2255
rect 35073 2185 35076 2199
rect 35128 2185 35131 2199
rect 35073 2175 35131 2185
rect 35073 2119 35074 2175
rect 35130 2119 35131 2175
rect 35073 2109 35131 2119
rect 35073 2095 35076 2109
rect 35128 2095 35131 2109
rect 35073 2039 35074 2095
rect 35130 2039 35131 2095
rect 35073 2015 35076 2039
rect 35128 2015 35131 2039
rect 35073 1959 35074 2015
rect 35130 1959 35131 2015
rect 35073 1935 35076 1959
rect 35128 1935 35131 1959
rect 35073 1879 35074 1935
rect 35130 1879 35131 1935
rect 35073 1865 35076 1879
rect 35128 1865 35131 1879
rect 35073 1855 35131 1865
rect 35073 1799 35074 1855
rect 35130 1799 35131 1855
rect 35073 1789 35131 1799
rect 35073 1775 35076 1789
rect 35128 1775 35131 1789
rect 35073 1719 35074 1775
rect 35130 1719 35131 1775
rect 35073 1695 35076 1719
rect 35128 1695 35131 1719
rect 35073 1639 35074 1695
rect 35130 1639 35131 1695
rect 35073 1615 35076 1639
rect 35128 1615 35131 1639
rect 35073 1559 35074 1615
rect 35130 1559 35131 1615
rect 35073 1545 35076 1559
rect 35128 1545 35131 1559
rect 35073 1535 35131 1545
rect 35073 1479 35074 1535
rect 35130 1479 35131 1535
rect 35073 1469 35131 1479
rect 35073 1455 35076 1469
rect 35128 1455 35131 1469
rect 35073 1399 35074 1455
rect 35130 1399 35131 1455
rect 35073 1375 35076 1399
rect 35128 1375 35131 1399
rect 35073 1319 35074 1375
rect 35130 1319 35131 1375
rect 35073 1295 35076 1319
rect 35128 1295 35131 1319
rect 35073 1239 35074 1295
rect 35130 1239 35131 1295
rect 35073 1225 35076 1239
rect 35128 1225 35131 1239
rect 35073 1215 35131 1225
rect 35073 1159 35074 1215
rect 35130 1159 35131 1215
rect 35073 1147 35131 1159
rect 35169 3133 35227 3147
rect 35169 3081 35172 3133
rect 35224 3081 35227 3133
rect 35169 3069 35227 3081
rect 35169 3017 35172 3069
rect 35224 3017 35227 3069
rect 35169 3005 35227 3017
rect 35169 2953 35172 3005
rect 35224 2953 35227 3005
rect 35169 2941 35227 2953
rect 35169 2889 35172 2941
rect 35224 2889 35227 2941
rect 35169 2877 35227 2889
rect 35169 2825 35172 2877
rect 35224 2825 35227 2877
rect 35169 2813 35227 2825
rect 35169 2761 35172 2813
rect 35224 2761 35227 2813
rect 35169 2749 35227 2761
rect 35169 2697 35172 2749
rect 35224 2697 35227 2749
rect 35169 2685 35227 2697
rect 35169 2633 35172 2685
rect 35224 2633 35227 2685
rect 35169 2621 35227 2633
rect 35169 2569 35172 2621
rect 35224 2569 35227 2621
rect 35169 2557 35227 2569
rect 35169 2505 35172 2557
rect 35224 2505 35227 2557
rect 35169 2493 35227 2505
rect 35169 2441 35172 2493
rect 35224 2441 35227 2493
rect 35169 2429 35227 2441
rect 35169 2377 35172 2429
rect 35224 2377 35227 2429
rect 35169 2365 35227 2377
rect 35169 2313 35172 2365
rect 35224 2313 35227 2365
rect 35169 2301 35227 2313
rect 35169 2249 35172 2301
rect 35224 2249 35227 2301
rect 35169 2237 35227 2249
rect 35169 2185 35172 2237
rect 35224 2185 35227 2237
rect 35169 2173 35227 2185
rect 35169 2121 35172 2173
rect 35224 2121 35227 2173
rect 35169 2109 35227 2121
rect 35169 2057 35172 2109
rect 35224 2057 35227 2109
rect 35169 2045 35227 2057
rect 35169 1993 35172 2045
rect 35224 1993 35227 2045
rect 35169 1981 35227 1993
rect 35169 1929 35172 1981
rect 35224 1929 35227 1981
rect 35169 1917 35227 1929
rect 35169 1865 35172 1917
rect 35224 1865 35227 1917
rect 35169 1853 35227 1865
rect 35169 1801 35172 1853
rect 35224 1801 35227 1853
rect 35169 1789 35227 1801
rect 35169 1737 35172 1789
rect 35224 1737 35227 1789
rect 35169 1725 35227 1737
rect 35169 1673 35172 1725
rect 35224 1673 35227 1725
rect 35169 1661 35227 1673
rect 35169 1609 35172 1661
rect 35224 1609 35227 1661
rect 35169 1597 35227 1609
rect 35169 1545 35172 1597
rect 35224 1545 35227 1597
rect 35169 1533 35227 1545
rect 35169 1481 35172 1533
rect 35224 1481 35227 1533
rect 35169 1469 35227 1481
rect 35169 1417 35172 1469
rect 35224 1417 35227 1469
rect 35169 1405 35227 1417
rect 35169 1353 35172 1405
rect 35224 1353 35227 1405
rect 35169 1341 35227 1353
rect 35169 1289 35172 1341
rect 35224 1289 35227 1341
rect 35169 1277 35227 1289
rect 35169 1225 35172 1277
rect 35224 1225 35227 1277
rect 35169 1213 35227 1225
rect 35169 1161 35172 1213
rect 35224 1161 35227 1213
rect 35169 830 35227 1161
rect 35265 3135 35323 3147
rect 35265 3079 35266 3135
rect 35322 3079 35323 3135
rect 35265 3069 35323 3079
rect 35265 3055 35268 3069
rect 35320 3055 35323 3069
rect 35265 2999 35266 3055
rect 35322 2999 35323 3055
rect 35265 2975 35268 2999
rect 35320 2975 35323 2999
rect 35265 2919 35266 2975
rect 35322 2919 35323 2975
rect 35265 2895 35268 2919
rect 35320 2895 35323 2919
rect 35265 2839 35266 2895
rect 35322 2839 35323 2895
rect 35265 2825 35268 2839
rect 35320 2825 35323 2839
rect 35265 2815 35323 2825
rect 35265 2759 35266 2815
rect 35322 2759 35323 2815
rect 35265 2749 35323 2759
rect 35265 2735 35268 2749
rect 35320 2735 35323 2749
rect 35265 2679 35266 2735
rect 35322 2679 35323 2735
rect 35265 2655 35268 2679
rect 35320 2655 35323 2679
rect 35265 2599 35266 2655
rect 35322 2599 35323 2655
rect 35265 2575 35268 2599
rect 35320 2575 35323 2599
rect 35265 2519 35266 2575
rect 35322 2519 35323 2575
rect 35265 2505 35268 2519
rect 35320 2505 35323 2519
rect 35265 2495 35323 2505
rect 35265 2439 35266 2495
rect 35322 2439 35323 2495
rect 35265 2429 35323 2439
rect 35265 2415 35268 2429
rect 35320 2415 35323 2429
rect 35265 2359 35266 2415
rect 35322 2359 35323 2415
rect 35265 2335 35268 2359
rect 35320 2335 35323 2359
rect 35265 2279 35266 2335
rect 35322 2279 35323 2335
rect 35265 2255 35268 2279
rect 35320 2255 35323 2279
rect 35265 2199 35266 2255
rect 35322 2199 35323 2255
rect 35265 2185 35268 2199
rect 35320 2185 35323 2199
rect 35265 2175 35323 2185
rect 35265 2119 35266 2175
rect 35322 2119 35323 2175
rect 35265 2109 35323 2119
rect 35265 2095 35268 2109
rect 35320 2095 35323 2109
rect 35265 2039 35266 2095
rect 35322 2039 35323 2095
rect 35265 2015 35268 2039
rect 35320 2015 35323 2039
rect 35265 1959 35266 2015
rect 35322 1959 35323 2015
rect 35265 1935 35268 1959
rect 35320 1935 35323 1959
rect 35265 1879 35266 1935
rect 35322 1879 35323 1935
rect 35265 1865 35268 1879
rect 35320 1865 35323 1879
rect 35265 1855 35323 1865
rect 35265 1799 35266 1855
rect 35322 1799 35323 1855
rect 35265 1789 35323 1799
rect 35265 1775 35268 1789
rect 35320 1775 35323 1789
rect 35265 1719 35266 1775
rect 35322 1719 35323 1775
rect 35265 1695 35268 1719
rect 35320 1695 35323 1719
rect 35265 1639 35266 1695
rect 35322 1639 35323 1695
rect 35265 1615 35268 1639
rect 35320 1615 35323 1639
rect 35265 1559 35266 1615
rect 35322 1559 35323 1615
rect 35265 1545 35268 1559
rect 35320 1545 35323 1559
rect 35265 1535 35323 1545
rect 35265 1479 35266 1535
rect 35322 1479 35323 1535
rect 35265 1469 35323 1479
rect 35265 1455 35268 1469
rect 35320 1455 35323 1469
rect 35265 1399 35266 1455
rect 35322 1399 35323 1455
rect 35265 1375 35268 1399
rect 35320 1375 35323 1399
rect 35265 1319 35266 1375
rect 35322 1319 35323 1375
rect 35265 1295 35268 1319
rect 35320 1295 35323 1319
rect 35265 1239 35266 1295
rect 35322 1239 35323 1295
rect 35265 1225 35268 1239
rect 35320 1225 35323 1239
rect 35265 1215 35323 1225
rect 35265 1159 35266 1215
rect 35322 1159 35323 1215
rect 35265 1147 35323 1159
rect 35361 3133 35419 3147
rect 35361 3081 35364 3133
rect 35416 3081 35419 3133
rect 35361 3069 35419 3081
rect 35361 3017 35364 3069
rect 35416 3017 35419 3069
rect 35361 3005 35419 3017
rect 35361 2953 35364 3005
rect 35416 2953 35419 3005
rect 35361 2941 35419 2953
rect 35361 2889 35364 2941
rect 35416 2889 35419 2941
rect 35361 2877 35419 2889
rect 35361 2825 35364 2877
rect 35416 2825 35419 2877
rect 35361 2813 35419 2825
rect 35361 2761 35364 2813
rect 35416 2761 35419 2813
rect 35361 2749 35419 2761
rect 35361 2697 35364 2749
rect 35416 2697 35419 2749
rect 35361 2685 35419 2697
rect 35361 2633 35364 2685
rect 35416 2633 35419 2685
rect 35361 2621 35419 2633
rect 35361 2569 35364 2621
rect 35416 2569 35419 2621
rect 35361 2557 35419 2569
rect 35361 2505 35364 2557
rect 35416 2505 35419 2557
rect 35361 2493 35419 2505
rect 35361 2441 35364 2493
rect 35416 2441 35419 2493
rect 35361 2429 35419 2441
rect 35361 2377 35364 2429
rect 35416 2377 35419 2429
rect 35361 2365 35419 2377
rect 35361 2313 35364 2365
rect 35416 2313 35419 2365
rect 35361 2301 35419 2313
rect 35361 2249 35364 2301
rect 35416 2249 35419 2301
rect 35361 2237 35419 2249
rect 35361 2185 35364 2237
rect 35416 2185 35419 2237
rect 35361 2173 35419 2185
rect 35361 2121 35364 2173
rect 35416 2121 35419 2173
rect 35361 2109 35419 2121
rect 35361 2057 35364 2109
rect 35416 2057 35419 2109
rect 35361 2045 35419 2057
rect 35361 1993 35364 2045
rect 35416 1993 35419 2045
rect 35361 1981 35419 1993
rect 35361 1929 35364 1981
rect 35416 1929 35419 1981
rect 35361 1917 35419 1929
rect 35361 1865 35364 1917
rect 35416 1865 35419 1917
rect 35361 1853 35419 1865
rect 35361 1801 35364 1853
rect 35416 1801 35419 1853
rect 35361 1789 35419 1801
rect 35361 1737 35364 1789
rect 35416 1737 35419 1789
rect 35361 1725 35419 1737
rect 35361 1673 35364 1725
rect 35416 1673 35419 1725
rect 35361 1661 35419 1673
rect 35361 1609 35364 1661
rect 35416 1609 35419 1661
rect 35361 1597 35419 1609
rect 35361 1545 35364 1597
rect 35416 1545 35419 1597
rect 35361 1533 35419 1545
rect 35361 1481 35364 1533
rect 35416 1481 35419 1533
rect 35361 1469 35419 1481
rect 35361 1417 35364 1469
rect 35416 1417 35419 1469
rect 35361 1405 35419 1417
rect 35361 1353 35364 1405
rect 35416 1353 35419 1405
rect 35361 1341 35419 1353
rect 35361 1289 35364 1341
rect 35416 1289 35419 1341
rect 35361 1277 35419 1289
rect 35361 1225 35364 1277
rect 35416 1225 35419 1277
rect 35361 1213 35419 1225
rect 35361 1161 35364 1213
rect 35416 1161 35419 1213
rect 35361 830 35419 1161
rect 35457 3135 35515 3147
rect 35457 3079 35458 3135
rect 35514 3079 35515 3135
rect 35457 3069 35515 3079
rect 35457 3055 35460 3069
rect 35512 3055 35515 3069
rect 35457 2999 35458 3055
rect 35514 2999 35515 3055
rect 35457 2975 35460 2999
rect 35512 2975 35515 2999
rect 35457 2919 35458 2975
rect 35514 2919 35515 2975
rect 35457 2895 35460 2919
rect 35512 2895 35515 2919
rect 35457 2839 35458 2895
rect 35514 2839 35515 2895
rect 35457 2825 35460 2839
rect 35512 2825 35515 2839
rect 35457 2815 35515 2825
rect 35457 2759 35458 2815
rect 35514 2759 35515 2815
rect 35457 2749 35515 2759
rect 35457 2735 35460 2749
rect 35512 2735 35515 2749
rect 35457 2679 35458 2735
rect 35514 2679 35515 2735
rect 35457 2655 35460 2679
rect 35512 2655 35515 2679
rect 35457 2599 35458 2655
rect 35514 2599 35515 2655
rect 35457 2575 35460 2599
rect 35512 2575 35515 2599
rect 35457 2519 35458 2575
rect 35514 2519 35515 2575
rect 35457 2505 35460 2519
rect 35512 2505 35515 2519
rect 35457 2495 35515 2505
rect 35457 2439 35458 2495
rect 35514 2439 35515 2495
rect 35457 2429 35515 2439
rect 35457 2415 35460 2429
rect 35512 2415 35515 2429
rect 35457 2359 35458 2415
rect 35514 2359 35515 2415
rect 35457 2335 35460 2359
rect 35512 2335 35515 2359
rect 35457 2279 35458 2335
rect 35514 2279 35515 2335
rect 35457 2255 35460 2279
rect 35512 2255 35515 2279
rect 35457 2199 35458 2255
rect 35514 2199 35515 2255
rect 35457 2185 35460 2199
rect 35512 2185 35515 2199
rect 35457 2175 35515 2185
rect 35457 2119 35458 2175
rect 35514 2119 35515 2175
rect 35457 2109 35515 2119
rect 35457 2095 35460 2109
rect 35512 2095 35515 2109
rect 35457 2039 35458 2095
rect 35514 2039 35515 2095
rect 35457 2015 35460 2039
rect 35512 2015 35515 2039
rect 35457 1959 35458 2015
rect 35514 1959 35515 2015
rect 35457 1935 35460 1959
rect 35512 1935 35515 1959
rect 35457 1879 35458 1935
rect 35514 1879 35515 1935
rect 35457 1865 35460 1879
rect 35512 1865 35515 1879
rect 35457 1855 35515 1865
rect 35457 1799 35458 1855
rect 35514 1799 35515 1855
rect 35457 1789 35515 1799
rect 35457 1775 35460 1789
rect 35512 1775 35515 1789
rect 35457 1719 35458 1775
rect 35514 1719 35515 1775
rect 35457 1695 35460 1719
rect 35512 1695 35515 1719
rect 35457 1639 35458 1695
rect 35514 1639 35515 1695
rect 35457 1615 35460 1639
rect 35512 1615 35515 1639
rect 35457 1559 35458 1615
rect 35514 1559 35515 1615
rect 35457 1545 35460 1559
rect 35512 1545 35515 1559
rect 35457 1535 35515 1545
rect 35457 1479 35458 1535
rect 35514 1479 35515 1535
rect 35457 1469 35515 1479
rect 35457 1455 35460 1469
rect 35512 1455 35515 1469
rect 35457 1399 35458 1455
rect 35514 1399 35515 1455
rect 35457 1375 35460 1399
rect 35512 1375 35515 1399
rect 35457 1319 35458 1375
rect 35514 1319 35515 1375
rect 35457 1295 35460 1319
rect 35512 1295 35515 1319
rect 35457 1239 35458 1295
rect 35514 1239 35515 1295
rect 35457 1225 35460 1239
rect 35512 1225 35515 1239
rect 35457 1215 35515 1225
rect 35457 1159 35458 1215
rect 35514 1159 35515 1215
rect 35457 1147 35515 1159
rect 35553 3133 35611 3147
rect 35553 3081 35556 3133
rect 35608 3081 35611 3133
rect 35553 3069 35611 3081
rect 35553 3017 35556 3069
rect 35608 3017 35611 3069
rect 35553 3005 35611 3017
rect 35553 2953 35556 3005
rect 35608 2953 35611 3005
rect 35553 2941 35611 2953
rect 35553 2889 35556 2941
rect 35608 2889 35611 2941
rect 35553 2877 35611 2889
rect 35553 2825 35556 2877
rect 35608 2825 35611 2877
rect 35553 2813 35611 2825
rect 35553 2761 35556 2813
rect 35608 2761 35611 2813
rect 35553 2749 35611 2761
rect 35553 2697 35556 2749
rect 35608 2697 35611 2749
rect 35553 2685 35611 2697
rect 35553 2633 35556 2685
rect 35608 2633 35611 2685
rect 35553 2621 35611 2633
rect 35553 2569 35556 2621
rect 35608 2569 35611 2621
rect 35553 2557 35611 2569
rect 35553 2505 35556 2557
rect 35608 2505 35611 2557
rect 35553 2493 35611 2505
rect 35553 2441 35556 2493
rect 35608 2441 35611 2493
rect 35553 2429 35611 2441
rect 35553 2377 35556 2429
rect 35608 2377 35611 2429
rect 35553 2365 35611 2377
rect 35553 2313 35556 2365
rect 35608 2313 35611 2365
rect 35553 2301 35611 2313
rect 35553 2249 35556 2301
rect 35608 2249 35611 2301
rect 35553 2237 35611 2249
rect 35553 2185 35556 2237
rect 35608 2185 35611 2237
rect 35553 2173 35611 2185
rect 35553 2121 35556 2173
rect 35608 2121 35611 2173
rect 35553 2109 35611 2121
rect 35553 2057 35556 2109
rect 35608 2057 35611 2109
rect 35553 2045 35611 2057
rect 35553 1993 35556 2045
rect 35608 1993 35611 2045
rect 35553 1981 35611 1993
rect 35553 1929 35556 1981
rect 35608 1929 35611 1981
rect 35553 1917 35611 1929
rect 35553 1865 35556 1917
rect 35608 1865 35611 1917
rect 35553 1853 35611 1865
rect 35553 1801 35556 1853
rect 35608 1801 35611 1853
rect 35553 1789 35611 1801
rect 35553 1737 35556 1789
rect 35608 1737 35611 1789
rect 35553 1725 35611 1737
rect 35553 1673 35556 1725
rect 35608 1673 35611 1725
rect 35553 1661 35611 1673
rect 35553 1609 35556 1661
rect 35608 1609 35611 1661
rect 35553 1597 35611 1609
rect 35553 1545 35556 1597
rect 35608 1545 35611 1597
rect 35553 1533 35611 1545
rect 35553 1481 35556 1533
rect 35608 1481 35611 1533
rect 35553 1469 35611 1481
rect 35553 1417 35556 1469
rect 35608 1417 35611 1469
rect 35553 1405 35611 1417
rect 35553 1353 35556 1405
rect 35608 1353 35611 1405
rect 35553 1341 35611 1353
rect 35553 1289 35556 1341
rect 35608 1289 35611 1341
rect 35553 1277 35611 1289
rect 35553 1225 35556 1277
rect 35608 1225 35611 1277
rect 35553 1213 35611 1225
rect 35553 1161 35556 1213
rect 35608 1161 35611 1213
rect 35553 830 35611 1161
rect 35649 3135 35707 3147
rect 35649 3079 35650 3135
rect 35706 3079 35707 3135
rect 35649 3069 35707 3079
rect 35649 3055 35652 3069
rect 35704 3055 35707 3069
rect 35649 2999 35650 3055
rect 35706 2999 35707 3055
rect 35649 2975 35652 2999
rect 35704 2975 35707 2999
rect 35649 2919 35650 2975
rect 35706 2919 35707 2975
rect 35649 2895 35652 2919
rect 35704 2895 35707 2919
rect 35649 2839 35650 2895
rect 35706 2839 35707 2895
rect 35649 2825 35652 2839
rect 35704 2825 35707 2839
rect 35649 2815 35707 2825
rect 35649 2759 35650 2815
rect 35706 2759 35707 2815
rect 35649 2749 35707 2759
rect 35649 2735 35652 2749
rect 35704 2735 35707 2749
rect 35649 2679 35650 2735
rect 35706 2679 35707 2735
rect 35649 2655 35652 2679
rect 35704 2655 35707 2679
rect 35649 2599 35650 2655
rect 35706 2599 35707 2655
rect 35649 2575 35652 2599
rect 35704 2575 35707 2599
rect 35649 2519 35650 2575
rect 35706 2519 35707 2575
rect 35649 2505 35652 2519
rect 35704 2505 35707 2519
rect 35649 2495 35707 2505
rect 35649 2439 35650 2495
rect 35706 2439 35707 2495
rect 35649 2429 35707 2439
rect 35649 2415 35652 2429
rect 35704 2415 35707 2429
rect 35649 2359 35650 2415
rect 35706 2359 35707 2415
rect 35649 2335 35652 2359
rect 35704 2335 35707 2359
rect 35649 2279 35650 2335
rect 35706 2279 35707 2335
rect 35649 2255 35652 2279
rect 35704 2255 35707 2279
rect 35649 2199 35650 2255
rect 35706 2199 35707 2255
rect 35649 2185 35652 2199
rect 35704 2185 35707 2199
rect 35649 2175 35707 2185
rect 35649 2119 35650 2175
rect 35706 2119 35707 2175
rect 35649 2109 35707 2119
rect 35649 2095 35652 2109
rect 35704 2095 35707 2109
rect 35649 2039 35650 2095
rect 35706 2039 35707 2095
rect 35649 2015 35652 2039
rect 35704 2015 35707 2039
rect 35649 1959 35650 2015
rect 35706 1959 35707 2015
rect 35649 1935 35652 1959
rect 35704 1935 35707 1959
rect 35649 1879 35650 1935
rect 35706 1879 35707 1935
rect 35649 1865 35652 1879
rect 35704 1865 35707 1879
rect 35649 1855 35707 1865
rect 35649 1799 35650 1855
rect 35706 1799 35707 1855
rect 35649 1789 35707 1799
rect 35649 1775 35652 1789
rect 35704 1775 35707 1789
rect 35649 1719 35650 1775
rect 35706 1719 35707 1775
rect 35649 1695 35652 1719
rect 35704 1695 35707 1719
rect 35649 1639 35650 1695
rect 35706 1639 35707 1695
rect 35649 1615 35652 1639
rect 35704 1615 35707 1639
rect 35649 1559 35650 1615
rect 35706 1559 35707 1615
rect 35649 1545 35652 1559
rect 35704 1545 35707 1559
rect 35649 1535 35707 1545
rect 35649 1479 35650 1535
rect 35706 1479 35707 1535
rect 35649 1469 35707 1479
rect 35649 1455 35652 1469
rect 35704 1455 35707 1469
rect 35649 1399 35650 1455
rect 35706 1399 35707 1455
rect 35649 1375 35652 1399
rect 35704 1375 35707 1399
rect 35649 1319 35650 1375
rect 35706 1319 35707 1375
rect 35649 1295 35652 1319
rect 35704 1295 35707 1319
rect 35649 1239 35650 1295
rect 35706 1239 35707 1295
rect 35649 1225 35652 1239
rect 35704 1225 35707 1239
rect 35649 1215 35707 1225
rect 35649 1159 35650 1215
rect 35706 1159 35707 1215
rect 35649 1147 35707 1159
rect 35745 3133 35803 3147
rect 35745 3081 35748 3133
rect 35800 3081 35803 3133
rect 35745 3069 35803 3081
rect 35745 3017 35748 3069
rect 35800 3017 35803 3069
rect 35745 3005 35803 3017
rect 35745 2953 35748 3005
rect 35800 2953 35803 3005
rect 35745 2941 35803 2953
rect 35745 2889 35748 2941
rect 35800 2889 35803 2941
rect 35745 2877 35803 2889
rect 35745 2825 35748 2877
rect 35800 2825 35803 2877
rect 35745 2813 35803 2825
rect 35745 2761 35748 2813
rect 35800 2761 35803 2813
rect 35745 2749 35803 2761
rect 35745 2697 35748 2749
rect 35800 2697 35803 2749
rect 35745 2685 35803 2697
rect 35745 2633 35748 2685
rect 35800 2633 35803 2685
rect 35745 2621 35803 2633
rect 35745 2569 35748 2621
rect 35800 2569 35803 2621
rect 35745 2557 35803 2569
rect 35745 2505 35748 2557
rect 35800 2505 35803 2557
rect 35745 2493 35803 2505
rect 35745 2441 35748 2493
rect 35800 2441 35803 2493
rect 35745 2429 35803 2441
rect 35745 2377 35748 2429
rect 35800 2377 35803 2429
rect 35745 2365 35803 2377
rect 35745 2313 35748 2365
rect 35800 2313 35803 2365
rect 35745 2301 35803 2313
rect 35745 2249 35748 2301
rect 35800 2249 35803 2301
rect 35745 2237 35803 2249
rect 35745 2185 35748 2237
rect 35800 2185 35803 2237
rect 35745 2173 35803 2185
rect 35745 2121 35748 2173
rect 35800 2121 35803 2173
rect 35745 2109 35803 2121
rect 35745 2057 35748 2109
rect 35800 2057 35803 2109
rect 35745 2045 35803 2057
rect 35745 1993 35748 2045
rect 35800 1993 35803 2045
rect 35745 1981 35803 1993
rect 35745 1929 35748 1981
rect 35800 1929 35803 1981
rect 35745 1917 35803 1929
rect 35745 1865 35748 1917
rect 35800 1865 35803 1917
rect 35745 1853 35803 1865
rect 35745 1801 35748 1853
rect 35800 1801 35803 1853
rect 35745 1789 35803 1801
rect 35745 1737 35748 1789
rect 35800 1737 35803 1789
rect 35745 1725 35803 1737
rect 35745 1673 35748 1725
rect 35800 1673 35803 1725
rect 35745 1661 35803 1673
rect 35745 1609 35748 1661
rect 35800 1609 35803 1661
rect 35745 1597 35803 1609
rect 35745 1545 35748 1597
rect 35800 1545 35803 1597
rect 35745 1533 35803 1545
rect 35745 1481 35748 1533
rect 35800 1481 35803 1533
rect 35745 1469 35803 1481
rect 35745 1417 35748 1469
rect 35800 1417 35803 1469
rect 35745 1405 35803 1417
rect 35745 1353 35748 1405
rect 35800 1353 35803 1405
rect 35745 1341 35803 1353
rect 35745 1289 35748 1341
rect 35800 1289 35803 1341
rect 35745 1277 35803 1289
rect 35745 1225 35748 1277
rect 35800 1225 35803 1277
rect 35745 1213 35803 1225
rect 35745 1161 35748 1213
rect 35800 1161 35803 1213
rect 35745 830 35803 1161
rect 35841 3135 35899 3147
rect 35841 3079 35842 3135
rect 35898 3079 35899 3135
rect 35841 3069 35899 3079
rect 35841 3055 35844 3069
rect 35896 3055 35899 3069
rect 35841 2999 35842 3055
rect 35898 2999 35899 3055
rect 35841 2975 35844 2999
rect 35896 2975 35899 2999
rect 35841 2919 35842 2975
rect 35898 2919 35899 2975
rect 35841 2895 35844 2919
rect 35896 2895 35899 2919
rect 35841 2839 35842 2895
rect 35898 2839 35899 2895
rect 35841 2825 35844 2839
rect 35896 2825 35899 2839
rect 35841 2815 35899 2825
rect 35841 2759 35842 2815
rect 35898 2759 35899 2815
rect 35841 2749 35899 2759
rect 35841 2735 35844 2749
rect 35896 2735 35899 2749
rect 35841 2679 35842 2735
rect 35898 2679 35899 2735
rect 35841 2655 35844 2679
rect 35896 2655 35899 2679
rect 35841 2599 35842 2655
rect 35898 2599 35899 2655
rect 35841 2575 35844 2599
rect 35896 2575 35899 2599
rect 35841 2519 35842 2575
rect 35898 2519 35899 2575
rect 35841 2505 35844 2519
rect 35896 2505 35899 2519
rect 35841 2495 35899 2505
rect 35841 2439 35842 2495
rect 35898 2439 35899 2495
rect 35841 2429 35899 2439
rect 35841 2415 35844 2429
rect 35896 2415 35899 2429
rect 35841 2359 35842 2415
rect 35898 2359 35899 2415
rect 35841 2335 35844 2359
rect 35896 2335 35899 2359
rect 35841 2279 35842 2335
rect 35898 2279 35899 2335
rect 35841 2255 35844 2279
rect 35896 2255 35899 2279
rect 35841 2199 35842 2255
rect 35898 2199 35899 2255
rect 35841 2185 35844 2199
rect 35896 2185 35899 2199
rect 35841 2175 35899 2185
rect 35841 2119 35842 2175
rect 35898 2119 35899 2175
rect 35841 2109 35899 2119
rect 35841 2095 35844 2109
rect 35896 2095 35899 2109
rect 35841 2039 35842 2095
rect 35898 2039 35899 2095
rect 35841 2015 35844 2039
rect 35896 2015 35899 2039
rect 35841 1959 35842 2015
rect 35898 1959 35899 2015
rect 35841 1935 35844 1959
rect 35896 1935 35899 1959
rect 35841 1879 35842 1935
rect 35898 1879 35899 1935
rect 35841 1865 35844 1879
rect 35896 1865 35899 1879
rect 35841 1855 35899 1865
rect 35841 1799 35842 1855
rect 35898 1799 35899 1855
rect 35841 1789 35899 1799
rect 35841 1775 35844 1789
rect 35896 1775 35899 1789
rect 35841 1719 35842 1775
rect 35898 1719 35899 1775
rect 35841 1695 35844 1719
rect 35896 1695 35899 1719
rect 35841 1639 35842 1695
rect 35898 1639 35899 1695
rect 35841 1615 35844 1639
rect 35896 1615 35899 1639
rect 35841 1559 35842 1615
rect 35898 1559 35899 1615
rect 35841 1545 35844 1559
rect 35896 1545 35899 1559
rect 35841 1535 35899 1545
rect 35841 1479 35842 1535
rect 35898 1479 35899 1535
rect 35841 1469 35899 1479
rect 35841 1455 35844 1469
rect 35896 1455 35899 1469
rect 35841 1399 35842 1455
rect 35898 1399 35899 1455
rect 35841 1375 35844 1399
rect 35896 1375 35899 1399
rect 35841 1319 35842 1375
rect 35898 1319 35899 1375
rect 35841 1295 35844 1319
rect 35896 1295 35899 1319
rect 35841 1239 35842 1295
rect 35898 1239 35899 1295
rect 35841 1225 35844 1239
rect 35896 1225 35899 1239
rect 35841 1215 35899 1225
rect 35841 1159 35842 1215
rect 35898 1159 35899 1215
rect 35841 1147 35899 1159
rect 35937 3133 35995 3147
rect 35937 3081 35940 3133
rect 35992 3081 35995 3133
rect 35937 3069 35995 3081
rect 35937 3017 35940 3069
rect 35992 3017 35995 3069
rect 35937 3005 35995 3017
rect 35937 2953 35940 3005
rect 35992 2953 35995 3005
rect 35937 2941 35995 2953
rect 35937 2889 35940 2941
rect 35992 2889 35995 2941
rect 35937 2877 35995 2889
rect 35937 2825 35940 2877
rect 35992 2825 35995 2877
rect 35937 2813 35995 2825
rect 35937 2761 35940 2813
rect 35992 2761 35995 2813
rect 35937 2749 35995 2761
rect 35937 2697 35940 2749
rect 35992 2697 35995 2749
rect 35937 2685 35995 2697
rect 35937 2633 35940 2685
rect 35992 2633 35995 2685
rect 35937 2621 35995 2633
rect 35937 2569 35940 2621
rect 35992 2569 35995 2621
rect 35937 2557 35995 2569
rect 35937 2505 35940 2557
rect 35992 2505 35995 2557
rect 35937 2493 35995 2505
rect 35937 2441 35940 2493
rect 35992 2441 35995 2493
rect 35937 2429 35995 2441
rect 35937 2377 35940 2429
rect 35992 2377 35995 2429
rect 35937 2365 35995 2377
rect 35937 2313 35940 2365
rect 35992 2313 35995 2365
rect 35937 2301 35995 2313
rect 35937 2249 35940 2301
rect 35992 2249 35995 2301
rect 35937 2237 35995 2249
rect 35937 2185 35940 2237
rect 35992 2185 35995 2237
rect 35937 2173 35995 2185
rect 35937 2121 35940 2173
rect 35992 2121 35995 2173
rect 35937 2109 35995 2121
rect 35937 2057 35940 2109
rect 35992 2057 35995 2109
rect 35937 2045 35995 2057
rect 35937 1993 35940 2045
rect 35992 1993 35995 2045
rect 35937 1981 35995 1993
rect 35937 1929 35940 1981
rect 35992 1929 35995 1981
rect 35937 1917 35995 1929
rect 35937 1865 35940 1917
rect 35992 1865 35995 1917
rect 35937 1853 35995 1865
rect 35937 1801 35940 1853
rect 35992 1801 35995 1853
rect 35937 1789 35995 1801
rect 35937 1737 35940 1789
rect 35992 1737 35995 1789
rect 35937 1725 35995 1737
rect 35937 1673 35940 1725
rect 35992 1673 35995 1725
rect 35937 1661 35995 1673
rect 35937 1609 35940 1661
rect 35992 1609 35995 1661
rect 35937 1597 35995 1609
rect 35937 1545 35940 1597
rect 35992 1545 35995 1597
rect 35937 1533 35995 1545
rect 35937 1481 35940 1533
rect 35992 1481 35995 1533
rect 35937 1469 35995 1481
rect 35937 1417 35940 1469
rect 35992 1417 35995 1469
rect 35937 1405 35995 1417
rect 35937 1353 35940 1405
rect 35992 1353 35995 1405
rect 35937 1341 35995 1353
rect 35937 1289 35940 1341
rect 35992 1289 35995 1341
rect 35937 1277 35995 1289
rect 35937 1225 35940 1277
rect 35992 1225 35995 1277
rect 35937 1213 35995 1225
rect 35937 1161 35940 1213
rect 35992 1161 35995 1213
rect 35937 830 35995 1161
rect 36033 3135 36091 3147
rect 36033 3079 36034 3135
rect 36090 3079 36091 3135
rect 36033 3069 36091 3079
rect 36033 3055 36036 3069
rect 36088 3055 36091 3069
rect 36033 2999 36034 3055
rect 36090 2999 36091 3055
rect 36033 2975 36036 2999
rect 36088 2975 36091 2999
rect 36033 2919 36034 2975
rect 36090 2919 36091 2975
rect 36033 2895 36036 2919
rect 36088 2895 36091 2919
rect 36033 2839 36034 2895
rect 36090 2839 36091 2895
rect 36033 2825 36036 2839
rect 36088 2825 36091 2839
rect 36033 2815 36091 2825
rect 36033 2759 36034 2815
rect 36090 2759 36091 2815
rect 36033 2749 36091 2759
rect 36033 2735 36036 2749
rect 36088 2735 36091 2749
rect 36033 2679 36034 2735
rect 36090 2679 36091 2735
rect 36033 2655 36036 2679
rect 36088 2655 36091 2679
rect 36033 2599 36034 2655
rect 36090 2599 36091 2655
rect 36033 2575 36036 2599
rect 36088 2575 36091 2599
rect 36033 2519 36034 2575
rect 36090 2519 36091 2575
rect 36033 2505 36036 2519
rect 36088 2505 36091 2519
rect 36033 2495 36091 2505
rect 36033 2439 36034 2495
rect 36090 2439 36091 2495
rect 36033 2429 36091 2439
rect 36033 2415 36036 2429
rect 36088 2415 36091 2429
rect 36033 2359 36034 2415
rect 36090 2359 36091 2415
rect 36033 2335 36036 2359
rect 36088 2335 36091 2359
rect 36033 2279 36034 2335
rect 36090 2279 36091 2335
rect 36033 2255 36036 2279
rect 36088 2255 36091 2279
rect 36033 2199 36034 2255
rect 36090 2199 36091 2255
rect 36033 2185 36036 2199
rect 36088 2185 36091 2199
rect 36033 2175 36091 2185
rect 36033 2119 36034 2175
rect 36090 2119 36091 2175
rect 36033 2109 36091 2119
rect 36033 2095 36036 2109
rect 36088 2095 36091 2109
rect 36033 2039 36034 2095
rect 36090 2039 36091 2095
rect 36033 2015 36036 2039
rect 36088 2015 36091 2039
rect 36033 1959 36034 2015
rect 36090 1959 36091 2015
rect 36033 1935 36036 1959
rect 36088 1935 36091 1959
rect 36033 1879 36034 1935
rect 36090 1879 36091 1935
rect 36033 1865 36036 1879
rect 36088 1865 36091 1879
rect 36033 1855 36091 1865
rect 36033 1799 36034 1855
rect 36090 1799 36091 1855
rect 36033 1789 36091 1799
rect 36033 1775 36036 1789
rect 36088 1775 36091 1789
rect 36033 1719 36034 1775
rect 36090 1719 36091 1775
rect 36033 1695 36036 1719
rect 36088 1695 36091 1719
rect 36033 1639 36034 1695
rect 36090 1639 36091 1695
rect 36033 1615 36036 1639
rect 36088 1615 36091 1639
rect 36033 1559 36034 1615
rect 36090 1559 36091 1615
rect 36033 1545 36036 1559
rect 36088 1545 36091 1559
rect 36033 1535 36091 1545
rect 36033 1479 36034 1535
rect 36090 1479 36091 1535
rect 36033 1469 36091 1479
rect 36033 1455 36036 1469
rect 36088 1455 36091 1469
rect 36033 1399 36034 1455
rect 36090 1399 36091 1455
rect 36033 1375 36036 1399
rect 36088 1375 36091 1399
rect 36033 1319 36034 1375
rect 36090 1319 36091 1375
rect 36033 1295 36036 1319
rect 36088 1295 36091 1319
rect 36033 1239 36034 1295
rect 36090 1239 36091 1295
rect 36033 1225 36036 1239
rect 36088 1225 36091 1239
rect 36033 1215 36091 1225
rect 36033 1159 36034 1215
rect 36090 1159 36091 1215
rect 36033 1147 36091 1159
rect 36129 3133 36187 3147
rect 36129 3081 36132 3133
rect 36184 3081 36187 3133
rect 36129 3069 36187 3081
rect 36129 3017 36132 3069
rect 36184 3017 36187 3069
rect 36129 3005 36187 3017
rect 36129 2953 36132 3005
rect 36184 2953 36187 3005
rect 36129 2941 36187 2953
rect 36129 2889 36132 2941
rect 36184 2889 36187 2941
rect 36129 2877 36187 2889
rect 36129 2825 36132 2877
rect 36184 2825 36187 2877
rect 36129 2813 36187 2825
rect 36129 2761 36132 2813
rect 36184 2761 36187 2813
rect 36129 2749 36187 2761
rect 36129 2697 36132 2749
rect 36184 2697 36187 2749
rect 36129 2685 36187 2697
rect 36129 2633 36132 2685
rect 36184 2633 36187 2685
rect 36129 2621 36187 2633
rect 36129 2569 36132 2621
rect 36184 2569 36187 2621
rect 36129 2557 36187 2569
rect 36129 2505 36132 2557
rect 36184 2505 36187 2557
rect 36129 2493 36187 2505
rect 36129 2441 36132 2493
rect 36184 2441 36187 2493
rect 36129 2429 36187 2441
rect 36129 2377 36132 2429
rect 36184 2377 36187 2429
rect 36129 2365 36187 2377
rect 36129 2313 36132 2365
rect 36184 2313 36187 2365
rect 36129 2301 36187 2313
rect 36129 2249 36132 2301
rect 36184 2249 36187 2301
rect 36129 2237 36187 2249
rect 36129 2185 36132 2237
rect 36184 2185 36187 2237
rect 36129 2173 36187 2185
rect 36129 2121 36132 2173
rect 36184 2121 36187 2173
rect 36129 2109 36187 2121
rect 36129 2057 36132 2109
rect 36184 2057 36187 2109
rect 36129 2045 36187 2057
rect 36129 1993 36132 2045
rect 36184 1993 36187 2045
rect 36129 1981 36187 1993
rect 36129 1929 36132 1981
rect 36184 1929 36187 1981
rect 36129 1917 36187 1929
rect 36129 1865 36132 1917
rect 36184 1865 36187 1917
rect 36129 1853 36187 1865
rect 36129 1801 36132 1853
rect 36184 1801 36187 1853
rect 36129 1789 36187 1801
rect 36129 1737 36132 1789
rect 36184 1737 36187 1789
rect 36129 1725 36187 1737
rect 36129 1673 36132 1725
rect 36184 1673 36187 1725
rect 36129 1661 36187 1673
rect 36129 1609 36132 1661
rect 36184 1609 36187 1661
rect 36129 1597 36187 1609
rect 36129 1545 36132 1597
rect 36184 1545 36187 1597
rect 36129 1533 36187 1545
rect 36129 1481 36132 1533
rect 36184 1481 36187 1533
rect 36129 1469 36187 1481
rect 36129 1417 36132 1469
rect 36184 1417 36187 1469
rect 36129 1405 36187 1417
rect 36129 1353 36132 1405
rect 36184 1353 36187 1405
rect 36129 1341 36187 1353
rect 36129 1289 36132 1341
rect 36184 1289 36187 1341
rect 36129 1277 36187 1289
rect 36129 1225 36132 1277
rect 36184 1225 36187 1277
rect 36129 1213 36187 1225
rect 36129 1161 36132 1213
rect 36184 1161 36187 1213
rect 36129 830 36187 1161
rect 36225 3135 36283 3147
rect 36225 3079 36226 3135
rect 36282 3079 36283 3135
rect 36225 3069 36283 3079
rect 36225 3055 36228 3069
rect 36280 3055 36283 3069
rect 36225 2999 36226 3055
rect 36282 2999 36283 3055
rect 36225 2975 36228 2999
rect 36280 2975 36283 2999
rect 36225 2919 36226 2975
rect 36282 2919 36283 2975
rect 36225 2895 36228 2919
rect 36280 2895 36283 2919
rect 36225 2839 36226 2895
rect 36282 2839 36283 2895
rect 36225 2825 36228 2839
rect 36280 2825 36283 2839
rect 36225 2815 36283 2825
rect 36225 2759 36226 2815
rect 36282 2759 36283 2815
rect 36225 2749 36283 2759
rect 36225 2735 36228 2749
rect 36280 2735 36283 2749
rect 36225 2679 36226 2735
rect 36282 2679 36283 2735
rect 36225 2655 36228 2679
rect 36280 2655 36283 2679
rect 36225 2599 36226 2655
rect 36282 2599 36283 2655
rect 36225 2575 36228 2599
rect 36280 2575 36283 2599
rect 36225 2519 36226 2575
rect 36282 2519 36283 2575
rect 36225 2505 36228 2519
rect 36280 2505 36283 2519
rect 36225 2495 36283 2505
rect 36225 2439 36226 2495
rect 36282 2439 36283 2495
rect 36225 2429 36283 2439
rect 36225 2415 36228 2429
rect 36280 2415 36283 2429
rect 36225 2359 36226 2415
rect 36282 2359 36283 2415
rect 36225 2335 36228 2359
rect 36280 2335 36283 2359
rect 36225 2279 36226 2335
rect 36282 2279 36283 2335
rect 36225 2255 36228 2279
rect 36280 2255 36283 2279
rect 36225 2199 36226 2255
rect 36282 2199 36283 2255
rect 36225 2185 36228 2199
rect 36280 2185 36283 2199
rect 36225 2175 36283 2185
rect 36225 2119 36226 2175
rect 36282 2119 36283 2175
rect 36225 2109 36283 2119
rect 36225 2095 36228 2109
rect 36280 2095 36283 2109
rect 36225 2039 36226 2095
rect 36282 2039 36283 2095
rect 36225 2015 36228 2039
rect 36280 2015 36283 2039
rect 36225 1959 36226 2015
rect 36282 1959 36283 2015
rect 36225 1935 36228 1959
rect 36280 1935 36283 1959
rect 36225 1879 36226 1935
rect 36282 1879 36283 1935
rect 36225 1865 36228 1879
rect 36280 1865 36283 1879
rect 36225 1855 36283 1865
rect 36225 1799 36226 1855
rect 36282 1799 36283 1855
rect 36225 1789 36283 1799
rect 36225 1775 36228 1789
rect 36280 1775 36283 1789
rect 36225 1719 36226 1775
rect 36282 1719 36283 1775
rect 36225 1695 36228 1719
rect 36280 1695 36283 1719
rect 36225 1639 36226 1695
rect 36282 1639 36283 1695
rect 36225 1615 36228 1639
rect 36280 1615 36283 1639
rect 36225 1559 36226 1615
rect 36282 1559 36283 1615
rect 36225 1545 36228 1559
rect 36280 1545 36283 1559
rect 36225 1535 36283 1545
rect 36225 1479 36226 1535
rect 36282 1479 36283 1535
rect 36225 1469 36283 1479
rect 36225 1455 36228 1469
rect 36280 1455 36283 1469
rect 36225 1399 36226 1455
rect 36282 1399 36283 1455
rect 36225 1375 36228 1399
rect 36280 1375 36283 1399
rect 36225 1319 36226 1375
rect 36282 1319 36283 1375
rect 36225 1295 36228 1319
rect 36280 1295 36283 1319
rect 36225 1239 36226 1295
rect 36282 1239 36283 1295
rect 36225 1225 36228 1239
rect 36280 1225 36283 1239
rect 36225 1215 36283 1225
rect 36225 1159 36226 1215
rect 36282 1159 36283 1215
rect 36225 1147 36283 1159
rect 36321 3133 36379 3147
rect 36321 3081 36324 3133
rect 36376 3081 36379 3133
rect 36321 3069 36379 3081
rect 36321 3017 36324 3069
rect 36376 3017 36379 3069
rect 36321 3005 36379 3017
rect 36321 2953 36324 3005
rect 36376 2953 36379 3005
rect 36321 2941 36379 2953
rect 36321 2889 36324 2941
rect 36376 2889 36379 2941
rect 36321 2877 36379 2889
rect 36321 2825 36324 2877
rect 36376 2825 36379 2877
rect 36321 2813 36379 2825
rect 36321 2761 36324 2813
rect 36376 2761 36379 2813
rect 36321 2749 36379 2761
rect 36321 2697 36324 2749
rect 36376 2697 36379 2749
rect 36321 2685 36379 2697
rect 36321 2633 36324 2685
rect 36376 2633 36379 2685
rect 36321 2621 36379 2633
rect 36321 2569 36324 2621
rect 36376 2569 36379 2621
rect 36321 2557 36379 2569
rect 36321 2505 36324 2557
rect 36376 2505 36379 2557
rect 36321 2493 36379 2505
rect 36321 2441 36324 2493
rect 36376 2441 36379 2493
rect 36321 2429 36379 2441
rect 36321 2377 36324 2429
rect 36376 2377 36379 2429
rect 36321 2365 36379 2377
rect 36321 2313 36324 2365
rect 36376 2313 36379 2365
rect 36321 2301 36379 2313
rect 36321 2249 36324 2301
rect 36376 2249 36379 2301
rect 36321 2237 36379 2249
rect 36321 2185 36324 2237
rect 36376 2185 36379 2237
rect 36321 2173 36379 2185
rect 36321 2121 36324 2173
rect 36376 2121 36379 2173
rect 36321 2109 36379 2121
rect 36321 2057 36324 2109
rect 36376 2057 36379 2109
rect 36321 2045 36379 2057
rect 36321 1993 36324 2045
rect 36376 1993 36379 2045
rect 36321 1981 36379 1993
rect 36321 1929 36324 1981
rect 36376 1929 36379 1981
rect 36321 1917 36379 1929
rect 36321 1865 36324 1917
rect 36376 1865 36379 1917
rect 36321 1853 36379 1865
rect 36321 1801 36324 1853
rect 36376 1801 36379 1853
rect 36321 1789 36379 1801
rect 36321 1737 36324 1789
rect 36376 1737 36379 1789
rect 36321 1725 36379 1737
rect 36321 1673 36324 1725
rect 36376 1673 36379 1725
rect 36321 1661 36379 1673
rect 36321 1609 36324 1661
rect 36376 1609 36379 1661
rect 36321 1597 36379 1609
rect 36321 1545 36324 1597
rect 36376 1545 36379 1597
rect 36321 1533 36379 1545
rect 36321 1481 36324 1533
rect 36376 1481 36379 1533
rect 36321 1469 36379 1481
rect 36321 1417 36324 1469
rect 36376 1417 36379 1469
rect 36321 1405 36379 1417
rect 36321 1353 36324 1405
rect 36376 1353 36379 1405
rect 36321 1341 36379 1353
rect 36321 1289 36324 1341
rect 36376 1289 36379 1341
rect 36321 1277 36379 1289
rect 36321 1225 36324 1277
rect 36376 1225 36379 1277
rect 36321 1213 36379 1225
rect 36321 1161 36324 1213
rect 36376 1161 36379 1213
rect 36321 830 36379 1161
rect 36417 3135 36475 3147
rect 36417 3079 36418 3135
rect 36474 3079 36475 3135
rect 36417 3069 36475 3079
rect 36417 3055 36420 3069
rect 36472 3055 36475 3069
rect 36417 2999 36418 3055
rect 36474 2999 36475 3055
rect 36417 2975 36420 2999
rect 36472 2975 36475 2999
rect 36417 2919 36418 2975
rect 36474 2919 36475 2975
rect 36417 2895 36420 2919
rect 36472 2895 36475 2919
rect 36417 2839 36418 2895
rect 36474 2839 36475 2895
rect 36417 2825 36420 2839
rect 36472 2825 36475 2839
rect 36417 2815 36475 2825
rect 36417 2759 36418 2815
rect 36474 2759 36475 2815
rect 36417 2749 36475 2759
rect 36417 2735 36420 2749
rect 36472 2735 36475 2749
rect 36417 2679 36418 2735
rect 36474 2679 36475 2735
rect 36417 2655 36420 2679
rect 36472 2655 36475 2679
rect 36417 2599 36418 2655
rect 36474 2599 36475 2655
rect 36417 2575 36420 2599
rect 36472 2575 36475 2599
rect 36417 2519 36418 2575
rect 36474 2519 36475 2575
rect 36417 2505 36420 2519
rect 36472 2505 36475 2519
rect 36417 2495 36475 2505
rect 36417 2439 36418 2495
rect 36474 2439 36475 2495
rect 36417 2429 36475 2439
rect 36417 2415 36420 2429
rect 36472 2415 36475 2429
rect 36417 2359 36418 2415
rect 36474 2359 36475 2415
rect 36417 2335 36420 2359
rect 36472 2335 36475 2359
rect 36417 2279 36418 2335
rect 36474 2279 36475 2335
rect 36417 2255 36420 2279
rect 36472 2255 36475 2279
rect 36417 2199 36418 2255
rect 36474 2199 36475 2255
rect 36417 2185 36420 2199
rect 36472 2185 36475 2199
rect 36417 2175 36475 2185
rect 36417 2119 36418 2175
rect 36474 2119 36475 2175
rect 36417 2109 36475 2119
rect 36417 2095 36420 2109
rect 36472 2095 36475 2109
rect 36417 2039 36418 2095
rect 36474 2039 36475 2095
rect 36417 2015 36420 2039
rect 36472 2015 36475 2039
rect 36417 1959 36418 2015
rect 36474 1959 36475 2015
rect 36417 1935 36420 1959
rect 36472 1935 36475 1959
rect 36417 1879 36418 1935
rect 36474 1879 36475 1935
rect 36417 1865 36420 1879
rect 36472 1865 36475 1879
rect 36417 1855 36475 1865
rect 36417 1799 36418 1855
rect 36474 1799 36475 1855
rect 36417 1789 36475 1799
rect 36417 1775 36420 1789
rect 36472 1775 36475 1789
rect 36417 1719 36418 1775
rect 36474 1719 36475 1775
rect 36417 1695 36420 1719
rect 36472 1695 36475 1719
rect 36417 1639 36418 1695
rect 36474 1639 36475 1695
rect 36417 1615 36420 1639
rect 36472 1615 36475 1639
rect 36417 1559 36418 1615
rect 36474 1559 36475 1615
rect 36417 1545 36420 1559
rect 36472 1545 36475 1559
rect 36417 1535 36475 1545
rect 36417 1479 36418 1535
rect 36474 1479 36475 1535
rect 36417 1469 36475 1479
rect 36417 1455 36420 1469
rect 36472 1455 36475 1469
rect 36417 1399 36418 1455
rect 36474 1399 36475 1455
rect 36417 1375 36420 1399
rect 36472 1375 36475 1399
rect 36417 1319 36418 1375
rect 36474 1319 36475 1375
rect 36417 1295 36420 1319
rect 36472 1295 36475 1319
rect 36417 1239 36418 1295
rect 36474 1239 36475 1295
rect 36417 1225 36420 1239
rect 36472 1225 36475 1239
rect 36417 1215 36475 1225
rect 36417 1159 36418 1215
rect 36474 1159 36475 1215
rect 36417 1147 36475 1159
rect 36513 3133 36571 3147
rect 36513 3081 36516 3133
rect 36568 3081 36571 3133
rect 36513 3069 36571 3081
rect 36513 3017 36516 3069
rect 36568 3017 36571 3069
rect 36513 3005 36571 3017
rect 36513 2953 36516 3005
rect 36568 2953 36571 3005
rect 36513 2941 36571 2953
rect 36513 2889 36516 2941
rect 36568 2889 36571 2941
rect 36513 2877 36571 2889
rect 36513 2825 36516 2877
rect 36568 2825 36571 2877
rect 36513 2813 36571 2825
rect 36513 2761 36516 2813
rect 36568 2761 36571 2813
rect 36513 2749 36571 2761
rect 36513 2697 36516 2749
rect 36568 2697 36571 2749
rect 36513 2685 36571 2697
rect 36513 2633 36516 2685
rect 36568 2633 36571 2685
rect 36513 2621 36571 2633
rect 36513 2569 36516 2621
rect 36568 2569 36571 2621
rect 36513 2557 36571 2569
rect 36513 2505 36516 2557
rect 36568 2505 36571 2557
rect 36513 2493 36571 2505
rect 36513 2441 36516 2493
rect 36568 2441 36571 2493
rect 36513 2429 36571 2441
rect 36513 2377 36516 2429
rect 36568 2377 36571 2429
rect 36513 2365 36571 2377
rect 36513 2313 36516 2365
rect 36568 2313 36571 2365
rect 36513 2301 36571 2313
rect 36513 2249 36516 2301
rect 36568 2249 36571 2301
rect 36513 2237 36571 2249
rect 36513 2185 36516 2237
rect 36568 2185 36571 2237
rect 36513 2173 36571 2185
rect 36513 2121 36516 2173
rect 36568 2121 36571 2173
rect 36513 2109 36571 2121
rect 36513 2057 36516 2109
rect 36568 2057 36571 2109
rect 36513 2045 36571 2057
rect 36513 1993 36516 2045
rect 36568 1993 36571 2045
rect 36513 1981 36571 1993
rect 36513 1929 36516 1981
rect 36568 1929 36571 1981
rect 36513 1917 36571 1929
rect 36513 1865 36516 1917
rect 36568 1865 36571 1917
rect 36513 1853 36571 1865
rect 36513 1801 36516 1853
rect 36568 1801 36571 1853
rect 36513 1789 36571 1801
rect 36513 1737 36516 1789
rect 36568 1737 36571 1789
rect 36513 1725 36571 1737
rect 36513 1673 36516 1725
rect 36568 1673 36571 1725
rect 36513 1661 36571 1673
rect 36513 1609 36516 1661
rect 36568 1609 36571 1661
rect 36513 1597 36571 1609
rect 36513 1545 36516 1597
rect 36568 1545 36571 1597
rect 36513 1533 36571 1545
rect 36513 1481 36516 1533
rect 36568 1481 36571 1533
rect 36513 1469 36571 1481
rect 36513 1417 36516 1469
rect 36568 1417 36571 1469
rect 36513 1405 36571 1417
rect 36513 1353 36516 1405
rect 36568 1353 36571 1405
rect 36513 1341 36571 1353
rect 36513 1289 36516 1341
rect 36568 1289 36571 1341
rect 36513 1277 36571 1289
rect 36513 1225 36516 1277
rect 36568 1225 36571 1277
rect 36513 1213 36571 1225
rect 36513 1161 36516 1213
rect 36568 1161 36571 1213
rect 36513 830 36571 1161
rect 36609 3135 36667 3147
rect 36609 3079 36610 3135
rect 36666 3079 36667 3135
rect 36609 3069 36667 3079
rect 36609 3055 36612 3069
rect 36664 3055 36667 3069
rect 36609 2999 36610 3055
rect 36666 2999 36667 3055
rect 36609 2975 36612 2999
rect 36664 2975 36667 2999
rect 36609 2919 36610 2975
rect 36666 2919 36667 2975
rect 36609 2895 36612 2919
rect 36664 2895 36667 2919
rect 36609 2839 36610 2895
rect 36666 2839 36667 2895
rect 36609 2825 36612 2839
rect 36664 2825 36667 2839
rect 36609 2815 36667 2825
rect 36609 2759 36610 2815
rect 36666 2759 36667 2815
rect 36609 2749 36667 2759
rect 36609 2735 36612 2749
rect 36664 2735 36667 2749
rect 36609 2679 36610 2735
rect 36666 2679 36667 2735
rect 36609 2655 36612 2679
rect 36664 2655 36667 2679
rect 36609 2599 36610 2655
rect 36666 2599 36667 2655
rect 36609 2575 36612 2599
rect 36664 2575 36667 2599
rect 36609 2519 36610 2575
rect 36666 2519 36667 2575
rect 36609 2505 36612 2519
rect 36664 2505 36667 2519
rect 36609 2495 36667 2505
rect 36609 2439 36610 2495
rect 36666 2439 36667 2495
rect 36609 2429 36667 2439
rect 36609 2415 36612 2429
rect 36664 2415 36667 2429
rect 36609 2359 36610 2415
rect 36666 2359 36667 2415
rect 36609 2335 36612 2359
rect 36664 2335 36667 2359
rect 36609 2279 36610 2335
rect 36666 2279 36667 2335
rect 36609 2255 36612 2279
rect 36664 2255 36667 2279
rect 36609 2199 36610 2255
rect 36666 2199 36667 2255
rect 36609 2185 36612 2199
rect 36664 2185 36667 2199
rect 36609 2175 36667 2185
rect 36609 2119 36610 2175
rect 36666 2119 36667 2175
rect 36609 2109 36667 2119
rect 36609 2095 36612 2109
rect 36664 2095 36667 2109
rect 36609 2039 36610 2095
rect 36666 2039 36667 2095
rect 36609 2015 36612 2039
rect 36664 2015 36667 2039
rect 36609 1959 36610 2015
rect 36666 1959 36667 2015
rect 36609 1935 36612 1959
rect 36664 1935 36667 1959
rect 36609 1879 36610 1935
rect 36666 1879 36667 1935
rect 36609 1865 36612 1879
rect 36664 1865 36667 1879
rect 36609 1855 36667 1865
rect 36609 1799 36610 1855
rect 36666 1799 36667 1855
rect 36609 1789 36667 1799
rect 36609 1775 36612 1789
rect 36664 1775 36667 1789
rect 36609 1719 36610 1775
rect 36666 1719 36667 1775
rect 36609 1695 36612 1719
rect 36664 1695 36667 1719
rect 36609 1639 36610 1695
rect 36666 1639 36667 1695
rect 36609 1615 36612 1639
rect 36664 1615 36667 1639
rect 36609 1559 36610 1615
rect 36666 1559 36667 1615
rect 36609 1545 36612 1559
rect 36664 1545 36667 1559
rect 36609 1535 36667 1545
rect 36609 1479 36610 1535
rect 36666 1479 36667 1535
rect 36609 1469 36667 1479
rect 36609 1455 36612 1469
rect 36664 1455 36667 1469
rect 36609 1399 36610 1455
rect 36666 1399 36667 1455
rect 36609 1375 36612 1399
rect 36664 1375 36667 1399
rect 36609 1319 36610 1375
rect 36666 1319 36667 1375
rect 36609 1295 36612 1319
rect 36664 1295 36667 1319
rect 36609 1239 36610 1295
rect 36666 1239 36667 1295
rect 36609 1225 36612 1239
rect 36664 1225 36667 1239
rect 36609 1215 36667 1225
rect 36609 1159 36610 1215
rect 36666 1159 36667 1215
rect 36609 1147 36667 1159
rect 36705 3133 36763 3147
rect 36705 3081 36708 3133
rect 36760 3081 36763 3133
rect 36705 3069 36763 3081
rect 36705 3017 36708 3069
rect 36760 3017 36763 3069
rect 36705 3005 36763 3017
rect 36705 2953 36708 3005
rect 36760 2953 36763 3005
rect 36705 2941 36763 2953
rect 36705 2889 36708 2941
rect 36760 2889 36763 2941
rect 36705 2877 36763 2889
rect 36705 2825 36708 2877
rect 36760 2825 36763 2877
rect 36705 2813 36763 2825
rect 36705 2761 36708 2813
rect 36760 2761 36763 2813
rect 36705 2749 36763 2761
rect 36705 2697 36708 2749
rect 36760 2697 36763 2749
rect 36705 2685 36763 2697
rect 36705 2633 36708 2685
rect 36760 2633 36763 2685
rect 36705 2621 36763 2633
rect 36705 2569 36708 2621
rect 36760 2569 36763 2621
rect 36705 2557 36763 2569
rect 36705 2505 36708 2557
rect 36760 2505 36763 2557
rect 36705 2493 36763 2505
rect 36705 2441 36708 2493
rect 36760 2441 36763 2493
rect 36705 2429 36763 2441
rect 36705 2377 36708 2429
rect 36760 2377 36763 2429
rect 36705 2365 36763 2377
rect 36705 2313 36708 2365
rect 36760 2313 36763 2365
rect 36705 2301 36763 2313
rect 36705 2249 36708 2301
rect 36760 2249 36763 2301
rect 36705 2237 36763 2249
rect 36705 2185 36708 2237
rect 36760 2185 36763 2237
rect 36705 2173 36763 2185
rect 36705 2121 36708 2173
rect 36760 2121 36763 2173
rect 36705 2109 36763 2121
rect 36705 2057 36708 2109
rect 36760 2057 36763 2109
rect 36705 2045 36763 2057
rect 36705 1993 36708 2045
rect 36760 1993 36763 2045
rect 36705 1981 36763 1993
rect 36705 1929 36708 1981
rect 36760 1929 36763 1981
rect 36705 1917 36763 1929
rect 36705 1865 36708 1917
rect 36760 1865 36763 1917
rect 36705 1853 36763 1865
rect 36705 1801 36708 1853
rect 36760 1801 36763 1853
rect 36705 1789 36763 1801
rect 36705 1737 36708 1789
rect 36760 1737 36763 1789
rect 36705 1725 36763 1737
rect 36705 1673 36708 1725
rect 36760 1673 36763 1725
rect 36705 1661 36763 1673
rect 36705 1609 36708 1661
rect 36760 1609 36763 1661
rect 36705 1597 36763 1609
rect 36705 1545 36708 1597
rect 36760 1545 36763 1597
rect 36705 1533 36763 1545
rect 36705 1481 36708 1533
rect 36760 1481 36763 1533
rect 36705 1469 36763 1481
rect 36705 1417 36708 1469
rect 36760 1417 36763 1469
rect 36705 1405 36763 1417
rect 36705 1353 36708 1405
rect 36760 1353 36763 1405
rect 36705 1341 36763 1353
rect 36705 1289 36708 1341
rect 36760 1289 36763 1341
rect 36705 1277 36763 1289
rect 36705 1225 36708 1277
rect 36760 1225 36763 1277
rect 36705 1213 36763 1225
rect 36705 1161 36708 1213
rect 36760 1161 36763 1213
rect 36705 830 36763 1161
rect 36801 3135 36859 3147
rect 36801 3079 36802 3135
rect 36858 3079 36859 3135
rect 36801 3069 36859 3079
rect 36801 3055 36804 3069
rect 36856 3055 36859 3069
rect 36801 2999 36802 3055
rect 36858 2999 36859 3055
rect 36801 2975 36804 2999
rect 36856 2975 36859 2999
rect 36801 2919 36802 2975
rect 36858 2919 36859 2975
rect 36801 2895 36804 2919
rect 36856 2895 36859 2919
rect 36801 2839 36802 2895
rect 36858 2839 36859 2895
rect 36801 2825 36804 2839
rect 36856 2825 36859 2839
rect 36801 2815 36859 2825
rect 36801 2759 36802 2815
rect 36858 2759 36859 2815
rect 36801 2749 36859 2759
rect 36801 2735 36804 2749
rect 36856 2735 36859 2749
rect 36801 2679 36802 2735
rect 36858 2679 36859 2735
rect 36801 2655 36804 2679
rect 36856 2655 36859 2679
rect 36801 2599 36802 2655
rect 36858 2599 36859 2655
rect 36801 2575 36804 2599
rect 36856 2575 36859 2599
rect 36801 2519 36802 2575
rect 36858 2519 36859 2575
rect 36801 2505 36804 2519
rect 36856 2505 36859 2519
rect 36801 2495 36859 2505
rect 36801 2439 36802 2495
rect 36858 2439 36859 2495
rect 36801 2429 36859 2439
rect 36801 2415 36804 2429
rect 36856 2415 36859 2429
rect 36801 2359 36802 2415
rect 36858 2359 36859 2415
rect 36801 2335 36804 2359
rect 36856 2335 36859 2359
rect 36801 2279 36802 2335
rect 36858 2279 36859 2335
rect 36801 2255 36804 2279
rect 36856 2255 36859 2279
rect 36801 2199 36802 2255
rect 36858 2199 36859 2255
rect 36801 2185 36804 2199
rect 36856 2185 36859 2199
rect 36801 2175 36859 2185
rect 36801 2119 36802 2175
rect 36858 2119 36859 2175
rect 36801 2109 36859 2119
rect 36801 2095 36804 2109
rect 36856 2095 36859 2109
rect 36801 2039 36802 2095
rect 36858 2039 36859 2095
rect 36801 2015 36804 2039
rect 36856 2015 36859 2039
rect 36801 1959 36802 2015
rect 36858 1959 36859 2015
rect 36801 1935 36804 1959
rect 36856 1935 36859 1959
rect 36801 1879 36802 1935
rect 36858 1879 36859 1935
rect 36801 1865 36804 1879
rect 36856 1865 36859 1879
rect 36801 1855 36859 1865
rect 36801 1799 36802 1855
rect 36858 1799 36859 1855
rect 36801 1789 36859 1799
rect 36801 1775 36804 1789
rect 36856 1775 36859 1789
rect 36801 1719 36802 1775
rect 36858 1719 36859 1775
rect 36801 1695 36804 1719
rect 36856 1695 36859 1719
rect 36801 1639 36802 1695
rect 36858 1639 36859 1695
rect 36801 1615 36804 1639
rect 36856 1615 36859 1639
rect 36801 1559 36802 1615
rect 36858 1559 36859 1615
rect 36801 1545 36804 1559
rect 36856 1545 36859 1559
rect 36801 1535 36859 1545
rect 36801 1479 36802 1535
rect 36858 1479 36859 1535
rect 36801 1469 36859 1479
rect 36801 1455 36804 1469
rect 36856 1455 36859 1469
rect 36801 1399 36802 1455
rect 36858 1399 36859 1455
rect 36801 1375 36804 1399
rect 36856 1375 36859 1399
rect 36801 1319 36802 1375
rect 36858 1319 36859 1375
rect 36801 1295 36804 1319
rect 36856 1295 36859 1319
rect 36801 1239 36802 1295
rect 36858 1239 36859 1295
rect 36801 1225 36804 1239
rect 36856 1225 36859 1239
rect 36801 1215 36859 1225
rect 36801 1159 36802 1215
rect 36858 1159 36859 1215
rect 36801 1147 36859 1159
rect 36897 3133 36955 3147
rect 36897 3081 36900 3133
rect 36952 3081 36955 3133
rect 36897 3069 36955 3081
rect 36897 3017 36900 3069
rect 36952 3017 36955 3069
rect 36897 3005 36955 3017
rect 36897 2953 36900 3005
rect 36952 2953 36955 3005
rect 36897 2941 36955 2953
rect 36897 2889 36900 2941
rect 36952 2889 36955 2941
rect 36897 2877 36955 2889
rect 36897 2825 36900 2877
rect 36952 2825 36955 2877
rect 36897 2813 36955 2825
rect 36897 2761 36900 2813
rect 36952 2761 36955 2813
rect 36897 2749 36955 2761
rect 36897 2697 36900 2749
rect 36952 2697 36955 2749
rect 36897 2685 36955 2697
rect 36897 2633 36900 2685
rect 36952 2633 36955 2685
rect 36897 2621 36955 2633
rect 36897 2569 36900 2621
rect 36952 2569 36955 2621
rect 36897 2557 36955 2569
rect 36897 2505 36900 2557
rect 36952 2505 36955 2557
rect 36897 2493 36955 2505
rect 36897 2441 36900 2493
rect 36952 2441 36955 2493
rect 36897 2429 36955 2441
rect 36897 2377 36900 2429
rect 36952 2377 36955 2429
rect 36897 2365 36955 2377
rect 36897 2313 36900 2365
rect 36952 2313 36955 2365
rect 36897 2301 36955 2313
rect 36897 2249 36900 2301
rect 36952 2249 36955 2301
rect 36897 2237 36955 2249
rect 36897 2185 36900 2237
rect 36952 2185 36955 2237
rect 36897 2173 36955 2185
rect 36897 2121 36900 2173
rect 36952 2121 36955 2173
rect 36897 2109 36955 2121
rect 36897 2057 36900 2109
rect 36952 2057 36955 2109
rect 36897 2045 36955 2057
rect 36897 1993 36900 2045
rect 36952 1993 36955 2045
rect 36897 1981 36955 1993
rect 36897 1929 36900 1981
rect 36952 1929 36955 1981
rect 36897 1917 36955 1929
rect 36897 1865 36900 1917
rect 36952 1865 36955 1917
rect 36897 1853 36955 1865
rect 36897 1801 36900 1853
rect 36952 1801 36955 1853
rect 36897 1789 36955 1801
rect 36897 1737 36900 1789
rect 36952 1737 36955 1789
rect 36897 1725 36955 1737
rect 36897 1673 36900 1725
rect 36952 1673 36955 1725
rect 36897 1661 36955 1673
rect 36897 1609 36900 1661
rect 36952 1609 36955 1661
rect 36897 1597 36955 1609
rect 36897 1545 36900 1597
rect 36952 1545 36955 1597
rect 36897 1533 36955 1545
rect 36897 1481 36900 1533
rect 36952 1481 36955 1533
rect 36897 1469 36955 1481
rect 36897 1417 36900 1469
rect 36952 1417 36955 1469
rect 36897 1405 36955 1417
rect 36897 1353 36900 1405
rect 36952 1353 36955 1405
rect 36897 1341 36955 1353
rect 36897 1289 36900 1341
rect 36952 1289 36955 1341
rect 36897 1277 36955 1289
rect 36897 1225 36900 1277
rect 36952 1225 36955 1277
rect 36897 1213 36955 1225
rect 36897 1161 36900 1213
rect 36952 1161 36955 1213
rect 36897 830 36955 1161
rect 36993 3135 37051 3147
rect 36993 3079 36994 3135
rect 37050 3079 37051 3135
rect 36993 3069 37051 3079
rect 36993 3055 36996 3069
rect 37048 3055 37051 3069
rect 36993 2999 36994 3055
rect 37050 2999 37051 3055
rect 36993 2975 36996 2999
rect 37048 2975 37051 2999
rect 36993 2919 36994 2975
rect 37050 2919 37051 2975
rect 36993 2895 36996 2919
rect 37048 2895 37051 2919
rect 36993 2839 36994 2895
rect 37050 2839 37051 2895
rect 36993 2825 36996 2839
rect 37048 2825 37051 2839
rect 36993 2815 37051 2825
rect 36993 2759 36994 2815
rect 37050 2759 37051 2815
rect 36993 2749 37051 2759
rect 36993 2735 36996 2749
rect 37048 2735 37051 2749
rect 36993 2679 36994 2735
rect 37050 2679 37051 2735
rect 36993 2655 36996 2679
rect 37048 2655 37051 2679
rect 36993 2599 36994 2655
rect 37050 2599 37051 2655
rect 36993 2575 36996 2599
rect 37048 2575 37051 2599
rect 36993 2519 36994 2575
rect 37050 2519 37051 2575
rect 36993 2505 36996 2519
rect 37048 2505 37051 2519
rect 36993 2495 37051 2505
rect 36993 2439 36994 2495
rect 37050 2439 37051 2495
rect 36993 2429 37051 2439
rect 36993 2415 36996 2429
rect 37048 2415 37051 2429
rect 36993 2359 36994 2415
rect 37050 2359 37051 2415
rect 36993 2335 36996 2359
rect 37048 2335 37051 2359
rect 36993 2279 36994 2335
rect 37050 2279 37051 2335
rect 36993 2255 36996 2279
rect 37048 2255 37051 2279
rect 36993 2199 36994 2255
rect 37050 2199 37051 2255
rect 36993 2185 36996 2199
rect 37048 2185 37051 2199
rect 36993 2175 37051 2185
rect 36993 2119 36994 2175
rect 37050 2119 37051 2175
rect 36993 2109 37051 2119
rect 36993 2095 36996 2109
rect 37048 2095 37051 2109
rect 36993 2039 36994 2095
rect 37050 2039 37051 2095
rect 36993 2015 36996 2039
rect 37048 2015 37051 2039
rect 36993 1959 36994 2015
rect 37050 1959 37051 2015
rect 36993 1935 36996 1959
rect 37048 1935 37051 1959
rect 36993 1879 36994 1935
rect 37050 1879 37051 1935
rect 36993 1865 36996 1879
rect 37048 1865 37051 1879
rect 36993 1855 37051 1865
rect 36993 1799 36994 1855
rect 37050 1799 37051 1855
rect 36993 1789 37051 1799
rect 36993 1775 36996 1789
rect 37048 1775 37051 1789
rect 36993 1719 36994 1775
rect 37050 1719 37051 1775
rect 36993 1695 36996 1719
rect 37048 1695 37051 1719
rect 36993 1639 36994 1695
rect 37050 1639 37051 1695
rect 36993 1615 36996 1639
rect 37048 1615 37051 1639
rect 36993 1559 36994 1615
rect 37050 1559 37051 1615
rect 36993 1545 36996 1559
rect 37048 1545 37051 1559
rect 36993 1535 37051 1545
rect 36993 1479 36994 1535
rect 37050 1479 37051 1535
rect 36993 1469 37051 1479
rect 36993 1455 36996 1469
rect 37048 1455 37051 1469
rect 36993 1399 36994 1455
rect 37050 1399 37051 1455
rect 36993 1375 36996 1399
rect 37048 1375 37051 1399
rect 36993 1319 36994 1375
rect 37050 1319 37051 1375
rect 36993 1295 36996 1319
rect 37048 1295 37051 1319
rect 36993 1239 36994 1295
rect 37050 1239 37051 1295
rect 36993 1225 36996 1239
rect 37048 1225 37051 1239
rect 36993 1215 37051 1225
rect 36993 1159 36994 1215
rect 37050 1159 37051 1215
rect 36993 1147 37051 1159
rect 37089 3133 37147 3147
rect 37089 3081 37092 3133
rect 37144 3081 37147 3133
rect 37089 3069 37147 3081
rect 37089 3017 37092 3069
rect 37144 3017 37147 3069
rect 37089 3005 37147 3017
rect 37089 2953 37092 3005
rect 37144 2953 37147 3005
rect 37089 2941 37147 2953
rect 37089 2889 37092 2941
rect 37144 2889 37147 2941
rect 37089 2877 37147 2889
rect 37089 2825 37092 2877
rect 37144 2825 37147 2877
rect 37089 2813 37147 2825
rect 37089 2761 37092 2813
rect 37144 2761 37147 2813
rect 37089 2749 37147 2761
rect 37089 2697 37092 2749
rect 37144 2697 37147 2749
rect 37089 2685 37147 2697
rect 37089 2633 37092 2685
rect 37144 2633 37147 2685
rect 37089 2621 37147 2633
rect 37089 2569 37092 2621
rect 37144 2569 37147 2621
rect 37089 2557 37147 2569
rect 37089 2505 37092 2557
rect 37144 2505 37147 2557
rect 37089 2493 37147 2505
rect 37089 2441 37092 2493
rect 37144 2441 37147 2493
rect 37089 2429 37147 2441
rect 37089 2377 37092 2429
rect 37144 2377 37147 2429
rect 37089 2365 37147 2377
rect 37089 2313 37092 2365
rect 37144 2313 37147 2365
rect 37089 2301 37147 2313
rect 37089 2249 37092 2301
rect 37144 2249 37147 2301
rect 37089 2237 37147 2249
rect 37089 2185 37092 2237
rect 37144 2185 37147 2237
rect 37089 2173 37147 2185
rect 37089 2121 37092 2173
rect 37144 2121 37147 2173
rect 37089 2109 37147 2121
rect 37089 2057 37092 2109
rect 37144 2057 37147 2109
rect 37089 2045 37147 2057
rect 37089 1993 37092 2045
rect 37144 1993 37147 2045
rect 37089 1981 37147 1993
rect 37089 1929 37092 1981
rect 37144 1929 37147 1981
rect 37089 1917 37147 1929
rect 37089 1865 37092 1917
rect 37144 1865 37147 1917
rect 37089 1853 37147 1865
rect 37089 1801 37092 1853
rect 37144 1801 37147 1853
rect 37089 1789 37147 1801
rect 37089 1737 37092 1789
rect 37144 1737 37147 1789
rect 37089 1725 37147 1737
rect 37089 1673 37092 1725
rect 37144 1673 37147 1725
rect 37089 1661 37147 1673
rect 37089 1609 37092 1661
rect 37144 1609 37147 1661
rect 37089 1597 37147 1609
rect 37089 1545 37092 1597
rect 37144 1545 37147 1597
rect 37089 1533 37147 1545
rect 37089 1481 37092 1533
rect 37144 1481 37147 1533
rect 37089 1469 37147 1481
rect 37089 1417 37092 1469
rect 37144 1417 37147 1469
rect 37089 1405 37147 1417
rect 37089 1353 37092 1405
rect 37144 1353 37147 1405
rect 37089 1341 37147 1353
rect 37089 1289 37092 1341
rect 37144 1289 37147 1341
rect 37089 1277 37147 1289
rect 37089 1225 37092 1277
rect 37144 1225 37147 1277
rect 37089 1213 37147 1225
rect 37089 1161 37092 1213
rect 37144 1161 37147 1213
rect 37089 830 37147 1161
rect 37185 3135 37243 3147
rect 37185 3079 37186 3135
rect 37242 3079 37243 3135
rect 37185 3069 37243 3079
rect 37185 3055 37188 3069
rect 37240 3055 37243 3069
rect 37185 2999 37186 3055
rect 37242 2999 37243 3055
rect 37185 2975 37188 2999
rect 37240 2975 37243 2999
rect 37185 2919 37186 2975
rect 37242 2919 37243 2975
rect 37185 2895 37188 2919
rect 37240 2895 37243 2919
rect 37185 2839 37186 2895
rect 37242 2839 37243 2895
rect 37185 2825 37188 2839
rect 37240 2825 37243 2839
rect 37185 2815 37243 2825
rect 37185 2759 37186 2815
rect 37242 2759 37243 2815
rect 37185 2749 37243 2759
rect 37185 2735 37188 2749
rect 37240 2735 37243 2749
rect 37185 2679 37186 2735
rect 37242 2679 37243 2735
rect 37185 2655 37188 2679
rect 37240 2655 37243 2679
rect 37185 2599 37186 2655
rect 37242 2599 37243 2655
rect 37185 2575 37188 2599
rect 37240 2575 37243 2599
rect 37185 2519 37186 2575
rect 37242 2519 37243 2575
rect 37185 2505 37188 2519
rect 37240 2505 37243 2519
rect 37185 2495 37243 2505
rect 37185 2439 37186 2495
rect 37242 2439 37243 2495
rect 37185 2429 37243 2439
rect 37185 2415 37188 2429
rect 37240 2415 37243 2429
rect 37185 2359 37186 2415
rect 37242 2359 37243 2415
rect 37185 2335 37188 2359
rect 37240 2335 37243 2359
rect 37185 2279 37186 2335
rect 37242 2279 37243 2335
rect 37185 2255 37188 2279
rect 37240 2255 37243 2279
rect 37185 2199 37186 2255
rect 37242 2199 37243 2255
rect 37185 2185 37188 2199
rect 37240 2185 37243 2199
rect 37185 2175 37243 2185
rect 37185 2119 37186 2175
rect 37242 2119 37243 2175
rect 37185 2109 37243 2119
rect 37185 2095 37188 2109
rect 37240 2095 37243 2109
rect 37185 2039 37186 2095
rect 37242 2039 37243 2095
rect 37185 2015 37188 2039
rect 37240 2015 37243 2039
rect 37185 1959 37186 2015
rect 37242 1959 37243 2015
rect 37185 1935 37188 1959
rect 37240 1935 37243 1959
rect 37185 1879 37186 1935
rect 37242 1879 37243 1935
rect 37185 1865 37188 1879
rect 37240 1865 37243 1879
rect 37185 1855 37243 1865
rect 37185 1799 37186 1855
rect 37242 1799 37243 1855
rect 37185 1789 37243 1799
rect 37185 1775 37188 1789
rect 37240 1775 37243 1789
rect 37185 1719 37186 1775
rect 37242 1719 37243 1775
rect 37185 1695 37188 1719
rect 37240 1695 37243 1719
rect 37185 1639 37186 1695
rect 37242 1639 37243 1695
rect 37185 1615 37188 1639
rect 37240 1615 37243 1639
rect 37185 1559 37186 1615
rect 37242 1559 37243 1615
rect 37185 1545 37188 1559
rect 37240 1545 37243 1559
rect 37185 1535 37243 1545
rect 37185 1479 37186 1535
rect 37242 1479 37243 1535
rect 37185 1469 37243 1479
rect 37185 1455 37188 1469
rect 37240 1455 37243 1469
rect 37185 1399 37186 1455
rect 37242 1399 37243 1455
rect 37185 1375 37188 1399
rect 37240 1375 37243 1399
rect 37185 1319 37186 1375
rect 37242 1319 37243 1375
rect 37185 1295 37188 1319
rect 37240 1295 37243 1319
rect 37185 1239 37186 1295
rect 37242 1239 37243 1295
rect 37185 1225 37188 1239
rect 37240 1225 37243 1239
rect 37185 1215 37243 1225
rect 37185 1159 37186 1215
rect 37242 1159 37243 1215
rect 37185 1147 37243 1159
rect 37281 3133 37339 3147
rect 37281 3081 37284 3133
rect 37336 3081 37339 3133
rect 37281 3069 37339 3081
rect 37281 3017 37284 3069
rect 37336 3017 37339 3069
rect 37281 3005 37339 3017
rect 37281 2953 37284 3005
rect 37336 2953 37339 3005
rect 37281 2941 37339 2953
rect 37281 2889 37284 2941
rect 37336 2889 37339 2941
rect 37281 2877 37339 2889
rect 37281 2825 37284 2877
rect 37336 2825 37339 2877
rect 37281 2813 37339 2825
rect 37281 2761 37284 2813
rect 37336 2761 37339 2813
rect 37281 2749 37339 2761
rect 37281 2697 37284 2749
rect 37336 2697 37339 2749
rect 37281 2685 37339 2697
rect 37281 2633 37284 2685
rect 37336 2633 37339 2685
rect 37281 2621 37339 2633
rect 37281 2569 37284 2621
rect 37336 2569 37339 2621
rect 37281 2557 37339 2569
rect 37281 2505 37284 2557
rect 37336 2505 37339 2557
rect 37281 2493 37339 2505
rect 37281 2441 37284 2493
rect 37336 2441 37339 2493
rect 37281 2429 37339 2441
rect 37281 2377 37284 2429
rect 37336 2377 37339 2429
rect 37281 2365 37339 2377
rect 37281 2313 37284 2365
rect 37336 2313 37339 2365
rect 37281 2301 37339 2313
rect 37281 2249 37284 2301
rect 37336 2249 37339 2301
rect 37281 2237 37339 2249
rect 37281 2185 37284 2237
rect 37336 2185 37339 2237
rect 37281 2173 37339 2185
rect 37281 2121 37284 2173
rect 37336 2121 37339 2173
rect 37281 2109 37339 2121
rect 37281 2057 37284 2109
rect 37336 2057 37339 2109
rect 37281 2045 37339 2057
rect 37281 1993 37284 2045
rect 37336 1993 37339 2045
rect 37281 1981 37339 1993
rect 37281 1929 37284 1981
rect 37336 1929 37339 1981
rect 37281 1917 37339 1929
rect 37281 1865 37284 1917
rect 37336 1865 37339 1917
rect 37281 1853 37339 1865
rect 37281 1801 37284 1853
rect 37336 1801 37339 1853
rect 37281 1789 37339 1801
rect 37281 1737 37284 1789
rect 37336 1737 37339 1789
rect 37281 1725 37339 1737
rect 37281 1673 37284 1725
rect 37336 1673 37339 1725
rect 37281 1661 37339 1673
rect 37281 1609 37284 1661
rect 37336 1609 37339 1661
rect 37281 1597 37339 1609
rect 37281 1545 37284 1597
rect 37336 1545 37339 1597
rect 37281 1533 37339 1545
rect 37281 1481 37284 1533
rect 37336 1481 37339 1533
rect 37281 1469 37339 1481
rect 37281 1417 37284 1469
rect 37336 1417 37339 1469
rect 37281 1405 37339 1417
rect 37281 1353 37284 1405
rect 37336 1353 37339 1405
rect 37281 1341 37339 1353
rect 37281 1289 37284 1341
rect 37336 1289 37339 1341
rect 37281 1277 37339 1289
rect 37281 1225 37284 1277
rect 37336 1225 37339 1277
rect 37281 1213 37339 1225
rect 37281 1161 37284 1213
rect 37336 1161 37339 1213
rect 37281 830 37339 1161
rect 37377 3135 37435 3147
rect 37377 3079 37378 3135
rect 37434 3079 37435 3135
rect 37377 3069 37435 3079
rect 37377 3055 37380 3069
rect 37432 3055 37435 3069
rect 37377 2999 37378 3055
rect 37434 2999 37435 3055
rect 37377 2975 37380 2999
rect 37432 2975 37435 2999
rect 37377 2919 37378 2975
rect 37434 2919 37435 2975
rect 37377 2895 37380 2919
rect 37432 2895 37435 2919
rect 37377 2839 37378 2895
rect 37434 2839 37435 2895
rect 37377 2825 37380 2839
rect 37432 2825 37435 2839
rect 37377 2815 37435 2825
rect 37377 2759 37378 2815
rect 37434 2759 37435 2815
rect 37377 2749 37435 2759
rect 37377 2735 37380 2749
rect 37432 2735 37435 2749
rect 37377 2679 37378 2735
rect 37434 2679 37435 2735
rect 37377 2655 37380 2679
rect 37432 2655 37435 2679
rect 37377 2599 37378 2655
rect 37434 2599 37435 2655
rect 37377 2575 37380 2599
rect 37432 2575 37435 2599
rect 37377 2519 37378 2575
rect 37434 2519 37435 2575
rect 37377 2505 37380 2519
rect 37432 2505 37435 2519
rect 37377 2495 37435 2505
rect 37377 2439 37378 2495
rect 37434 2439 37435 2495
rect 37377 2429 37435 2439
rect 37377 2415 37380 2429
rect 37432 2415 37435 2429
rect 37377 2359 37378 2415
rect 37434 2359 37435 2415
rect 37377 2335 37380 2359
rect 37432 2335 37435 2359
rect 37377 2279 37378 2335
rect 37434 2279 37435 2335
rect 37377 2255 37380 2279
rect 37432 2255 37435 2279
rect 37377 2199 37378 2255
rect 37434 2199 37435 2255
rect 37377 2185 37380 2199
rect 37432 2185 37435 2199
rect 37377 2175 37435 2185
rect 37377 2119 37378 2175
rect 37434 2119 37435 2175
rect 37377 2109 37435 2119
rect 37377 2095 37380 2109
rect 37432 2095 37435 2109
rect 37377 2039 37378 2095
rect 37434 2039 37435 2095
rect 37377 2015 37380 2039
rect 37432 2015 37435 2039
rect 37377 1959 37378 2015
rect 37434 1959 37435 2015
rect 37377 1935 37380 1959
rect 37432 1935 37435 1959
rect 37377 1879 37378 1935
rect 37434 1879 37435 1935
rect 37377 1865 37380 1879
rect 37432 1865 37435 1879
rect 37377 1855 37435 1865
rect 37377 1799 37378 1855
rect 37434 1799 37435 1855
rect 37377 1789 37435 1799
rect 37377 1775 37380 1789
rect 37432 1775 37435 1789
rect 37377 1719 37378 1775
rect 37434 1719 37435 1775
rect 37377 1695 37380 1719
rect 37432 1695 37435 1719
rect 37377 1639 37378 1695
rect 37434 1639 37435 1695
rect 37377 1615 37380 1639
rect 37432 1615 37435 1639
rect 37377 1559 37378 1615
rect 37434 1559 37435 1615
rect 37377 1545 37380 1559
rect 37432 1545 37435 1559
rect 37377 1535 37435 1545
rect 37377 1479 37378 1535
rect 37434 1479 37435 1535
rect 37377 1469 37435 1479
rect 37377 1455 37380 1469
rect 37432 1455 37435 1469
rect 37377 1399 37378 1455
rect 37434 1399 37435 1455
rect 37377 1375 37380 1399
rect 37432 1375 37435 1399
rect 37377 1319 37378 1375
rect 37434 1319 37435 1375
rect 37377 1295 37380 1319
rect 37432 1295 37435 1319
rect 37377 1239 37378 1295
rect 37434 1239 37435 1295
rect 37377 1225 37380 1239
rect 37432 1225 37435 1239
rect 37377 1215 37435 1225
rect 37377 1159 37378 1215
rect 37434 1159 37435 1215
rect 37377 1147 37435 1159
rect 37473 3133 37531 3147
rect 37473 3081 37476 3133
rect 37528 3081 37531 3133
rect 37473 3069 37531 3081
rect 37473 3017 37476 3069
rect 37528 3017 37531 3069
rect 37473 3005 37531 3017
rect 37473 2953 37476 3005
rect 37528 2953 37531 3005
rect 37473 2941 37531 2953
rect 37473 2889 37476 2941
rect 37528 2889 37531 2941
rect 37473 2877 37531 2889
rect 37473 2825 37476 2877
rect 37528 2825 37531 2877
rect 37473 2813 37531 2825
rect 37473 2761 37476 2813
rect 37528 2761 37531 2813
rect 37473 2749 37531 2761
rect 37473 2697 37476 2749
rect 37528 2697 37531 2749
rect 37473 2685 37531 2697
rect 37473 2633 37476 2685
rect 37528 2633 37531 2685
rect 37473 2621 37531 2633
rect 37473 2569 37476 2621
rect 37528 2569 37531 2621
rect 37473 2557 37531 2569
rect 37473 2505 37476 2557
rect 37528 2505 37531 2557
rect 37473 2493 37531 2505
rect 37473 2441 37476 2493
rect 37528 2441 37531 2493
rect 37473 2429 37531 2441
rect 37473 2377 37476 2429
rect 37528 2377 37531 2429
rect 37473 2365 37531 2377
rect 37473 2313 37476 2365
rect 37528 2313 37531 2365
rect 37473 2301 37531 2313
rect 37473 2249 37476 2301
rect 37528 2249 37531 2301
rect 37473 2237 37531 2249
rect 37473 2185 37476 2237
rect 37528 2185 37531 2237
rect 37473 2173 37531 2185
rect 37473 2121 37476 2173
rect 37528 2121 37531 2173
rect 37473 2109 37531 2121
rect 37473 2057 37476 2109
rect 37528 2057 37531 2109
rect 37473 2045 37531 2057
rect 37473 1993 37476 2045
rect 37528 1993 37531 2045
rect 37473 1981 37531 1993
rect 37473 1929 37476 1981
rect 37528 1929 37531 1981
rect 37473 1917 37531 1929
rect 37473 1865 37476 1917
rect 37528 1865 37531 1917
rect 37473 1853 37531 1865
rect 37473 1801 37476 1853
rect 37528 1801 37531 1853
rect 37473 1789 37531 1801
rect 37473 1737 37476 1789
rect 37528 1737 37531 1789
rect 37473 1725 37531 1737
rect 37473 1673 37476 1725
rect 37528 1673 37531 1725
rect 37473 1661 37531 1673
rect 37473 1609 37476 1661
rect 37528 1609 37531 1661
rect 37473 1597 37531 1609
rect 37473 1545 37476 1597
rect 37528 1545 37531 1597
rect 37473 1533 37531 1545
rect 37473 1481 37476 1533
rect 37528 1481 37531 1533
rect 37473 1469 37531 1481
rect 37473 1417 37476 1469
rect 37528 1417 37531 1469
rect 37473 1405 37531 1417
rect 37473 1353 37476 1405
rect 37528 1353 37531 1405
rect 37473 1341 37531 1353
rect 37473 1289 37476 1341
rect 37528 1289 37531 1341
rect 37473 1277 37531 1289
rect 37473 1225 37476 1277
rect 37528 1225 37531 1277
rect 37473 1213 37531 1225
rect 37473 1161 37476 1213
rect 37528 1161 37531 1213
rect 37473 830 37531 1161
rect 37569 3135 37627 3147
rect 37569 3079 37570 3135
rect 37626 3079 37627 3135
rect 37569 3069 37627 3079
rect 37569 3055 37572 3069
rect 37624 3055 37627 3069
rect 37569 2999 37570 3055
rect 37626 2999 37627 3055
rect 37569 2975 37572 2999
rect 37624 2975 37627 2999
rect 37569 2919 37570 2975
rect 37626 2919 37627 2975
rect 37569 2895 37572 2919
rect 37624 2895 37627 2919
rect 37569 2839 37570 2895
rect 37626 2839 37627 2895
rect 37569 2825 37572 2839
rect 37624 2825 37627 2839
rect 37569 2815 37627 2825
rect 37569 2759 37570 2815
rect 37626 2759 37627 2815
rect 37569 2749 37627 2759
rect 37569 2735 37572 2749
rect 37624 2735 37627 2749
rect 37569 2679 37570 2735
rect 37626 2679 37627 2735
rect 37569 2655 37572 2679
rect 37624 2655 37627 2679
rect 37569 2599 37570 2655
rect 37626 2599 37627 2655
rect 37569 2575 37572 2599
rect 37624 2575 37627 2599
rect 37569 2519 37570 2575
rect 37626 2519 37627 2575
rect 37569 2505 37572 2519
rect 37624 2505 37627 2519
rect 37569 2495 37627 2505
rect 37569 2439 37570 2495
rect 37626 2439 37627 2495
rect 37569 2429 37627 2439
rect 37569 2415 37572 2429
rect 37624 2415 37627 2429
rect 37569 2359 37570 2415
rect 37626 2359 37627 2415
rect 37569 2335 37572 2359
rect 37624 2335 37627 2359
rect 37569 2279 37570 2335
rect 37626 2279 37627 2335
rect 37569 2255 37572 2279
rect 37624 2255 37627 2279
rect 37569 2199 37570 2255
rect 37626 2199 37627 2255
rect 37569 2185 37572 2199
rect 37624 2185 37627 2199
rect 37569 2175 37627 2185
rect 37569 2119 37570 2175
rect 37626 2119 37627 2175
rect 37569 2109 37627 2119
rect 37569 2095 37572 2109
rect 37624 2095 37627 2109
rect 37569 2039 37570 2095
rect 37626 2039 37627 2095
rect 37569 2015 37572 2039
rect 37624 2015 37627 2039
rect 37569 1959 37570 2015
rect 37626 1959 37627 2015
rect 37569 1935 37572 1959
rect 37624 1935 37627 1959
rect 37569 1879 37570 1935
rect 37626 1879 37627 1935
rect 37569 1865 37572 1879
rect 37624 1865 37627 1879
rect 37569 1855 37627 1865
rect 37569 1799 37570 1855
rect 37626 1799 37627 1855
rect 37569 1789 37627 1799
rect 37569 1775 37572 1789
rect 37624 1775 37627 1789
rect 37569 1719 37570 1775
rect 37626 1719 37627 1775
rect 37569 1695 37572 1719
rect 37624 1695 37627 1719
rect 37569 1639 37570 1695
rect 37626 1639 37627 1695
rect 37569 1615 37572 1639
rect 37624 1615 37627 1639
rect 37569 1559 37570 1615
rect 37626 1559 37627 1615
rect 37569 1545 37572 1559
rect 37624 1545 37627 1559
rect 37569 1535 37627 1545
rect 37569 1479 37570 1535
rect 37626 1479 37627 1535
rect 37569 1469 37627 1479
rect 37569 1455 37572 1469
rect 37624 1455 37627 1469
rect 37569 1399 37570 1455
rect 37626 1399 37627 1455
rect 37569 1375 37572 1399
rect 37624 1375 37627 1399
rect 37569 1319 37570 1375
rect 37626 1319 37627 1375
rect 37569 1295 37572 1319
rect 37624 1295 37627 1319
rect 37569 1239 37570 1295
rect 37626 1239 37627 1295
rect 37569 1225 37572 1239
rect 37624 1225 37627 1239
rect 37569 1215 37627 1225
rect 37569 1159 37570 1215
rect 37626 1159 37627 1215
rect 37569 1147 37627 1159
rect 37665 3133 37723 3147
rect 37665 3081 37668 3133
rect 37720 3081 37723 3133
rect 37665 3069 37723 3081
rect 37665 3017 37668 3069
rect 37720 3017 37723 3069
rect 37665 3005 37723 3017
rect 37665 2953 37668 3005
rect 37720 2953 37723 3005
rect 37665 2941 37723 2953
rect 37665 2889 37668 2941
rect 37720 2889 37723 2941
rect 37665 2877 37723 2889
rect 37665 2825 37668 2877
rect 37720 2825 37723 2877
rect 37665 2813 37723 2825
rect 37665 2761 37668 2813
rect 37720 2761 37723 2813
rect 37665 2749 37723 2761
rect 37665 2697 37668 2749
rect 37720 2697 37723 2749
rect 37665 2685 37723 2697
rect 37665 2633 37668 2685
rect 37720 2633 37723 2685
rect 37665 2621 37723 2633
rect 37665 2569 37668 2621
rect 37720 2569 37723 2621
rect 37665 2557 37723 2569
rect 37665 2505 37668 2557
rect 37720 2505 37723 2557
rect 37665 2493 37723 2505
rect 37665 2441 37668 2493
rect 37720 2441 37723 2493
rect 37665 2429 37723 2441
rect 37665 2377 37668 2429
rect 37720 2377 37723 2429
rect 37665 2365 37723 2377
rect 37665 2313 37668 2365
rect 37720 2313 37723 2365
rect 37665 2301 37723 2313
rect 37665 2249 37668 2301
rect 37720 2249 37723 2301
rect 37665 2237 37723 2249
rect 37665 2185 37668 2237
rect 37720 2185 37723 2237
rect 37665 2173 37723 2185
rect 37665 2121 37668 2173
rect 37720 2121 37723 2173
rect 37665 2109 37723 2121
rect 37665 2057 37668 2109
rect 37720 2057 37723 2109
rect 37665 2045 37723 2057
rect 37665 1993 37668 2045
rect 37720 1993 37723 2045
rect 37665 1981 37723 1993
rect 37665 1929 37668 1981
rect 37720 1929 37723 1981
rect 37665 1917 37723 1929
rect 37665 1865 37668 1917
rect 37720 1865 37723 1917
rect 37665 1853 37723 1865
rect 37665 1801 37668 1853
rect 37720 1801 37723 1853
rect 37665 1789 37723 1801
rect 37665 1737 37668 1789
rect 37720 1737 37723 1789
rect 37665 1725 37723 1737
rect 37665 1673 37668 1725
rect 37720 1673 37723 1725
rect 37665 1661 37723 1673
rect 37665 1609 37668 1661
rect 37720 1609 37723 1661
rect 37665 1597 37723 1609
rect 37665 1545 37668 1597
rect 37720 1545 37723 1597
rect 37665 1533 37723 1545
rect 37665 1481 37668 1533
rect 37720 1481 37723 1533
rect 37665 1469 37723 1481
rect 37665 1417 37668 1469
rect 37720 1417 37723 1469
rect 37665 1405 37723 1417
rect 37665 1353 37668 1405
rect 37720 1353 37723 1405
rect 37665 1341 37723 1353
rect 37665 1289 37668 1341
rect 37720 1289 37723 1341
rect 37665 1277 37723 1289
rect 37665 1225 37668 1277
rect 37720 1225 37723 1277
rect 37665 1213 37723 1225
rect 37665 1161 37668 1213
rect 37720 1161 37723 1213
rect 37665 830 37723 1161
rect 37761 3135 37819 3147
rect 37761 3079 37762 3135
rect 37818 3079 37819 3135
rect 37761 3069 37819 3079
rect 37761 3055 37764 3069
rect 37816 3055 37819 3069
rect 37761 2999 37762 3055
rect 37818 2999 37819 3055
rect 37761 2975 37764 2999
rect 37816 2975 37819 2999
rect 37761 2919 37762 2975
rect 37818 2919 37819 2975
rect 37761 2895 37764 2919
rect 37816 2895 37819 2919
rect 37761 2839 37762 2895
rect 37818 2839 37819 2895
rect 37761 2825 37764 2839
rect 37816 2825 37819 2839
rect 37761 2815 37819 2825
rect 37761 2759 37762 2815
rect 37818 2759 37819 2815
rect 37761 2749 37819 2759
rect 37761 2735 37764 2749
rect 37816 2735 37819 2749
rect 37761 2679 37762 2735
rect 37818 2679 37819 2735
rect 37761 2655 37764 2679
rect 37816 2655 37819 2679
rect 37761 2599 37762 2655
rect 37818 2599 37819 2655
rect 37761 2575 37764 2599
rect 37816 2575 37819 2599
rect 37761 2519 37762 2575
rect 37818 2519 37819 2575
rect 37761 2505 37764 2519
rect 37816 2505 37819 2519
rect 37761 2495 37819 2505
rect 37761 2439 37762 2495
rect 37818 2439 37819 2495
rect 37761 2429 37819 2439
rect 37761 2415 37764 2429
rect 37816 2415 37819 2429
rect 37761 2359 37762 2415
rect 37818 2359 37819 2415
rect 37761 2335 37764 2359
rect 37816 2335 37819 2359
rect 37761 2279 37762 2335
rect 37818 2279 37819 2335
rect 37761 2255 37764 2279
rect 37816 2255 37819 2279
rect 37761 2199 37762 2255
rect 37818 2199 37819 2255
rect 37761 2185 37764 2199
rect 37816 2185 37819 2199
rect 37761 2175 37819 2185
rect 37761 2119 37762 2175
rect 37818 2119 37819 2175
rect 37761 2109 37819 2119
rect 37761 2095 37764 2109
rect 37816 2095 37819 2109
rect 37761 2039 37762 2095
rect 37818 2039 37819 2095
rect 37761 2015 37764 2039
rect 37816 2015 37819 2039
rect 37761 1959 37762 2015
rect 37818 1959 37819 2015
rect 37761 1935 37764 1959
rect 37816 1935 37819 1959
rect 37761 1879 37762 1935
rect 37818 1879 37819 1935
rect 37761 1865 37764 1879
rect 37816 1865 37819 1879
rect 37761 1855 37819 1865
rect 37761 1799 37762 1855
rect 37818 1799 37819 1855
rect 37761 1789 37819 1799
rect 37761 1775 37764 1789
rect 37816 1775 37819 1789
rect 37761 1719 37762 1775
rect 37818 1719 37819 1775
rect 37761 1695 37764 1719
rect 37816 1695 37819 1719
rect 37761 1639 37762 1695
rect 37818 1639 37819 1695
rect 37761 1615 37764 1639
rect 37816 1615 37819 1639
rect 37761 1559 37762 1615
rect 37818 1559 37819 1615
rect 37761 1545 37764 1559
rect 37816 1545 37819 1559
rect 37761 1535 37819 1545
rect 37761 1479 37762 1535
rect 37818 1479 37819 1535
rect 37761 1469 37819 1479
rect 37761 1455 37764 1469
rect 37816 1455 37819 1469
rect 37761 1399 37762 1455
rect 37818 1399 37819 1455
rect 37761 1375 37764 1399
rect 37816 1375 37819 1399
rect 37761 1319 37762 1375
rect 37818 1319 37819 1375
rect 37761 1295 37764 1319
rect 37816 1295 37819 1319
rect 37761 1239 37762 1295
rect 37818 1239 37819 1295
rect 37761 1225 37764 1239
rect 37816 1225 37819 1239
rect 37761 1215 37819 1225
rect 37761 1159 37762 1215
rect 37818 1159 37819 1215
rect 37761 1147 37819 1159
rect 37857 3133 37915 3147
rect 37857 3081 37860 3133
rect 37912 3081 37915 3133
rect 37857 3069 37915 3081
rect 37857 3017 37860 3069
rect 37912 3017 37915 3069
rect 37857 3005 37915 3017
rect 37857 2953 37860 3005
rect 37912 2953 37915 3005
rect 37857 2941 37915 2953
rect 37857 2889 37860 2941
rect 37912 2889 37915 2941
rect 37857 2877 37915 2889
rect 37857 2825 37860 2877
rect 37912 2825 37915 2877
rect 37857 2813 37915 2825
rect 37857 2761 37860 2813
rect 37912 2761 37915 2813
rect 37857 2749 37915 2761
rect 37857 2697 37860 2749
rect 37912 2697 37915 2749
rect 37857 2685 37915 2697
rect 37857 2633 37860 2685
rect 37912 2633 37915 2685
rect 37857 2621 37915 2633
rect 37857 2569 37860 2621
rect 37912 2569 37915 2621
rect 37857 2557 37915 2569
rect 37857 2505 37860 2557
rect 37912 2505 37915 2557
rect 37857 2493 37915 2505
rect 37857 2441 37860 2493
rect 37912 2441 37915 2493
rect 37857 2429 37915 2441
rect 37857 2377 37860 2429
rect 37912 2377 37915 2429
rect 37857 2365 37915 2377
rect 37857 2313 37860 2365
rect 37912 2313 37915 2365
rect 37857 2301 37915 2313
rect 37857 2249 37860 2301
rect 37912 2249 37915 2301
rect 37857 2237 37915 2249
rect 37857 2185 37860 2237
rect 37912 2185 37915 2237
rect 37857 2173 37915 2185
rect 37857 2121 37860 2173
rect 37912 2121 37915 2173
rect 37857 2109 37915 2121
rect 37857 2057 37860 2109
rect 37912 2057 37915 2109
rect 37857 2045 37915 2057
rect 37857 1993 37860 2045
rect 37912 1993 37915 2045
rect 37857 1981 37915 1993
rect 37857 1929 37860 1981
rect 37912 1929 37915 1981
rect 37857 1917 37915 1929
rect 37857 1865 37860 1917
rect 37912 1865 37915 1917
rect 37857 1853 37915 1865
rect 37857 1801 37860 1853
rect 37912 1801 37915 1853
rect 37857 1789 37915 1801
rect 37857 1737 37860 1789
rect 37912 1737 37915 1789
rect 37857 1725 37915 1737
rect 37857 1673 37860 1725
rect 37912 1673 37915 1725
rect 37857 1661 37915 1673
rect 37857 1609 37860 1661
rect 37912 1609 37915 1661
rect 37857 1597 37915 1609
rect 37857 1545 37860 1597
rect 37912 1545 37915 1597
rect 37857 1533 37915 1545
rect 37857 1481 37860 1533
rect 37912 1481 37915 1533
rect 37857 1469 37915 1481
rect 37857 1417 37860 1469
rect 37912 1417 37915 1469
rect 37857 1405 37915 1417
rect 37857 1353 37860 1405
rect 37912 1353 37915 1405
rect 37857 1341 37915 1353
rect 37857 1289 37860 1341
rect 37912 1289 37915 1341
rect 37857 1277 37915 1289
rect 37857 1225 37860 1277
rect 37912 1225 37915 1277
rect 37857 1213 37915 1225
rect 37857 1161 37860 1213
rect 37912 1161 37915 1213
rect 37857 830 37915 1161
rect 37953 3135 38011 3147
rect 37953 3079 37954 3135
rect 38010 3079 38011 3135
rect 37953 3069 38011 3079
rect 37953 3055 37956 3069
rect 38008 3055 38011 3069
rect 37953 2999 37954 3055
rect 38010 2999 38011 3055
rect 37953 2975 37956 2999
rect 38008 2975 38011 2999
rect 37953 2919 37954 2975
rect 38010 2919 38011 2975
rect 37953 2895 37956 2919
rect 38008 2895 38011 2919
rect 37953 2839 37954 2895
rect 38010 2839 38011 2895
rect 37953 2825 37956 2839
rect 38008 2825 38011 2839
rect 37953 2815 38011 2825
rect 37953 2759 37954 2815
rect 38010 2759 38011 2815
rect 37953 2749 38011 2759
rect 37953 2735 37956 2749
rect 38008 2735 38011 2749
rect 37953 2679 37954 2735
rect 38010 2679 38011 2735
rect 37953 2655 37956 2679
rect 38008 2655 38011 2679
rect 37953 2599 37954 2655
rect 38010 2599 38011 2655
rect 37953 2575 37956 2599
rect 38008 2575 38011 2599
rect 37953 2519 37954 2575
rect 38010 2519 38011 2575
rect 37953 2505 37956 2519
rect 38008 2505 38011 2519
rect 37953 2495 38011 2505
rect 37953 2439 37954 2495
rect 38010 2439 38011 2495
rect 37953 2429 38011 2439
rect 37953 2415 37956 2429
rect 38008 2415 38011 2429
rect 37953 2359 37954 2415
rect 38010 2359 38011 2415
rect 37953 2335 37956 2359
rect 38008 2335 38011 2359
rect 37953 2279 37954 2335
rect 38010 2279 38011 2335
rect 37953 2255 37956 2279
rect 38008 2255 38011 2279
rect 37953 2199 37954 2255
rect 38010 2199 38011 2255
rect 37953 2185 37956 2199
rect 38008 2185 38011 2199
rect 37953 2175 38011 2185
rect 37953 2119 37954 2175
rect 38010 2119 38011 2175
rect 37953 2109 38011 2119
rect 37953 2095 37956 2109
rect 38008 2095 38011 2109
rect 37953 2039 37954 2095
rect 38010 2039 38011 2095
rect 37953 2015 37956 2039
rect 38008 2015 38011 2039
rect 37953 1959 37954 2015
rect 38010 1959 38011 2015
rect 37953 1935 37956 1959
rect 38008 1935 38011 1959
rect 37953 1879 37954 1935
rect 38010 1879 38011 1935
rect 37953 1865 37956 1879
rect 38008 1865 38011 1879
rect 37953 1855 38011 1865
rect 37953 1799 37954 1855
rect 38010 1799 38011 1855
rect 37953 1789 38011 1799
rect 37953 1775 37956 1789
rect 38008 1775 38011 1789
rect 37953 1719 37954 1775
rect 38010 1719 38011 1775
rect 37953 1695 37956 1719
rect 38008 1695 38011 1719
rect 37953 1639 37954 1695
rect 38010 1639 38011 1695
rect 37953 1615 37956 1639
rect 38008 1615 38011 1639
rect 37953 1559 37954 1615
rect 38010 1559 38011 1615
rect 37953 1545 37956 1559
rect 38008 1545 38011 1559
rect 37953 1535 38011 1545
rect 37953 1479 37954 1535
rect 38010 1479 38011 1535
rect 37953 1469 38011 1479
rect 37953 1455 37956 1469
rect 38008 1455 38011 1469
rect 37953 1399 37954 1455
rect 38010 1399 38011 1455
rect 37953 1375 37956 1399
rect 38008 1375 38011 1399
rect 37953 1319 37954 1375
rect 38010 1319 38011 1375
rect 37953 1295 37956 1319
rect 38008 1295 38011 1319
rect 37953 1239 37954 1295
rect 38010 1239 38011 1295
rect 37953 1225 37956 1239
rect 38008 1225 38011 1239
rect 37953 1215 38011 1225
rect 37953 1159 37954 1215
rect 38010 1159 38011 1215
rect 37953 1147 38011 1159
rect 38049 3133 38107 3147
rect 38049 3081 38052 3133
rect 38104 3081 38107 3133
rect 38049 3069 38107 3081
rect 38049 3017 38052 3069
rect 38104 3017 38107 3069
rect 38049 3005 38107 3017
rect 38049 2953 38052 3005
rect 38104 2953 38107 3005
rect 38049 2941 38107 2953
rect 38049 2889 38052 2941
rect 38104 2889 38107 2941
rect 38049 2877 38107 2889
rect 38049 2825 38052 2877
rect 38104 2825 38107 2877
rect 38049 2813 38107 2825
rect 38049 2761 38052 2813
rect 38104 2761 38107 2813
rect 38049 2749 38107 2761
rect 38049 2697 38052 2749
rect 38104 2697 38107 2749
rect 38049 2685 38107 2697
rect 38049 2633 38052 2685
rect 38104 2633 38107 2685
rect 38049 2621 38107 2633
rect 38049 2569 38052 2621
rect 38104 2569 38107 2621
rect 38049 2557 38107 2569
rect 38049 2505 38052 2557
rect 38104 2505 38107 2557
rect 38049 2493 38107 2505
rect 38049 2441 38052 2493
rect 38104 2441 38107 2493
rect 38049 2429 38107 2441
rect 38049 2377 38052 2429
rect 38104 2377 38107 2429
rect 38049 2365 38107 2377
rect 38049 2313 38052 2365
rect 38104 2313 38107 2365
rect 38049 2301 38107 2313
rect 38049 2249 38052 2301
rect 38104 2249 38107 2301
rect 38049 2237 38107 2249
rect 38049 2185 38052 2237
rect 38104 2185 38107 2237
rect 38049 2173 38107 2185
rect 38049 2121 38052 2173
rect 38104 2121 38107 2173
rect 38049 2109 38107 2121
rect 38049 2057 38052 2109
rect 38104 2057 38107 2109
rect 38049 2045 38107 2057
rect 38049 1993 38052 2045
rect 38104 1993 38107 2045
rect 38049 1981 38107 1993
rect 38049 1929 38052 1981
rect 38104 1929 38107 1981
rect 38049 1917 38107 1929
rect 38049 1865 38052 1917
rect 38104 1865 38107 1917
rect 38049 1853 38107 1865
rect 38049 1801 38052 1853
rect 38104 1801 38107 1853
rect 38049 1789 38107 1801
rect 38049 1737 38052 1789
rect 38104 1737 38107 1789
rect 38049 1725 38107 1737
rect 38049 1673 38052 1725
rect 38104 1673 38107 1725
rect 38049 1661 38107 1673
rect 38049 1609 38052 1661
rect 38104 1609 38107 1661
rect 38049 1597 38107 1609
rect 38049 1545 38052 1597
rect 38104 1545 38107 1597
rect 38049 1533 38107 1545
rect 38049 1481 38052 1533
rect 38104 1481 38107 1533
rect 38049 1469 38107 1481
rect 38049 1417 38052 1469
rect 38104 1417 38107 1469
rect 38049 1405 38107 1417
rect 38049 1353 38052 1405
rect 38104 1353 38107 1405
rect 38049 1341 38107 1353
rect 38049 1289 38052 1341
rect 38104 1289 38107 1341
rect 38049 1277 38107 1289
rect 38049 1225 38052 1277
rect 38104 1225 38107 1277
rect 38049 1213 38107 1225
rect 38049 1161 38052 1213
rect 38104 1161 38107 1213
rect 38049 830 38107 1161
rect 38145 3135 38203 3147
rect 38145 3079 38146 3135
rect 38202 3079 38203 3135
rect 38145 3069 38203 3079
rect 38145 3055 38148 3069
rect 38200 3055 38203 3069
rect 38145 2999 38146 3055
rect 38202 2999 38203 3055
rect 38145 2975 38148 2999
rect 38200 2975 38203 2999
rect 38145 2919 38146 2975
rect 38202 2919 38203 2975
rect 38145 2895 38148 2919
rect 38200 2895 38203 2919
rect 38145 2839 38146 2895
rect 38202 2839 38203 2895
rect 38145 2825 38148 2839
rect 38200 2825 38203 2839
rect 38145 2815 38203 2825
rect 38145 2759 38146 2815
rect 38202 2759 38203 2815
rect 38145 2749 38203 2759
rect 38145 2735 38148 2749
rect 38200 2735 38203 2749
rect 38145 2679 38146 2735
rect 38202 2679 38203 2735
rect 38145 2655 38148 2679
rect 38200 2655 38203 2679
rect 38145 2599 38146 2655
rect 38202 2599 38203 2655
rect 38145 2575 38148 2599
rect 38200 2575 38203 2599
rect 38145 2519 38146 2575
rect 38202 2519 38203 2575
rect 38145 2505 38148 2519
rect 38200 2505 38203 2519
rect 38145 2495 38203 2505
rect 38145 2439 38146 2495
rect 38202 2439 38203 2495
rect 38145 2429 38203 2439
rect 38145 2415 38148 2429
rect 38200 2415 38203 2429
rect 38145 2359 38146 2415
rect 38202 2359 38203 2415
rect 38145 2335 38148 2359
rect 38200 2335 38203 2359
rect 38145 2279 38146 2335
rect 38202 2279 38203 2335
rect 38145 2255 38148 2279
rect 38200 2255 38203 2279
rect 38145 2199 38146 2255
rect 38202 2199 38203 2255
rect 38145 2185 38148 2199
rect 38200 2185 38203 2199
rect 38145 2175 38203 2185
rect 38145 2119 38146 2175
rect 38202 2119 38203 2175
rect 38145 2109 38203 2119
rect 38145 2095 38148 2109
rect 38200 2095 38203 2109
rect 38145 2039 38146 2095
rect 38202 2039 38203 2095
rect 38145 2015 38148 2039
rect 38200 2015 38203 2039
rect 38145 1959 38146 2015
rect 38202 1959 38203 2015
rect 38145 1935 38148 1959
rect 38200 1935 38203 1959
rect 38145 1879 38146 1935
rect 38202 1879 38203 1935
rect 38145 1865 38148 1879
rect 38200 1865 38203 1879
rect 38145 1855 38203 1865
rect 38145 1799 38146 1855
rect 38202 1799 38203 1855
rect 38145 1789 38203 1799
rect 38145 1775 38148 1789
rect 38200 1775 38203 1789
rect 38145 1719 38146 1775
rect 38202 1719 38203 1775
rect 38145 1695 38148 1719
rect 38200 1695 38203 1719
rect 38145 1639 38146 1695
rect 38202 1639 38203 1695
rect 38145 1615 38148 1639
rect 38200 1615 38203 1639
rect 38145 1559 38146 1615
rect 38202 1559 38203 1615
rect 38145 1545 38148 1559
rect 38200 1545 38203 1559
rect 38145 1535 38203 1545
rect 38145 1479 38146 1535
rect 38202 1479 38203 1535
rect 38145 1469 38203 1479
rect 38145 1455 38148 1469
rect 38200 1455 38203 1469
rect 38145 1399 38146 1455
rect 38202 1399 38203 1455
rect 38145 1375 38148 1399
rect 38200 1375 38203 1399
rect 38145 1319 38146 1375
rect 38202 1319 38203 1375
rect 38145 1295 38148 1319
rect 38200 1295 38203 1319
rect 38145 1239 38146 1295
rect 38202 1239 38203 1295
rect 38145 1225 38148 1239
rect 38200 1225 38203 1239
rect 38145 1215 38203 1225
rect 38145 1159 38146 1215
rect 38202 1159 38203 1215
rect 38145 1147 38203 1159
rect 38241 3133 38299 3147
rect 38241 3081 38244 3133
rect 38296 3081 38299 3133
rect 38241 3069 38299 3081
rect 38241 3017 38244 3069
rect 38296 3017 38299 3069
rect 38241 3005 38299 3017
rect 38241 2953 38244 3005
rect 38296 2953 38299 3005
rect 38241 2941 38299 2953
rect 38241 2889 38244 2941
rect 38296 2889 38299 2941
rect 38241 2877 38299 2889
rect 38241 2825 38244 2877
rect 38296 2825 38299 2877
rect 38241 2813 38299 2825
rect 38241 2761 38244 2813
rect 38296 2761 38299 2813
rect 38241 2749 38299 2761
rect 38241 2697 38244 2749
rect 38296 2697 38299 2749
rect 38241 2685 38299 2697
rect 38241 2633 38244 2685
rect 38296 2633 38299 2685
rect 38241 2621 38299 2633
rect 38241 2569 38244 2621
rect 38296 2569 38299 2621
rect 38241 2557 38299 2569
rect 38241 2505 38244 2557
rect 38296 2505 38299 2557
rect 38241 2493 38299 2505
rect 38241 2441 38244 2493
rect 38296 2441 38299 2493
rect 38241 2429 38299 2441
rect 38241 2377 38244 2429
rect 38296 2377 38299 2429
rect 38241 2365 38299 2377
rect 38241 2313 38244 2365
rect 38296 2313 38299 2365
rect 38241 2301 38299 2313
rect 38241 2249 38244 2301
rect 38296 2249 38299 2301
rect 38241 2237 38299 2249
rect 38241 2185 38244 2237
rect 38296 2185 38299 2237
rect 38241 2173 38299 2185
rect 38241 2121 38244 2173
rect 38296 2121 38299 2173
rect 38241 2109 38299 2121
rect 38241 2057 38244 2109
rect 38296 2057 38299 2109
rect 38241 2045 38299 2057
rect 38241 1993 38244 2045
rect 38296 1993 38299 2045
rect 38241 1981 38299 1993
rect 38241 1929 38244 1981
rect 38296 1929 38299 1981
rect 38241 1917 38299 1929
rect 38241 1865 38244 1917
rect 38296 1865 38299 1917
rect 38241 1853 38299 1865
rect 38241 1801 38244 1853
rect 38296 1801 38299 1853
rect 38241 1789 38299 1801
rect 38241 1737 38244 1789
rect 38296 1737 38299 1789
rect 38241 1725 38299 1737
rect 38241 1673 38244 1725
rect 38296 1673 38299 1725
rect 38241 1661 38299 1673
rect 38241 1609 38244 1661
rect 38296 1609 38299 1661
rect 38241 1597 38299 1609
rect 38241 1545 38244 1597
rect 38296 1545 38299 1597
rect 38241 1533 38299 1545
rect 38241 1481 38244 1533
rect 38296 1481 38299 1533
rect 38241 1469 38299 1481
rect 38241 1417 38244 1469
rect 38296 1417 38299 1469
rect 38241 1405 38299 1417
rect 38241 1353 38244 1405
rect 38296 1353 38299 1405
rect 38241 1341 38299 1353
rect 38241 1289 38244 1341
rect 38296 1289 38299 1341
rect 38241 1277 38299 1289
rect 38241 1225 38244 1277
rect 38296 1225 38299 1277
rect 38241 1213 38299 1225
rect 38241 1161 38244 1213
rect 38296 1161 38299 1213
rect 38241 830 38299 1161
rect 38337 3135 38395 3147
rect 38337 3079 38338 3135
rect 38394 3079 38395 3135
rect 38337 3069 38395 3079
rect 38337 3055 38340 3069
rect 38392 3055 38395 3069
rect 38337 2999 38338 3055
rect 38394 2999 38395 3055
rect 38337 2975 38340 2999
rect 38392 2975 38395 2999
rect 38337 2919 38338 2975
rect 38394 2919 38395 2975
rect 38337 2895 38340 2919
rect 38392 2895 38395 2919
rect 38337 2839 38338 2895
rect 38394 2839 38395 2895
rect 38337 2825 38340 2839
rect 38392 2825 38395 2839
rect 38337 2815 38395 2825
rect 38337 2759 38338 2815
rect 38394 2759 38395 2815
rect 38337 2749 38395 2759
rect 38337 2735 38340 2749
rect 38392 2735 38395 2749
rect 38337 2679 38338 2735
rect 38394 2679 38395 2735
rect 38337 2655 38340 2679
rect 38392 2655 38395 2679
rect 38337 2599 38338 2655
rect 38394 2599 38395 2655
rect 38337 2575 38340 2599
rect 38392 2575 38395 2599
rect 38337 2519 38338 2575
rect 38394 2519 38395 2575
rect 38337 2505 38340 2519
rect 38392 2505 38395 2519
rect 38337 2495 38395 2505
rect 38337 2439 38338 2495
rect 38394 2439 38395 2495
rect 38337 2429 38395 2439
rect 38337 2415 38340 2429
rect 38392 2415 38395 2429
rect 38337 2359 38338 2415
rect 38394 2359 38395 2415
rect 38337 2335 38340 2359
rect 38392 2335 38395 2359
rect 38337 2279 38338 2335
rect 38394 2279 38395 2335
rect 38337 2255 38340 2279
rect 38392 2255 38395 2279
rect 38337 2199 38338 2255
rect 38394 2199 38395 2255
rect 38337 2185 38340 2199
rect 38392 2185 38395 2199
rect 38337 2175 38395 2185
rect 38337 2119 38338 2175
rect 38394 2119 38395 2175
rect 38337 2109 38395 2119
rect 38337 2095 38340 2109
rect 38392 2095 38395 2109
rect 38337 2039 38338 2095
rect 38394 2039 38395 2095
rect 38337 2015 38340 2039
rect 38392 2015 38395 2039
rect 38337 1959 38338 2015
rect 38394 1959 38395 2015
rect 38337 1935 38340 1959
rect 38392 1935 38395 1959
rect 38337 1879 38338 1935
rect 38394 1879 38395 1935
rect 38337 1865 38340 1879
rect 38392 1865 38395 1879
rect 38337 1855 38395 1865
rect 38337 1799 38338 1855
rect 38394 1799 38395 1855
rect 38337 1789 38395 1799
rect 38337 1775 38340 1789
rect 38392 1775 38395 1789
rect 38337 1719 38338 1775
rect 38394 1719 38395 1775
rect 38337 1695 38340 1719
rect 38392 1695 38395 1719
rect 38337 1639 38338 1695
rect 38394 1639 38395 1695
rect 38337 1615 38340 1639
rect 38392 1615 38395 1639
rect 38337 1559 38338 1615
rect 38394 1559 38395 1615
rect 38337 1545 38340 1559
rect 38392 1545 38395 1559
rect 38337 1535 38395 1545
rect 38337 1479 38338 1535
rect 38394 1479 38395 1535
rect 38337 1469 38395 1479
rect 38337 1455 38340 1469
rect 38392 1455 38395 1469
rect 38337 1399 38338 1455
rect 38394 1399 38395 1455
rect 38337 1375 38340 1399
rect 38392 1375 38395 1399
rect 38337 1319 38338 1375
rect 38394 1319 38395 1375
rect 38337 1295 38340 1319
rect 38392 1295 38395 1319
rect 38337 1239 38338 1295
rect 38394 1239 38395 1295
rect 38337 1225 38340 1239
rect 38392 1225 38395 1239
rect 38337 1215 38395 1225
rect 38337 1159 38338 1215
rect 38394 1159 38395 1215
rect 38337 1147 38395 1159
rect 38433 3133 38491 3147
rect 38433 3081 38436 3133
rect 38488 3081 38491 3133
rect 38433 3069 38491 3081
rect 38433 3017 38436 3069
rect 38488 3017 38491 3069
rect 38433 3005 38491 3017
rect 38433 2953 38436 3005
rect 38488 2953 38491 3005
rect 38433 2941 38491 2953
rect 38433 2889 38436 2941
rect 38488 2889 38491 2941
rect 38433 2877 38491 2889
rect 38433 2825 38436 2877
rect 38488 2825 38491 2877
rect 38433 2813 38491 2825
rect 38433 2761 38436 2813
rect 38488 2761 38491 2813
rect 38433 2749 38491 2761
rect 38433 2697 38436 2749
rect 38488 2697 38491 2749
rect 38433 2685 38491 2697
rect 38433 2633 38436 2685
rect 38488 2633 38491 2685
rect 38433 2621 38491 2633
rect 38433 2569 38436 2621
rect 38488 2569 38491 2621
rect 38433 2557 38491 2569
rect 38433 2505 38436 2557
rect 38488 2505 38491 2557
rect 38433 2493 38491 2505
rect 38433 2441 38436 2493
rect 38488 2441 38491 2493
rect 38433 2429 38491 2441
rect 38433 2377 38436 2429
rect 38488 2377 38491 2429
rect 38433 2365 38491 2377
rect 38433 2313 38436 2365
rect 38488 2313 38491 2365
rect 38433 2301 38491 2313
rect 38433 2249 38436 2301
rect 38488 2249 38491 2301
rect 38433 2237 38491 2249
rect 38433 2185 38436 2237
rect 38488 2185 38491 2237
rect 38433 2173 38491 2185
rect 38433 2121 38436 2173
rect 38488 2121 38491 2173
rect 38433 2109 38491 2121
rect 38433 2057 38436 2109
rect 38488 2057 38491 2109
rect 38433 2045 38491 2057
rect 38433 1993 38436 2045
rect 38488 1993 38491 2045
rect 38433 1981 38491 1993
rect 38433 1929 38436 1981
rect 38488 1929 38491 1981
rect 38433 1917 38491 1929
rect 38433 1865 38436 1917
rect 38488 1865 38491 1917
rect 38433 1853 38491 1865
rect 38433 1801 38436 1853
rect 38488 1801 38491 1853
rect 38433 1789 38491 1801
rect 38433 1737 38436 1789
rect 38488 1737 38491 1789
rect 38433 1725 38491 1737
rect 38433 1673 38436 1725
rect 38488 1673 38491 1725
rect 38433 1661 38491 1673
rect 38433 1609 38436 1661
rect 38488 1609 38491 1661
rect 38433 1597 38491 1609
rect 38433 1545 38436 1597
rect 38488 1545 38491 1597
rect 38433 1533 38491 1545
rect 38433 1481 38436 1533
rect 38488 1481 38491 1533
rect 38433 1469 38491 1481
rect 38433 1417 38436 1469
rect 38488 1417 38491 1469
rect 38433 1405 38491 1417
rect 38433 1353 38436 1405
rect 38488 1353 38491 1405
rect 38433 1341 38491 1353
rect 38433 1289 38436 1341
rect 38488 1289 38491 1341
rect 38433 1277 38491 1289
rect 38433 1225 38436 1277
rect 38488 1225 38491 1277
rect 38433 1213 38491 1225
rect 38433 1161 38436 1213
rect 38488 1161 38491 1213
rect 38433 830 38491 1161
rect 38529 3135 38587 3147
rect 38529 3079 38530 3135
rect 38586 3079 38587 3135
rect 38529 3069 38587 3079
rect 38529 3055 38532 3069
rect 38584 3055 38587 3069
rect 38529 2999 38530 3055
rect 38586 2999 38587 3055
rect 38529 2975 38532 2999
rect 38584 2975 38587 2999
rect 38529 2919 38530 2975
rect 38586 2919 38587 2975
rect 38529 2895 38532 2919
rect 38584 2895 38587 2919
rect 38529 2839 38530 2895
rect 38586 2839 38587 2895
rect 38529 2825 38532 2839
rect 38584 2825 38587 2839
rect 38529 2815 38587 2825
rect 38529 2759 38530 2815
rect 38586 2759 38587 2815
rect 38529 2749 38587 2759
rect 38529 2735 38532 2749
rect 38584 2735 38587 2749
rect 38529 2679 38530 2735
rect 38586 2679 38587 2735
rect 38529 2655 38532 2679
rect 38584 2655 38587 2679
rect 38529 2599 38530 2655
rect 38586 2599 38587 2655
rect 38529 2575 38532 2599
rect 38584 2575 38587 2599
rect 38529 2519 38530 2575
rect 38586 2519 38587 2575
rect 38529 2505 38532 2519
rect 38584 2505 38587 2519
rect 38529 2495 38587 2505
rect 38529 2439 38530 2495
rect 38586 2439 38587 2495
rect 38529 2429 38587 2439
rect 38529 2415 38532 2429
rect 38584 2415 38587 2429
rect 38529 2359 38530 2415
rect 38586 2359 38587 2415
rect 38529 2335 38532 2359
rect 38584 2335 38587 2359
rect 38529 2279 38530 2335
rect 38586 2279 38587 2335
rect 38529 2255 38532 2279
rect 38584 2255 38587 2279
rect 38529 2199 38530 2255
rect 38586 2199 38587 2255
rect 38529 2185 38532 2199
rect 38584 2185 38587 2199
rect 38529 2175 38587 2185
rect 38529 2119 38530 2175
rect 38586 2119 38587 2175
rect 38529 2109 38587 2119
rect 38529 2095 38532 2109
rect 38584 2095 38587 2109
rect 38529 2039 38530 2095
rect 38586 2039 38587 2095
rect 38529 2015 38532 2039
rect 38584 2015 38587 2039
rect 38529 1959 38530 2015
rect 38586 1959 38587 2015
rect 38529 1935 38532 1959
rect 38584 1935 38587 1959
rect 38529 1879 38530 1935
rect 38586 1879 38587 1935
rect 38529 1865 38532 1879
rect 38584 1865 38587 1879
rect 38529 1855 38587 1865
rect 38529 1799 38530 1855
rect 38586 1799 38587 1855
rect 38529 1789 38587 1799
rect 38529 1775 38532 1789
rect 38584 1775 38587 1789
rect 38529 1719 38530 1775
rect 38586 1719 38587 1775
rect 38529 1695 38532 1719
rect 38584 1695 38587 1719
rect 38529 1639 38530 1695
rect 38586 1639 38587 1695
rect 38529 1615 38532 1639
rect 38584 1615 38587 1639
rect 38529 1559 38530 1615
rect 38586 1559 38587 1615
rect 38529 1545 38532 1559
rect 38584 1545 38587 1559
rect 38529 1535 38587 1545
rect 38529 1479 38530 1535
rect 38586 1479 38587 1535
rect 38529 1469 38587 1479
rect 38529 1455 38532 1469
rect 38584 1455 38587 1469
rect 38529 1399 38530 1455
rect 38586 1399 38587 1455
rect 38529 1375 38532 1399
rect 38584 1375 38587 1399
rect 38529 1319 38530 1375
rect 38586 1319 38587 1375
rect 38529 1295 38532 1319
rect 38584 1295 38587 1319
rect 38529 1239 38530 1295
rect 38586 1239 38587 1295
rect 38529 1225 38532 1239
rect 38584 1225 38587 1239
rect 38529 1215 38587 1225
rect 38529 1159 38530 1215
rect 38586 1159 38587 1215
rect 38529 1147 38587 1159
rect 38625 3132 38683 3146
rect 38625 3080 38628 3132
rect 38680 3080 38683 3132
rect 38625 3068 38683 3080
rect 38625 3016 38628 3068
rect 38680 3016 38683 3068
rect 38625 3004 38683 3016
rect 38625 2952 38628 3004
rect 38680 2952 38683 3004
rect 38625 2940 38683 2952
rect 38625 2888 38628 2940
rect 38680 2888 38683 2940
rect 38625 2876 38683 2888
rect 38625 2824 38628 2876
rect 38680 2824 38683 2876
rect 38625 2812 38683 2824
rect 38625 2760 38628 2812
rect 38680 2760 38683 2812
rect 38625 2748 38683 2760
rect 38625 2696 38628 2748
rect 38680 2696 38683 2748
rect 38625 2684 38683 2696
rect 38625 2632 38628 2684
rect 38680 2632 38683 2684
rect 38625 2620 38683 2632
rect 38625 2568 38628 2620
rect 38680 2568 38683 2620
rect 38625 2556 38683 2568
rect 38625 2504 38628 2556
rect 38680 2504 38683 2556
rect 38625 2492 38683 2504
rect 38625 2440 38628 2492
rect 38680 2440 38683 2492
rect 38625 2428 38683 2440
rect 38625 2376 38628 2428
rect 38680 2376 38683 2428
rect 38625 2364 38683 2376
rect 38625 2312 38628 2364
rect 38680 2312 38683 2364
rect 38625 2300 38683 2312
rect 38625 2248 38628 2300
rect 38680 2248 38683 2300
rect 38625 2236 38683 2248
rect 38625 2184 38628 2236
rect 38680 2184 38683 2236
rect 38625 2172 38683 2184
rect 38625 2120 38628 2172
rect 38680 2120 38683 2172
rect 38625 2108 38683 2120
rect 38625 2056 38628 2108
rect 38680 2056 38683 2108
rect 38625 2044 38683 2056
rect 38625 1992 38628 2044
rect 38680 1992 38683 2044
rect 38625 1980 38683 1992
rect 38625 1928 38628 1980
rect 38680 1928 38683 1980
rect 38625 1916 38683 1928
rect 38625 1864 38628 1916
rect 38680 1864 38683 1916
rect 38625 1852 38683 1864
rect 38625 1800 38628 1852
rect 38680 1800 38683 1852
rect 38625 1788 38683 1800
rect 38625 1736 38628 1788
rect 38680 1736 38683 1788
rect 38625 1724 38683 1736
rect 38625 1672 38628 1724
rect 38680 1672 38683 1724
rect 38625 1660 38683 1672
rect 38625 1608 38628 1660
rect 38680 1608 38683 1660
rect 38625 1596 38683 1608
rect 38625 1544 38628 1596
rect 38680 1544 38683 1596
rect 38625 1532 38683 1544
rect 38625 1480 38628 1532
rect 38680 1480 38683 1532
rect 38625 1468 38683 1480
rect 38625 1416 38628 1468
rect 38680 1416 38683 1468
rect 38625 1404 38683 1416
rect 38625 1352 38628 1404
rect 38680 1352 38683 1404
rect 38625 1340 38683 1352
rect 38625 1288 38628 1340
rect 38680 1288 38683 1340
rect 38625 1276 38683 1288
rect 38625 1224 38628 1276
rect 38680 1224 38683 1276
rect 38625 1212 38683 1224
rect 38625 1160 38628 1212
rect 38680 1160 38683 1212
rect 38625 830 38683 1160
rect 29025 746 38684 830
rect 38625 745 38683 746
<< via2 >>
rect 29122 3133 29178 3135
rect 29122 3081 29124 3133
rect 29124 3081 29176 3133
rect 29176 3081 29178 3133
rect 29122 3079 29178 3081
rect 29122 3017 29124 3055
rect 29124 3017 29176 3055
rect 29176 3017 29178 3055
rect 29122 3005 29178 3017
rect 29122 2999 29124 3005
rect 29124 2999 29176 3005
rect 29176 2999 29178 3005
rect 29122 2953 29124 2975
rect 29124 2953 29176 2975
rect 29176 2953 29178 2975
rect 29122 2941 29178 2953
rect 29122 2919 29124 2941
rect 29124 2919 29176 2941
rect 29176 2919 29178 2941
rect 29122 2889 29124 2895
rect 29124 2889 29176 2895
rect 29176 2889 29178 2895
rect 29122 2877 29178 2889
rect 29122 2839 29124 2877
rect 29124 2839 29176 2877
rect 29176 2839 29178 2877
rect 29122 2813 29178 2815
rect 29122 2761 29124 2813
rect 29124 2761 29176 2813
rect 29176 2761 29178 2813
rect 29122 2759 29178 2761
rect 29122 2697 29124 2735
rect 29124 2697 29176 2735
rect 29176 2697 29178 2735
rect 29122 2685 29178 2697
rect 29122 2679 29124 2685
rect 29124 2679 29176 2685
rect 29176 2679 29178 2685
rect 29122 2633 29124 2655
rect 29124 2633 29176 2655
rect 29176 2633 29178 2655
rect 29122 2621 29178 2633
rect 29122 2599 29124 2621
rect 29124 2599 29176 2621
rect 29176 2599 29178 2621
rect 29122 2569 29124 2575
rect 29124 2569 29176 2575
rect 29176 2569 29178 2575
rect 29122 2557 29178 2569
rect 29122 2519 29124 2557
rect 29124 2519 29176 2557
rect 29176 2519 29178 2557
rect 29122 2493 29178 2495
rect 29122 2441 29124 2493
rect 29124 2441 29176 2493
rect 29176 2441 29178 2493
rect 29122 2439 29178 2441
rect 29122 2377 29124 2415
rect 29124 2377 29176 2415
rect 29176 2377 29178 2415
rect 29122 2365 29178 2377
rect 29122 2359 29124 2365
rect 29124 2359 29176 2365
rect 29176 2359 29178 2365
rect 29122 2313 29124 2335
rect 29124 2313 29176 2335
rect 29176 2313 29178 2335
rect 29122 2301 29178 2313
rect 29122 2279 29124 2301
rect 29124 2279 29176 2301
rect 29176 2279 29178 2301
rect 29122 2249 29124 2255
rect 29124 2249 29176 2255
rect 29176 2249 29178 2255
rect 29122 2237 29178 2249
rect 29122 2199 29124 2237
rect 29124 2199 29176 2237
rect 29176 2199 29178 2237
rect 29122 2173 29178 2175
rect 29122 2121 29124 2173
rect 29124 2121 29176 2173
rect 29176 2121 29178 2173
rect 29122 2119 29178 2121
rect 29122 2057 29124 2095
rect 29124 2057 29176 2095
rect 29176 2057 29178 2095
rect 29122 2045 29178 2057
rect 29122 2039 29124 2045
rect 29124 2039 29176 2045
rect 29176 2039 29178 2045
rect 29122 1993 29124 2015
rect 29124 1993 29176 2015
rect 29176 1993 29178 2015
rect 29122 1981 29178 1993
rect 29122 1959 29124 1981
rect 29124 1959 29176 1981
rect 29176 1959 29178 1981
rect 29122 1929 29124 1935
rect 29124 1929 29176 1935
rect 29176 1929 29178 1935
rect 29122 1917 29178 1929
rect 29122 1879 29124 1917
rect 29124 1879 29176 1917
rect 29176 1879 29178 1917
rect 29122 1853 29178 1855
rect 29122 1801 29124 1853
rect 29124 1801 29176 1853
rect 29176 1801 29178 1853
rect 29122 1799 29178 1801
rect 29122 1737 29124 1775
rect 29124 1737 29176 1775
rect 29176 1737 29178 1775
rect 29122 1725 29178 1737
rect 29122 1719 29124 1725
rect 29124 1719 29176 1725
rect 29176 1719 29178 1725
rect 29122 1673 29124 1695
rect 29124 1673 29176 1695
rect 29176 1673 29178 1695
rect 29122 1661 29178 1673
rect 29122 1639 29124 1661
rect 29124 1639 29176 1661
rect 29176 1639 29178 1661
rect 29122 1609 29124 1615
rect 29124 1609 29176 1615
rect 29176 1609 29178 1615
rect 29122 1597 29178 1609
rect 29122 1559 29124 1597
rect 29124 1559 29176 1597
rect 29176 1559 29178 1597
rect 29122 1533 29178 1535
rect 29122 1481 29124 1533
rect 29124 1481 29176 1533
rect 29176 1481 29178 1533
rect 29122 1479 29178 1481
rect 29122 1417 29124 1455
rect 29124 1417 29176 1455
rect 29176 1417 29178 1455
rect 29122 1405 29178 1417
rect 29122 1399 29124 1405
rect 29124 1399 29176 1405
rect 29176 1399 29178 1405
rect 29122 1353 29124 1375
rect 29124 1353 29176 1375
rect 29176 1353 29178 1375
rect 29122 1341 29178 1353
rect 29122 1319 29124 1341
rect 29124 1319 29176 1341
rect 29176 1319 29178 1341
rect 29122 1289 29124 1295
rect 29124 1289 29176 1295
rect 29176 1289 29178 1295
rect 29122 1277 29178 1289
rect 29122 1239 29124 1277
rect 29124 1239 29176 1277
rect 29176 1239 29178 1277
rect 29122 1213 29178 1215
rect 29122 1161 29124 1213
rect 29124 1161 29176 1213
rect 29176 1161 29178 1213
rect 29122 1159 29178 1161
rect 29314 3133 29370 3135
rect 29314 3081 29316 3133
rect 29316 3081 29368 3133
rect 29368 3081 29370 3133
rect 29314 3079 29370 3081
rect 29314 3017 29316 3055
rect 29316 3017 29368 3055
rect 29368 3017 29370 3055
rect 29314 3005 29370 3017
rect 29314 2999 29316 3005
rect 29316 2999 29368 3005
rect 29368 2999 29370 3005
rect 29314 2953 29316 2975
rect 29316 2953 29368 2975
rect 29368 2953 29370 2975
rect 29314 2941 29370 2953
rect 29314 2919 29316 2941
rect 29316 2919 29368 2941
rect 29368 2919 29370 2941
rect 29314 2889 29316 2895
rect 29316 2889 29368 2895
rect 29368 2889 29370 2895
rect 29314 2877 29370 2889
rect 29314 2839 29316 2877
rect 29316 2839 29368 2877
rect 29368 2839 29370 2877
rect 29314 2813 29370 2815
rect 29314 2761 29316 2813
rect 29316 2761 29368 2813
rect 29368 2761 29370 2813
rect 29314 2759 29370 2761
rect 29314 2697 29316 2735
rect 29316 2697 29368 2735
rect 29368 2697 29370 2735
rect 29314 2685 29370 2697
rect 29314 2679 29316 2685
rect 29316 2679 29368 2685
rect 29368 2679 29370 2685
rect 29314 2633 29316 2655
rect 29316 2633 29368 2655
rect 29368 2633 29370 2655
rect 29314 2621 29370 2633
rect 29314 2599 29316 2621
rect 29316 2599 29368 2621
rect 29368 2599 29370 2621
rect 29314 2569 29316 2575
rect 29316 2569 29368 2575
rect 29368 2569 29370 2575
rect 29314 2557 29370 2569
rect 29314 2519 29316 2557
rect 29316 2519 29368 2557
rect 29368 2519 29370 2557
rect 29314 2493 29370 2495
rect 29314 2441 29316 2493
rect 29316 2441 29368 2493
rect 29368 2441 29370 2493
rect 29314 2439 29370 2441
rect 29314 2377 29316 2415
rect 29316 2377 29368 2415
rect 29368 2377 29370 2415
rect 29314 2365 29370 2377
rect 29314 2359 29316 2365
rect 29316 2359 29368 2365
rect 29368 2359 29370 2365
rect 29314 2313 29316 2335
rect 29316 2313 29368 2335
rect 29368 2313 29370 2335
rect 29314 2301 29370 2313
rect 29314 2279 29316 2301
rect 29316 2279 29368 2301
rect 29368 2279 29370 2301
rect 29314 2249 29316 2255
rect 29316 2249 29368 2255
rect 29368 2249 29370 2255
rect 29314 2237 29370 2249
rect 29314 2199 29316 2237
rect 29316 2199 29368 2237
rect 29368 2199 29370 2237
rect 29314 2173 29370 2175
rect 29314 2121 29316 2173
rect 29316 2121 29368 2173
rect 29368 2121 29370 2173
rect 29314 2119 29370 2121
rect 29314 2057 29316 2095
rect 29316 2057 29368 2095
rect 29368 2057 29370 2095
rect 29314 2045 29370 2057
rect 29314 2039 29316 2045
rect 29316 2039 29368 2045
rect 29368 2039 29370 2045
rect 29314 1993 29316 2015
rect 29316 1993 29368 2015
rect 29368 1993 29370 2015
rect 29314 1981 29370 1993
rect 29314 1959 29316 1981
rect 29316 1959 29368 1981
rect 29368 1959 29370 1981
rect 29314 1929 29316 1935
rect 29316 1929 29368 1935
rect 29368 1929 29370 1935
rect 29314 1917 29370 1929
rect 29314 1879 29316 1917
rect 29316 1879 29368 1917
rect 29368 1879 29370 1917
rect 29314 1853 29370 1855
rect 29314 1801 29316 1853
rect 29316 1801 29368 1853
rect 29368 1801 29370 1853
rect 29314 1799 29370 1801
rect 29314 1737 29316 1775
rect 29316 1737 29368 1775
rect 29368 1737 29370 1775
rect 29314 1725 29370 1737
rect 29314 1719 29316 1725
rect 29316 1719 29368 1725
rect 29368 1719 29370 1725
rect 29314 1673 29316 1695
rect 29316 1673 29368 1695
rect 29368 1673 29370 1695
rect 29314 1661 29370 1673
rect 29314 1639 29316 1661
rect 29316 1639 29368 1661
rect 29368 1639 29370 1661
rect 29314 1609 29316 1615
rect 29316 1609 29368 1615
rect 29368 1609 29370 1615
rect 29314 1597 29370 1609
rect 29314 1559 29316 1597
rect 29316 1559 29368 1597
rect 29368 1559 29370 1597
rect 29314 1533 29370 1535
rect 29314 1481 29316 1533
rect 29316 1481 29368 1533
rect 29368 1481 29370 1533
rect 29314 1479 29370 1481
rect 29314 1417 29316 1455
rect 29316 1417 29368 1455
rect 29368 1417 29370 1455
rect 29314 1405 29370 1417
rect 29314 1399 29316 1405
rect 29316 1399 29368 1405
rect 29368 1399 29370 1405
rect 29314 1353 29316 1375
rect 29316 1353 29368 1375
rect 29368 1353 29370 1375
rect 29314 1341 29370 1353
rect 29314 1319 29316 1341
rect 29316 1319 29368 1341
rect 29368 1319 29370 1341
rect 29314 1289 29316 1295
rect 29316 1289 29368 1295
rect 29368 1289 29370 1295
rect 29314 1277 29370 1289
rect 29314 1239 29316 1277
rect 29316 1239 29368 1277
rect 29368 1239 29370 1277
rect 29314 1213 29370 1215
rect 29314 1161 29316 1213
rect 29316 1161 29368 1213
rect 29368 1161 29370 1213
rect 29314 1159 29370 1161
rect 29506 3133 29562 3135
rect 29506 3081 29508 3133
rect 29508 3081 29560 3133
rect 29560 3081 29562 3133
rect 29506 3079 29562 3081
rect 29506 3017 29508 3055
rect 29508 3017 29560 3055
rect 29560 3017 29562 3055
rect 29506 3005 29562 3017
rect 29506 2999 29508 3005
rect 29508 2999 29560 3005
rect 29560 2999 29562 3005
rect 29506 2953 29508 2975
rect 29508 2953 29560 2975
rect 29560 2953 29562 2975
rect 29506 2941 29562 2953
rect 29506 2919 29508 2941
rect 29508 2919 29560 2941
rect 29560 2919 29562 2941
rect 29506 2889 29508 2895
rect 29508 2889 29560 2895
rect 29560 2889 29562 2895
rect 29506 2877 29562 2889
rect 29506 2839 29508 2877
rect 29508 2839 29560 2877
rect 29560 2839 29562 2877
rect 29506 2813 29562 2815
rect 29506 2761 29508 2813
rect 29508 2761 29560 2813
rect 29560 2761 29562 2813
rect 29506 2759 29562 2761
rect 29506 2697 29508 2735
rect 29508 2697 29560 2735
rect 29560 2697 29562 2735
rect 29506 2685 29562 2697
rect 29506 2679 29508 2685
rect 29508 2679 29560 2685
rect 29560 2679 29562 2685
rect 29506 2633 29508 2655
rect 29508 2633 29560 2655
rect 29560 2633 29562 2655
rect 29506 2621 29562 2633
rect 29506 2599 29508 2621
rect 29508 2599 29560 2621
rect 29560 2599 29562 2621
rect 29506 2569 29508 2575
rect 29508 2569 29560 2575
rect 29560 2569 29562 2575
rect 29506 2557 29562 2569
rect 29506 2519 29508 2557
rect 29508 2519 29560 2557
rect 29560 2519 29562 2557
rect 29506 2493 29562 2495
rect 29506 2441 29508 2493
rect 29508 2441 29560 2493
rect 29560 2441 29562 2493
rect 29506 2439 29562 2441
rect 29506 2377 29508 2415
rect 29508 2377 29560 2415
rect 29560 2377 29562 2415
rect 29506 2365 29562 2377
rect 29506 2359 29508 2365
rect 29508 2359 29560 2365
rect 29560 2359 29562 2365
rect 29506 2313 29508 2335
rect 29508 2313 29560 2335
rect 29560 2313 29562 2335
rect 29506 2301 29562 2313
rect 29506 2279 29508 2301
rect 29508 2279 29560 2301
rect 29560 2279 29562 2301
rect 29506 2249 29508 2255
rect 29508 2249 29560 2255
rect 29560 2249 29562 2255
rect 29506 2237 29562 2249
rect 29506 2199 29508 2237
rect 29508 2199 29560 2237
rect 29560 2199 29562 2237
rect 29506 2173 29562 2175
rect 29506 2121 29508 2173
rect 29508 2121 29560 2173
rect 29560 2121 29562 2173
rect 29506 2119 29562 2121
rect 29506 2057 29508 2095
rect 29508 2057 29560 2095
rect 29560 2057 29562 2095
rect 29506 2045 29562 2057
rect 29506 2039 29508 2045
rect 29508 2039 29560 2045
rect 29560 2039 29562 2045
rect 29506 1993 29508 2015
rect 29508 1993 29560 2015
rect 29560 1993 29562 2015
rect 29506 1981 29562 1993
rect 29506 1959 29508 1981
rect 29508 1959 29560 1981
rect 29560 1959 29562 1981
rect 29506 1929 29508 1935
rect 29508 1929 29560 1935
rect 29560 1929 29562 1935
rect 29506 1917 29562 1929
rect 29506 1879 29508 1917
rect 29508 1879 29560 1917
rect 29560 1879 29562 1917
rect 29506 1853 29562 1855
rect 29506 1801 29508 1853
rect 29508 1801 29560 1853
rect 29560 1801 29562 1853
rect 29506 1799 29562 1801
rect 29506 1737 29508 1775
rect 29508 1737 29560 1775
rect 29560 1737 29562 1775
rect 29506 1725 29562 1737
rect 29506 1719 29508 1725
rect 29508 1719 29560 1725
rect 29560 1719 29562 1725
rect 29506 1673 29508 1695
rect 29508 1673 29560 1695
rect 29560 1673 29562 1695
rect 29506 1661 29562 1673
rect 29506 1639 29508 1661
rect 29508 1639 29560 1661
rect 29560 1639 29562 1661
rect 29506 1609 29508 1615
rect 29508 1609 29560 1615
rect 29560 1609 29562 1615
rect 29506 1597 29562 1609
rect 29506 1559 29508 1597
rect 29508 1559 29560 1597
rect 29560 1559 29562 1597
rect 29506 1533 29562 1535
rect 29506 1481 29508 1533
rect 29508 1481 29560 1533
rect 29560 1481 29562 1533
rect 29506 1479 29562 1481
rect 29506 1417 29508 1455
rect 29508 1417 29560 1455
rect 29560 1417 29562 1455
rect 29506 1405 29562 1417
rect 29506 1399 29508 1405
rect 29508 1399 29560 1405
rect 29560 1399 29562 1405
rect 29506 1353 29508 1375
rect 29508 1353 29560 1375
rect 29560 1353 29562 1375
rect 29506 1341 29562 1353
rect 29506 1319 29508 1341
rect 29508 1319 29560 1341
rect 29560 1319 29562 1341
rect 29506 1289 29508 1295
rect 29508 1289 29560 1295
rect 29560 1289 29562 1295
rect 29506 1277 29562 1289
rect 29506 1239 29508 1277
rect 29508 1239 29560 1277
rect 29560 1239 29562 1277
rect 29506 1213 29562 1215
rect 29506 1161 29508 1213
rect 29508 1161 29560 1213
rect 29560 1161 29562 1213
rect 29506 1159 29562 1161
rect 29698 3133 29754 3135
rect 29698 3081 29700 3133
rect 29700 3081 29752 3133
rect 29752 3081 29754 3133
rect 29698 3079 29754 3081
rect 29698 3017 29700 3055
rect 29700 3017 29752 3055
rect 29752 3017 29754 3055
rect 29698 3005 29754 3017
rect 29698 2999 29700 3005
rect 29700 2999 29752 3005
rect 29752 2999 29754 3005
rect 29698 2953 29700 2975
rect 29700 2953 29752 2975
rect 29752 2953 29754 2975
rect 29698 2941 29754 2953
rect 29698 2919 29700 2941
rect 29700 2919 29752 2941
rect 29752 2919 29754 2941
rect 29698 2889 29700 2895
rect 29700 2889 29752 2895
rect 29752 2889 29754 2895
rect 29698 2877 29754 2889
rect 29698 2839 29700 2877
rect 29700 2839 29752 2877
rect 29752 2839 29754 2877
rect 29698 2813 29754 2815
rect 29698 2761 29700 2813
rect 29700 2761 29752 2813
rect 29752 2761 29754 2813
rect 29698 2759 29754 2761
rect 29698 2697 29700 2735
rect 29700 2697 29752 2735
rect 29752 2697 29754 2735
rect 29698 2685 29754 2697
rect 29698 2679 29700 2685
rect 29700 2679 29752 2685
rect 29752 2679 29754 2685
rect 29698 2633 29700 2655
rect 29700 2633 29752 2655
rect 29752 2633 29754 2655
rect 29698 2621 29754 2633
rect 29698 2599 29700 2621
rect 29700 2599 29752 2621
rect 29752 2599 29754 2621
rect 29698 2569 29700 2575
rect 29700 2569 29752 2575
rect 29752 2569 29754 2575
rect 29698 2557 29754 2569
rect 29698 2519 29700 2557
rect 29700 2519 29752 2557
rect 29752 2519 29754 2557
rect 29698 2493 29754 2495
rect 29698 2441 29700 2493
rect 29700 2441 29752 2493
rect 29752 2441 29754 2493
rect 29698 2439 29754 2441
rect 29698 2377 29700 2415
rect 29700 2377 29752 2415
rect 29752 2377 29754 2415
rect 29698 2365 29754 2377
rect 29698 2359 29700 2365
rect 29700 2359 29752 2365
rect 29752 2359 29754 2365
rect 29698 2313 29700 2335
rect 29700 2313 29752 2335
rect 29752 2313 29754 2335
rect 29698 2301 29754 2313
rect 29698 2279 29700 2301
rect 29700 2279 29752 2301
rect 29752 2279 29754 2301
rect 29698 2249 29700 2255
rect 29700 2249 29752 2255
rect 29752 2249 29754 2255
rect 29698 2237 29754 2249
rect 29698 2199 29700 2237
rect 29700 2199 29752 2237
rect 29752 2199 29754 2237
rect 29698 2173 29754 2175
rect 29698 2121 29700 2173
rect 29700 2121 29752 2173
rect 29752 2121 29754 2173
rect 29698 2119 29754 2121
rect 29698 2057 29700 2095
rect 29700 2057 29752 2095
rect 29752 2057 29754 2095
rect 29698 2045 29754 2057
rect 29698 2039 29700 2045
rect 29700 2039 29752 2045
rect 29752 2039 29754 2045
rect 29698 1993 29700 2015
rect 29700 1993 29752 2015
rect 29752 1993 29754 2015
rect 29698 1981 29754 1993
rect 29698 1959 29700 1981
rect 29700 1959 29752 1981
rect 29752 1959 29754 1981
rect 29698 1929 29700 1935
rect 29700 1929 29752 1935
rect 29752 1929 29754 1935
rect 29698 1917 29754 1929
rect 29698 1879 29700 1917
rect 29700 1879 29752 1917
rect 29752 1879 29754 1917
rect 29698 1853 29754 1855
rect 29698 1801 29700 1853
rect 29700 1801 29752 1853
rect 29752 1801 29754 1853
rect 29698 1799 29754 1801
rect 29698 1737 29700 1775
rect 29700 1737 29752 1775
rect 29752 1737 29754 1775
rect 29698 1725 29754 1737
rect 29698 1719 29700 1725
rect 29700 1719 29752 1725
rect 29752 1719 29754 1725
rect 29698 1673 29700 1695
rect 29700 1673 29752 1695
rect 29752 1673 29754 1695
rect 29698 1661 29754 1673
rect 29698 1639 29700 1661
rect 29700 1639 29752 1661
rect 29752 1639 29754 1661
rect 29698 1609 29700 1615
rect 29700 1609 29752 1615
rect 29752 1609 29754 1615
rect 29698 1597 29754 1609
rect 29698 1559 29700 1597
rect 29700 1559 29752 1597
rect 29752 1559 29754 1597
rect 29698 1533 29754 1535
rect 29698 1481 29700 1533
rect 29700 1481 29752 1533
rect 29752 1481 29754 1533
rect 29698 1479 29754 1481
rect 29698 1417 29700 1455
rect 29700 1417 29752 1455
rect 29752 1417 29754 1455
rect 29698 1405 29754 1417
rect 29698 1399 29700 1405
rect 29700 1399 29752 1405
rect 29752 1399 29754 1405
rect 29698 1353 29700 1375
rect 29700 1353 29752 1375
rect 29752 1353 29754 1375
rect 29698 1341 29754 1353
rect 29698 1319 29700 1341
rect 29700 1319 29752 1341
rect 29752 1319 29754 1341
rect 29698 1289 29700 1295
rect 29700 1289 29752 1295
rect 29752 1289 29754 1295
rect 29698 1277 29754 1289
rect 29698 1239 29700 1277
rect 29700 1239 29752 1277
rect 29752 1239 29754 1277
rect 29698 1213 29754 1215
rect 29698 1161 29700 1213
rect 29700 1161 29752 1213
rect 29752 1161 29754 1213
rect 29698 1159 29754 1161
rect 29890 3133 29946 3135
rect 29890 3081 29892 3133
rect 29892 3081 29944 3133
rect 29944 3081 29946 3133
rect 29890 3079 29946 3081
rect 29890 3017 29892 3055
rect 29892 3017 29944 3055
rect 29944 3017 29946 3055
rect 29890 3005 29946 3017
rect 29890 2999 29892 3005
rect 29892 2999 29944 3005
rect 29944 2999 29946 3005
rect 29890 2953 29892 2975
rect 29892 2953 29944 2975
rect 29944 2953 29946 2975
rect 29890 2941 29946 2953
rect 29890 2919 29892 2941
rect 29892 2919 29944 2941
rect 29944 2919 29946 2941
rect 29890 2889 29892 2895
rect 29892 2889 29944 2895
rect 29944 2889 29946 2895
rect 29890 2877 29946 2889
rect 29890 2839 29892 2877
rect 29892 2839 29944 2877
rect 29944 2839 29946 2877
rect 29890 2813 29946 2815
rect 29890 2761 29892 2813
rect 29892 2761 29944 2813
rect 29944 2761 29946 2813
rect 29890 2759 29946 2761
rect 29890 2697 29892 2735
rect 29892 2697 29944 2735
rect 29944 2697 29946 2735
rect 29890 2685 29946 2697
rect 29890 2679 29892 2685
rect 29892 2679 29944 2685
rect 29944 2679 29946 2685
rect 29890 2633 29892 2655
rect 29892 2633 29944 2655
rect 29944 2633 29946 2655
rect 29890 2621 29946 2633
rect 29890 2599 29892 2621
rect 29892 2599 29944 2621
rect 29944 2599 29946 2621
rect 29890 2569 29892 2575
rect 29892 2569 29944 2575
rect 29944 2569 29946 2575
rect 29890 2557 29946 2569
rect 29890 2519 29892 2557
rect 29892 2519 29944 2557
rect 29944 2519 29946 2557
rect 29890 2493 29946 2495
rect 29890 2441 29892 2493
rect 29892 2441 29944 2493
rect 29944 2441 29946 2493
rect 29890 2439 29946 2441
rect 29890 2377 29892 2415
rect 29892 2377 29944 2415
rect 29944 2377 29946 2415
rect 29890 2365 29946 2377
rect 29890 2359 29892 2365
rect 29892 2359 29944 2365
rect 29944 2359 29946 2365
rect 29890 2313 29892 2335
rect 29892 2313 29944 2335
rect 29944 2313 29946 2335
rect 29890 2301 29946 2313
rect 29890 2279 29892 2301
rect 29892 2279 29944 2301
rect 29944 2279 29946 2301
rect 29890 2249 29892 2255
rect 29892 2249 29944 2255
rect 29944 2249 29946 2255
rect 29890 2237 29946 2249
rect 29890 2199 29892 2237
rect 29892 2199 29944 2237
rect 29944 2199 29946 2237
rect 29890 2173 29946 2175
rect 29890 2121 29892 2173
rect 29892 2121 29944 2173
rect 29944 2121 29946 2173
rect 29890 2119 29946 2121
rect 29890 2057 29892 2095
rect 29892 2057 29944 2095
rect 29944 2057 29946 2095
rect 29890 2045 29946 2057
rect 29890 2039 29892 2045
rect 29892 2039 29944 2045
rect 29944 2039 29946 2045
rect 29890 1993 29892 2015
rect 29892 1993 29944 2015
rect 29944 1993 29946 2015
rect 29890 1981 29946 1993
rect 29890 1959 29892 1981
rect 29892 1959 29944 1981
rect 29944 1959 29946 1981
rect 29890 1929 29892 1935
rect 29892 1929 29944 1935
rect 29944 1929 29946 1935
rect 29890 1917 29946 1929
rect 29890 1879 29892 1917
rect 29892 1879 29944 1917
rect 29944 1879 29946 1917
rect 29890 1853 29946 1855
rect 29890 1801 29892 1853
rect 29892 1801 29944 1853
rect 29944 1801 29946 1853
rect 29890 1799 29946 1801
rect 29890 1737 29892 1775
rect 29892 1737 29944 1775
rect 29944 1737 29946 1775
rect 29890 1725 29946 1737
rect 29890 1719 29892 1725
rect 29892 1719 29944 1725
rect 29944 1719 29946 1725
rect 29890 1673 29892 1695
rect 29892 1673 29944 1695
rect 29944 1673 29946 1695
rect 29890 1661 29946 1673
rect 29890 1639 29892 1661
rect 29892 1639 29944 1661
rect 29944 1639 29946 1661
rect 29890 1609 29892 1615
rect 29892 1609 29944 1615
rect 29944 1609 29946 1615
rect 29890 1597 29946 1609
rect 29890 1559 29892 1597
rect 29892 1559 29944 1597
rect 29944 1559 29946 1597
rect 29890 1533 29946 1535
rect 29890 1481 29892 1533
rect 29892 1481 29944 1533
rect 29944 1481 29946 1533
rect 29890 1479 29946 1481
rect 29890 1417 29892 1455
rect 29892 1417 29944 1455
rect 29944 1417 29946 1455
rect 29890 1405 29946 1417
rect 29890 1399 29892 1405
rect 29892 1399 29944 1405
rect 29944 1399 29946 1405
rect 29890 1353 29892 1375
rect 29892 1353 29944 1375
rect 29944 1353 29946 1375
rect 29890 1341 29946 1353
rect 29890 1319 29892 1341
rect 29892 1319 29944 1341
rect 29944 1319 29946 1341
rect 29890 1289 29892 1295
rect 29892 1289 29944 1295
rect 29944 1289 29946 1295
rect 29890 1277 29946 1289
rect 29890 1239 29892 1277
rect 29892 1239 29944 1277
rect 29944 1239 29946 1277
rect 29890 1213 29946 1215
rect 29890 1161 29892 1213
rect 29892 1161 29944 1213
rect 29944 1161 29946 1213
rect 29890 1159 29946 1161
rect 30082 3133 30138 3135
rect 30082 3081 30084 3133
rect 30084 3081 30136 3133
rect 30136 3081 30138 3133
rect 30082 3079 30138 3081
rect 30082 3017 30084 3055
rect 30084 3017 30136 3055
rect 30136 3017 30138 3055
rect 30082 3005 30138 3017
rect 30082 2999 30084 3005
rect 30084 2999 30136 3005
rect 30136 2999 30138 3005
rect 30082 2953 30084 2975
rect 30084 2953 30136 2975
rect 30136 2953 30138 2975
rect 30082 2941 30138 2953
rect 30082 2919 30084 2941
rect 30084 2919 30136 2941
rect 30136 2919 30138 2941
rect 30082 2889 30084 2895
rect 30084 2889 30136 2895
rect 30136 2889 30138 2895
rect 30082 2877 30138 2889
rect 30082 2839 30084 2877
rect 30084 2839 30136 2877
rect 30136 2839 30138 2877
rect 30082 2813 30138 2815
rect 30082 2761 30084 2813
rect 30084 2761 30136 2813
rect 30136 2761 30138 2813
rect 30082 2759 30138 2761
rect 30082 2697 30084 2735
rect 30084 2697 30136 2735
rect 30136 2697 30138 2735
rect 30082 2685 30138 2697
rect 30082 2679 30084 2685
rect 30084 2679 30136 2685
rect 30136 2679 30138 2685
rect 30082 2633 30084 2655
rect 30084 2633 30136 2655
rect 30136 2633 30138 2655
rect 30082 2621 30138 2633
rect 30082 2599 30084 2621
rect 30084 2599 30136 2621
rect 30136 2599 30138 2621
rect 30082 2569 30084 2575
rect 30084 2569 30136 2575
rect 30136 2569 30138 2575
rect 30082 2557 30138 2569
rect 30082 2519 30084 2557
rect 30084 2519 30136 2557
rect 30136 2519 30138 2557
rect 30082 2493 30138 2495
rect 30082 2441 30084 2493
rect 30084 2441 30136 2493
rect 30136 2441 30138 2493
rect 30082 2439 30138 2441
rect 30082 2377 30084 2415
rect 30084 2377 30136 2415
rect 30136 2377 30138 2415
rect 30082 2365 30138 2377
rect 30082 2359 30084 2365
rect 30084 2359 30136 2365
rect 30136 2359 30138 2365
rect 30082 2313 30084 2335
rect 30084 2313 30136 2335
rect 30136 2313 30138 2335
rect 30082 2301 30138 2313
rect 30082 2279 30084 2301
rect 30084 2279 30136 2301
rect 30136 2279 30138 2301
rect 30082 2249 30084 2255
rect 30084 2249 30136 2255
rect 30136 2249 30138 2255
rect 30082 2237 30138 2249
rect 30082 2199 30084 2237
rect 30084 2199 30136 2237
rect 30136 2199 30138 2237
rect 30082 2173 30138 2175
rect 30082 2121 30084 2173
rect 30084 2121 30136 2173
rect 30136 2121 30138 2173
rect 30082 2119 30138 2121
rect 30082 2057 30084 2095
rect 30084 2057 30136 2095
rect 30136 2057 30138 2095
rect 30082 2045 30138 2057
rect 30082 2039 30084 2045
rect 30084 2039 30136 2045
rect 30136 2039 30138 2045
rect 30082 1993 30084 2015
rect 30084 1993 30136 2015
rect 30136 1993 30138 2015
rect 30082 1981 30138 1993
rect 30082 1959 30084 1981
rect 30084 1959 30136 1981
rect 30136 1959 30138 1981
rect 30082 1929 30084 1935
rect 30084 1929 30136 1935
rect 30136 1929 30138 1935
rect 30082 1917 30138 1929
rect 30082 1879 30084 1917
rect 30084 1879 30136 1917
rect 30136 1879 30138 1917
rect 30082 1853 30138 1855
rect 30082 1801 30084 1853
rect 30084 1801 30136 1853
rect 30136 1801 30138 1853
rect 30082 1799 30138 1801
rect 30082 1737 30084 1775
rect 30084 1737 30136 1775
rect 30136 1737 30138 1775
rect 30082 1725 30138 1737
rect 30082 1719 30084 1725
rect 30084 1719 30136 1725
rect 30136 1719 30138 1725
rect 30082 1673 30084 1695
rect 30084 1673 30136 1695
rect 30136 1673 30138 1695
rect 30082 1661 30138 1673
rect 30082 1639 30084 1661
rect 30084 1639 30136 1661
rect 30136 1639 30138 1661
rect 30082 1609 30084 1615
rect 30084 1609 30136 1615
rect 30136 1609 30138 1615
rect 30082 1597 30138 1609
rect 30082 1559 30084 1597
rect 30084 1559 30136 1597
rect 30136 1559 30138 1597
rect 30082 1533 30138 1535
rect 30082 1481 30084 1533
rect 30084 1481 30136 1533
rect 30136 1481 30138 1533
rect 30082 1479 30138 1481
rect 30082 1417 30084 1455
rect 30084 1417 30136 1455
rect 30136 1417 30138 1455
rect 30082 1405 30138 1417
rect 30082 1399 30084 1405
rect 30084 1399 30136 1405
rect 30136 1399 30138 1405
rect 30082 1353 30084 1375
rect 30084 1353 30136 1375
rect 30136 1353 30138 1375
rect 30082 1341 30138 1353
rect 30082 1319 30084 1341
rect 30084 1319 30136 1341
rect 30136 1319 30138 1341
rect 30082 1289 30084 1295
rect 30084 1289 30136 1295
rect 30136 1289 30138 1295
rect 30082 1277 30138 1289
rect 30082 1239 30084 1277
rect 30084 1239 30136 1277
rect 30136 1239 30138 1277
rect 30082 1213 30138 1215
rect 30082 1161 30084 1213
rect 30084 1161 30136 1213
rect 30136 1161 30138 1213
rect 30082 1159 30138 1161
rect 30274 3133 30330 3135
rect 30274 3081 30276 3133
rect 30276 3081 30328 3133
rect 30328 3081 30330 3133
rect 30274 3079 30330 3081
rect 30274 3017 30276 3055
rect 30276 3017 30328 3055
rect 30328 3017 30330 3055
rect 30274 3005 30330 3017
rect 30274 2999 30276 3005
rect 30276 2999 30328 3005
rect 30328 2999 30330 3005
rect 30274 2953 30276 2975
rect 30276 2953 30328 2975
rect 30328 2953 30330 2975
rect 30274 2941 30330 2953
rect 30274 2919 30276 2941
rect 30276 2919 30328 2941
rect 30328 2919 30330 2941
rect 30274 2889 30276 2895
rect 30276 2889 30328 2895
rect 30328 2889 30330 2895
rect 30274 2877 30330 2889
rect 30274 2839 30276 2877
rect 30276 2839 30328 2877
rect 30328 2839 30330 2877
rect 30274 2813 30330 2815
rect 30274 2761 30276 2813
rect 30276 2761 30328 2813
rect 30328 2761 30330 2813
rect 30274 2759 30330 2761
rect 30274 2697 30276 2735
rect 30276 2697 30328 2735
rect 30328 2697 30330 2735
rect 30274 2685 30330 2697
rect 30274 2679 30276 2685
rect 30276 2679 30328 2685
rect 30328 2679 30330 2685
rect 30274 2633 30276 2655
rect 30276 2633 30328 2655
rect 30328 2633 30330 2655
rect 30274 2621 30330 2633
rect 30274 2599 30276 2621
rect 30276 2599 30328 2621
rect 30328 2599 30330 2621
rect 30274 2569 30276 2575
rect 30276 2569 30328 2575
rect 30328 2569 30330 2575
rect 30274 2557 30330 2569
rect 30274 2519 30276 2557
rect 30276 2519 30328 2557
rect 30328 2519 30330 2557
rect 30274 2493 30330 2495
rect 30274 2441 30276 2493
rect 30276 2441 30328 2493
rect 30328 2441 30330 2493
rect 30274 2439 30330 2441
rect 30274 2377 30276 2415
rect 30276 2377 30328 2415
rect 30328 2377 30330 2415
rect 30274 2365 30330 2377
rect 30274 2359 30276 2365
rect 30276 2359 30328 2365
rect 30328 2359 30330 2365
rect 30274 2313 30276 2335
rect 30276 2313 30328 2335
rect 30328 2313 30330 2335
rect 30274 2301 30330 2313
rect 30274 2279 30276 2301
rect 30276 2279 30328 2301
rect 30328 2279 30330 2301
rect 30274 2249 30276 2255
rect 30276 2249 30328 2255
rect 30328 2249 30330 2255
rect 30274 2237 30330 2249
rect 30274 2199 30276 2237
rect 30276 2199 30328 2237
rect 30328 2199 30330 2237
rect 30274 2173 30330 2175
rect 30274 2121 30276 2173
rect 30276 2121 30328 2173
rect 30328 2121 30330 2173
rect 30274 2119 30330 2121
rect 30274 2057 30276 2095
rect 30276 2057 30328 2095
rect 30328 2057 30330 2095
rect 30274 2045 30330 2057
rect 30274 2039 30276 2045
rect 30276 2039 30328 2045
rect 30328 2039 30330 2045
rect 30274 1993 30276 2015
rect 30276 1993 30328 2015
rect 30328 1993 30330 2015
rect 30274 1981 30330 1993
rect 30274 1959 30276 1981
rect 30276 1959 30328 1981
rect 30328 1959 30330 1981
rect 30274 1929 30276 1935
rect 30276 1929 30328 1935
rect 30328 1929 30330 1935
rect 30274 1917 30330 1929
rect 30274 1879 30276 1917
rect 30276 1879 30328 1917
rect 30328 1879 30330 1917
rect 30274 1853 30330 1855
rect 30274 1801 30276 1853
rect 30276 1801 30328 1853
rect 30328 1801 30330 1853
rect 30274 1799 30330 1801
rect 30274 1737 30276 1775
rect 30276 1737 30328 1775
rect 30328 1737 30330 1775
rect 30274 1725 30330 1737
rect 30274 1719 30276 1725
rect 30276 1719 30328 1725
rect 30328 1719 30330 1725
rect 30274 1673 30276 1695
rect 30276 1673 30328 1695
rect 30328 1673 30330 1695
rect 30274 1661 30330 1673
rect 30274 1639 30276 1661
rect 30276 1639 30328 1661
rect 30328 1639 30330 1661
rect 30274 1609 30276 1615
rect 30276 1609 30328 1615
rect 30328 1609 30330 1615
rect 30274 1597 30330 1609
rect 30274 1559 30276 1597
rect 30276 1559 30328 1597
rect 30328 1559 30330 1597
rect 30274 1533 30330 1535
rect 30274 1481 30276 1533
rect 30276 1481 30328 1533
rect 30328 1481 30330 1533
rect 30274 1479 30330 1481
rect 30274 1417 30276 1455
rect 30276 1417 30328 1455
rect 30328 1417 30330 1455
rect 30274 1405 30330 1417
rect 30274 1399 30276 1405
rect 30276 1399 30328 1405
rect 30328 1399 30330 1405
rect 30274 1353 30276 1375
rect 30276 1353 30328 1375
rect 30328 1353 30330 1375
rect 30274 1341 30330 1353
rect 30274 1319 30276 1341
rect 30276 1319 30328 1341
rect 30328 1319 30330 1341
rect 30274 1289 30276 1295
rect 30276 1289 30328 1295
rect 30328 1289 30330 1295
rect 30274 1277 30330 1289
rect 30274 1239 30276 1277
rect 30276 1239 30328 1277
rect 30328 1239 30330 1277
rect 30274 1213 30330 1215
rect 30274 1161 30276 1213
rect 30276 1161 30328 1213
rect 30328 1161 30330 1213
rect 30274 1159 30330 1161
rect 30466 3133 30522 3135
rect 30466 3081 30468 3133
rect 30468 3081 30520 3133
rect 30520 3081 30522 3133
rect 30466 3079 30522 3081
rect 30466 3017 30468 3055
rect 30468 3017 30520 3055
rect 30520 3017 30522 3055
rect 30466 3005 30522 3017
rect 30466 2999 30468 3005
rect 30468 2999 30520 3005
rect 30520 2999 30522 3005
rect 30466 2953 30468 2975
rect 30468 2953 30520 2975
rect 30520 2953 30522 2975
rect 30466 2941 30522 2953
rect 30466 2919 30468 2941
rect 30468 2919 30520 2941
rect 30520 2919 30522 2941
rect 30466 2889 30468 2895
rect 30468 2889 30520 2895
rect 30520 2889 30522 2895
rect 30466 2877 30522 2889
rect 30466 2839 30468 2877
rect 30468 2839 30520 2877
rect 30520 2839 30522 2877
rect 30466 2813 30522 2815
rect 30466 2761 30468 2813
rect 30468 2761 30520 2813
rect 30520 2761 30522 2813
rect 30466 2759 30522 2761
rect 30466 2697 30468 2735
rect 30468 2697 30520 2735
rect 30520 2697 30522 2735
rect 30466 2685 30522 2697
rect 30466 2679 30468 2685
rect 30468 2679 30520 2685
rect 30520 2679 30522 2685
rect 30466 2633 30468 2655
rect 30468 2633 30520 2655
rect 30520 2633 30522 2655
rect 30466 2621 30522 2633
rect 30466 2599 30468 2621
rect 30468 2599 30520 2621
rect 30520 2599 30522 2621
rect 30466 2569 30468 2575
rect 30468 2569 30520 2575
rect 30520 2569 30522 2575
rect 30466 2557 30522 2569
rect 30466 2519 30468 2557
rect 30468 2519 30520 2557
rect 30520 2519 30522 2557
rect 30466 2493 30522 2495
rect 30466 2441 30468 2493
rect 30468 2441 30520 2493
rect 30520 2441 30522 2493
rect 30466 2439 30522 2441
rect 30466 2377 30468 2415
rect 30468 2377 30520 2415
rect 30520 2377 30522 2415
rect 30466 2365 30522 2377
rect 30466 2359 30468 2365
rect 30468 2359 30520 2365
rect 30520 2359 30522 2365
rect 30466 2313 30468 2335
rect 30468 2313 30520 2335
rect 30520 2313 30522 2335
rect 30466 2301 30522 2313
rect 30466 2279 30468 2301
rect 30468 2279 30520 2301
rect 30520 2279 30522 2301
rect 30466 2249 30468 2255
rect 30468 2249 30520 2255
rect 30520 2249 30522 2255
rect 30466 2237 30522 2249
rect 30466 2199 30468 2237
rect 30468 2199 30520 2237
rect 30520 2199 30522 2237
rect 30466 2173 30522 2175
rect 30466 2121 30468 2173
rect 30468 2121 30520 2173
rect 30520 2121 30522 2173
rect 30466 2119 30522 2121
rect 30466 2057 30468 2095
rect 30468 2057 30520 2095
rect 30520 2057 30522 2095
rect 30466 2045 30522 2057
rect 30466 2039 30468 2045
rect 30468 2039 30520 2045
rect 30520 2039 30522 2045
rect 30466 1993 30468 2015
rect 30468 1993 30520 2015
rect 30520 1993 30522 2015
rect 30466 1981 30522 1993
rect 30466 1959 30468 1981
rect 30468 1959 30520 1981
rect 30520 1959 30522 1981
rect 30466 1929 30468 1935
rect 30468 1929 30520 1935
rect 30520 1929 30522 1935
rect 30466 1917 30522 1929
rect 30466 1879 30468 1917
rect 30468 1879 30520 1917
rect 30520 1879 30522 1917
rect 30466 1853 30522 1855
rect 30466 1801 30468 1853
rect 30468 1801 30520 1853
rect 30520 1801 30522 1853
rect 30466 1799 30522 1801
rect 30466 1737 30468 1775
rect 30468 1737 30520 1775
rect 30520 1737 30522 1775
rect 30466 1725 30522 1737
rect 30466 1719 30468 1725
rect 30468 1719 30520 1725
rect 30520 1719 30522 1725
rect 30466 1673 30468 1695
rect 30468 1673 30520 1695
rect 30520 1673 30522 1695
rect 30466 1661 30522 1673
rect 30466 1639 30468 1661
rect 30468 1639 30520 1661
rect 30520 1639 30522 1661
rect 30466 1609 30468 1615
rect 30468 1609 30520 1615
rect 30520 1609 30522 1615
rect 30466 1597 30522 1609
rect 30466 1559 30468 1597
rect 30468 1559 30520 1597
rect 30520 1559 30522 1597
rect 30466 1533 30522 1535
rect 30466 1481 30468 1533
rect 30468 1481 30520 1533
rect 30520 1481 30522 1533
rect 30466 1479 30522 1481
rect 30466 1417 30468 1455
rect 30468 1417 30520 1455
rect 30520 1417 30522 1455
rect 30466 1405 30522 1417
rect 30466 1399 30468 1405
rect 30468 1399 30520 1405
rect 30520 1399 30522 1405
rect 30466 1353 30468 1375
rect 30468 1353 30520 1375
rect 30520 1353 30522 1375
rect 30466 1341 30522 1353
rect 30466 1319 30468 1341
rect 30468 1319 30520 1341
rect 30520 1319 30522 1341
rect 30466 1289 30468 1295
rect 30468 1289 30520 1295
rect 30520 1289 30522 1295
rect 30466 1277 30522 1289
rect 30466 1239 30468 1277
rect 30468 1239 30520 1277
rect 30520 1239 30522 1277
rect 30466 1213 30522 1215
rect 30466 1161 30468 1213
rect 30468 1161 30520 1213
rect 30520 1161 30522 1213
rect 30466 1159 30522 1161
rect 30658 3133 30714 3135
rect 30658 3081 30660 3133
rect 30660 3081 30712 3133
rect 30712 3081 30714 3133
rect 30658 3079 30714 3081
rect 30658 3017 30660 3055
rect 30660 3017 30712 3055
rect 30712 3017 30714 3055
rect 30658 3005 30714 3017
rect 30658 2999 30660 3005
rect 30660 2999 30712 3005
rect 30712 2999 30714 3005
rect 30658 2953 30660 2975
rect 30660 2953 30712 2975
rect 30712 2953 30714 2975
rect 30658 2941 30714 2953
rect 30658 2919 30660 2941
rect 30660 2919 30712 2941
rect 30712 2919 30714 2941
rect 30658 2889 30660 2895
rect 30660 2889 30712 2895
rect 30712 2889 30714 2895
rect 30658 2877 30714 2889
rect 30658 2839 30660 2877
rect 30660 2839 30712 2877
rect 30712 2839 30714 2877
rect 30658 2813 30714 2815
rect 30658 2761 30660 2813
rect 30660 2761 30712 2813
rect 30712 2761 30714 2813
rect 30658 2759 30714 2761
rect 30658 2697 30660 2735
rect 30660 2697 30712 2735
rect 30712 2697 30714 2735
rect 30658 2685 30714 2697
rect 30658 2679 30660 2685
rect 30660 2679 30712 2685
rect 30712 2679 30714 2685
rect 30658 2633 30660 2655
rect 30660 2633 30712 2655
rect 30712 2633 30714 2655
rect 30658 2621 30714 2633
rect 30658 2599 30660 2621
rect 30660 2599 30712 2621
rect 30712 2599 30714 2621
rect 30658 2569 30660 2575
rect 30660 2569 30712 2575
rect 30712 2569 30714 2575
rect 30658 2557 30714 2569
rect 30658 2519 30660 2557
rect 30660 2519 30712 2557
rect 30712 2519 30714 2557
rect 30658 2493 30714 2495
rect 30658 2441 30660 2493
rect 30660 2441 30712 2493
rect 30712 2441 30714 2493
rect 30658 2439 30714 2441
rect 30658 2377 30660 2415
rect 30660 2377 30712 2415
rect 30712 2377 30714 2415
rect 30658 2365 30714 2377
rect 30658 2359 30660 2365
rect 30660 2359 30712 2365
rect 30712 2359 30714 2365
rect 30658 2313 30660 2335
rect 30660 2313 30712 2335
rect 30712 2313 30714 2335
rect 30658 2301 30714 2313
rect 30658 2279 30660 2301
rect 30660 2279 30712 2301
rect 30712 2279 30714 2301
rect 30658 2249 30660 2255
rect 30660 2249 30712 2255
rect 30712 2249 30714 2255
rect 30658 2237 30714 2249
rect 30658 2199 30660 2237
rect 30660 2199 30712 2237
rect 30712 2199 30714 2237
rect 30658 2173 30714 2175
rect 30658 2121 30660 2173
rect 30660 2121 30712 2173
rect 30712 2121 30714 2173
rect 30658 2119 30714 2121
rect 30658 2057 30660 2095
rect 30660 2057 30712 2095
rect 30712 2057 30714 2095
rect 30658 2045 30714 2057
rect 30658 2039 30660 2045
rect 30660 2039 30712 2045
rect 30712 2039 30714 2045
rect 30658 1993 30660 2015
rect 30660 1993 30712 2015
rect 30712 1993 30714 2015
rect 30658 1981 30714 1993
rect 30658 1959 30660 1981
rect 30660 1959 30712 1981
rect 30712 1959 30714 1981
rect 30658 1929 30660 1935
rect 30660 1929 30712 1935
rect 30712 1929 30714 1935
rect 30658 1917 30714 1929
rect 30658 1879 30660 1917
rect 30660 1879 30712 1917
rect 30712 1879 30714 1917
rect 30658 1853 30714 1855
rect 30658 1801 30660 1853
rect 30660 1801 30712 1853
rect 30712 1801 30714 1853
rect 30658 1799 30714 1801
rect 30658 1737 30660 1775
rect 30660 1737 30712 1775
rect 30712 1737 30714 1775
rect 30658 1725 30714 1737
rect 30658 1719 30660 1725
rect 30660 1719 30712 1725
rect 30712 1719 30714 1725
rect 30658 1673 30660 1695
rect 30660 1673 30712 1695
rect 30712 1673 30714 1695
rect 30658 1661 30714 1673
rect 30658 1639 30660 1661
rect 30660 1639 30712 1661
rect 30712 1639 30714 1661
rect 30658 1609 30660 1615
rect 30660 1609 30712 1615
rect 30712 1609 30714 1615
rect 30658 1597 30714 1609
rect 30658 1559 30660 1597
rect 30660 1559 30712 1597
rect 30712 1559 30714 1597
rect 30658 1533 30714 1535
rect 30658 1481 30660 1533
rect 30660 1481 30712 1533
rect 30712 1481 30714 1533
rect 30658 1479 30714 1481
rect 30658 1417 30660 1455
rect 30660 1417 30712 1455
rect 30712 1417 30714 1455
rect 30658 1405 30714 1417
rect 30658 1399 30660 1405
rect 30660 1399 30712 1405
rect 30712 1399 30714 1405
rect 30658 1353 30660 1375
rect 30660 1353 30712 1375
rect 30712 1353 30714 1375
rect 30658 1341 30714 1353
rect 30658 1319 30660 1341
rect 30660 1319 30712 1341
rect 30712 1319 30714 1341
rect 30658 1289 30660 1295
rect 30660 1289 30712 1295
rect 30712 1289 30714 1295
rect 30658 1277 30714 1289
rect 30658 1239 30660 1277
rect 30660 1239 30712 1277
rect 30712 1239 30714 1277
rect 30658 1213 30714 1215
rect 30658 1161 30660 1213
rect 30660 1161 30712 1213
rect 30712 1161 30714 1213
rect 30658 1159 30714 1161
rect 30850 3133 30906 3135
rect 30850 3081 30852 3133
rect 30852 3081 30904 3133
rect 30904 3081 30906 3133
rect 30850 3079 30906 3081
rect 30850 3017 30852 3055
rect 30852 3017 30904 3055
rect 30904 3017 30906 3055
rect 30850 3005 30906 3017
rect 30850 2999 30852 3005
rect 30852 2999 30904 3005
rect 30904 2999 30906 3005
rect 30850 2953 30852 2975
rect 30852 2953 30904 2975
rect 30904 2953 30906 2975
rect 30850 2941 30906 2953
rect 30850 2919 30852 2941
rect 30852 2919 30904 2941
rect 30904 2919 30906 2941
rect 30850 2889 30852 2895
rect 30852 2889 30904 2895
rect 30904 2889 30906 2895
rect 30850 2877 30906 2889
rect 30850 2839 30852 2877
rect 30852 2839 30904 2877
rect 30904 2839 30906 2877
rect 30850 2813 30906 2815
rect 30850 2761 30852 2813
rect 30852 2761 30904 2813
rect 30904 2761 30906 2813
rect 30850 2759 30906 2761
rect 30850 2697 30852 2735
rect 30852 2697 30904 2735
rect 30904 2697 30906 2735
rect 30850 2685 30906 2697
rect 30850 2679 30852 2685
rect 30852 2679 30904 2685
rect 30904 2679 30906 2685
rect 30850 2633 30852 2655
rect 30852 2633 30904 2655
rect 30904 2633 30906 2655
rect 30850 2621 30906 2633
rect 30850 2599 30852 2621
rect 30852 2599 30904 2621
rect 30904 2599 30906 2621
rect 30850 2569 30852 2575
rect 30852 2569 30904 2575
rect 30904 2569 30906 2575
rect 30850 2557 30906 2569
rect 30850 2519 30852 2557
rect 30852 2519 30904 2557
rect 30904 2519 30906 2557
rect 30850 2493 30906 2495
rect 30850 2441 30852 2493
rect 30852 2441 30904 2493
rect 30904 2441 30906 2493
rect 30850 2439 30906 2441
rect 30850 2377 30852 2415
rect 30852 2377 30904 2415
rect 30904 2377 30906 2415
rect 30850 2365 30906 2377
rect 30850 2359 30852 2365
rect 30852 2359 30904 2365
rect 30904 2359 30906 2365
rect 30850 2313 30852 2335
rect 30852 2313 30904 2335
rect 30904 2313 30906 2335
rect 30850 2301 30906 2313
rect 30850 2279 30852 2301
rect 30852 2279 30904 2301
rect 30904 2279 30906 2301
rect 30850 2249 30852 2255
rect 30852 2249 30904 2255
rect 30904 2249 30906 2255
rect 30850 2237 30906 2249
rect 30850 2199 30852 2237
rect 30852 2199 30904 2237
rect 30904 2199 30906 2237
rect 30850 2173 30906 2175
rect 30850 2121 30852 2173
rect 30852 2121 30904 2173
rect 30904 2121 30906 2173
rect 30850 2119 30906 2121
rect 30850 2057 30852 2095
rect 30852 2057 30904 2095
rect 30904 2057 30906 2095
rect 30850 2045 30906 2057
rect 30850 2039 30852 2045
rect 30852 2039 30904 2045
rect 30904 2039 30906 2045
rect 30850 1993 30852 2015
rect 30852 1993 30904 2015
rect 30904 1993 30906 2015
rect 30850 1981 30906 1993
rect 30850 1959 30852 1981
rect 30852 1959 30904 1981
rect 30904 1959 30906 1981
rect 30850 1929 30852 1935
rect 30852 1929 30904 1935
rect 30904 1929 30906 1935
rect 30850 1917 30906 1929
rect 30850 1879 30852 1917
rect 30852 1879 30904 1917
rect 30904 1879 30906 1917
rect 30850 1853 30906 1855
rect 30850 1801 30852 1853
rect 30852 1801 30904 1853
rect 30904 1801 30906 1853
rect 30850 1799 30906 1801
rect 30850 1737 30852 1775
rect 30852 1737 30904 1775
rect 30904 1737 30906 1775
rect 30850 1725 30906 1737
rect 30850 1719 30852 1725
rect 30852 1719 30904 1725
rect 30904 1719 30906 1725
rect 30850 1673 30852 1695
rect 30852 1673 30904 1695
rect 30904 1673 30906 1695
rect 30850 1661 30906 1673
rect 30850 1639 30852 1661
rect 30852 1639 30904 1661
rect 30904 1639 30906 1661
rect 30850 1609 30852 1615
rect 30852 1609 30904 1615
rect 30904 1609 30906 1615
rect 30850 1597 30906 1609
rect 30850 1559 30852 1597
rect 30852 1559 30904 1597
rect 30904 1559 30906 1597
rect 30850 1533 30906 1535
rect 30850 1481 30852 1533
rect 30852 1481 30904 1533
rect 30904 1481 30906 1533
rect 30850 1479 30906 1481
rect 30850 1417 30852 1455
rect 30852 1417 30904 1455
rect 30904 1417 30906 1455
rect 30850 1405 30906 1417
rect 30850 1399 30852 1405
rect 30852 1399 30904 1405
rect 30904 1399 30906 1405
rect 30850 1353 30852 1375
rect 30852 1353 30904 1375
rect 30904 1353 30906 1375
rect 30850 1341 30906 1353
rect 30850 1319 30852 1341
rect 30852 1319 30904 1341
rect 30904 1319 30906 1341
rect 30850 1289 30852 1295
rect 30852 1289 30904 1295
rect 30904 1289 30906 1295
rect 30850 1277 30906 1289
rect 30850 1239 30852 1277
rect 30852 1239 30904 1277
rect 30904 1239 30906 1277
rect 30850 1213 30906 1215
rect 30850 1161 30852 1213
rect 30852 1161 30904 1213
rect 30904 1161 30906 1213
rect 30850 1159 30906 1161
rect 31042 3133 31098 3135
rect 31042 3081 31044 3133
rect 31044 3081 31096 3133
rect 31096 3081 31098 3133
rect 31042 3079 31098 3081
rect 31042 3017 31044 3055
rect 31044 3017 31096 3055
rect 31096 3017 31098 3055
rect 31042 3005 31098 3017
rect 31042 2999 31044 3005
rect 31044 2999 31096 3005
rect 31096 2999 31098 3005
rect 31042 2953 31044 2975
rect 31044 2953 31096 2975
rect 31096 2953 31098 2975
rect 31042 2941 31098 2953
rect 31042 2919 31044 2941
rect 31044 2919 31096 2941
rect 31096 2919 31098 2941
rect 31042 2889 31044 2895
rect 31044 2889 31096 2895
rect 31096 2889 31098 2895
rect 31042 2877 31098 2889
rect 31042 2839 31044 2877
rect 31044 2839 31096 2877
rect 31096 2839 31098 2877
rect 31042 2813 31098 2815
rect 31042 2761 31044 2813
rect 31044 2761 31096 2813
rect 31096 2761 31098 2813
rect 31042 2759 31098 2761
rect 31042 2697 31044 2735
rect 31044 2697 31096 2735
rect 31096 2697 31098 2735
rect 31042 2685 31098 2697
rect 31042 2679 31044 2685
rect 31044 2679 31096 2685
rect 31096 2679 31098 2685
rect 31042 2633 31044 2655
rect 31044 2633 31096 2655
rect 31096 2633 31098 2655
rect 31042 2621 31098 2633
rect 31042 2599 31044 2621
rect 31044 2599 31096 2621
rect 31096 2599 31098 2621
rect 31042 2569 31044 2575
rect 31044 2569 31096 2575
rect 31096 2569 31098 2575
rect 31042 2557 31098 2569
rect 31042 2519 31044 2557
rect 31044 2519 31096 2557
rect 31096 2519 31098 2557
rect 31042 2493 31098 2495
rect 31042 2441 31044 2493
rect 31044 2441 31096 2493
rect 31096 2441 31098 2493
rect 31042 2439 31098 2441
rect 31042 2377 31044 2415
rect 31044 2377 31096 2415
rect 31096 2377 31098 2415
rect 31042 2365 31098 2377
rect 31042 2359 31044 2365
rect 31044 2359 31096 2365
rect 31096 2359 31098 2365
rect 31042 2313 31044 2335
rect 31044 2313 31096 2335
rect 31096 2313 31098 2335
rect 31042 2301 31098 2313
rect 31042 2279 31044 2301
rect 31044 2279 31096 2301
rect 31096 2279 31098 2301
rect 31042 2249 31044 2255
rect 31044 2249 31096 2255
rect 31096 2249 31098 2255
rect 31042 2237 31098 2249
rect 31042 2199 31044 2237
rect 31044 2199 31096 2237
rect 31096 2199 31098 2237
rect 31042 2173 31098 2175
rect 31042 2121 31044 2173
rect 31044 2121 31096 2173
rect 31096 2121 31098 2173
rect 31042 2119 31098 2121
rect 31042 2057 31044 2095
rect 31044 2057 31096 2095
rect 31096 2057 31098 2095
rect 31042 2045 31098 2057
rect 31042 2039 31044 2045
rect 31044 2039 31096 2045
rect 31096 2039 31098 2045
rect 31042 1993 31044 2015
rect 31044 1993 31096 2015
rect 31096 1993 31098 2015
rect 31042 1981 31098 1993
rect 31042 1959 31044 1981
rect 31044 1959 31096 1981
rect 31096 1959 31098 1981
rect 31042 1929 31044 1935
rect 31044 1929 31096 1935
rect 31096 1929 31098 1935
rect 31042 1917 31098 1929
rect 31042 1879 31044 1917
rect 31044 1879 31096 1917
rect 31096 1879 31098 1917
rect 31042 1853 31098 1855
rect 31042 1801 31044 1853
rect 31044 1801 31096 1853
rect 31096 1801 31098 1853
rect 31042 1799 31098 1801
rect 31042 1737 31044 1775
rect 31044 1737 31096 1775
rect 31096 1737 31098 1775
rect 31042 1725 31098 1737
rect 31042 1719 31044 1725
rect 31044 1719 31096 1725
rect 31096 1719 31098 1725
rect 31042 1673 31044 1695
rect 31044 1673 31096 1695
rect 31096 1673 31098 1695
rect 31042 1661 31098 1673
rect 31042 1639 31044 1661
rect 31044 1639 31096 1661
rect 31096 1639 31098 1661
rect 31042 1609 31044 1615
rect 31044 1609 31096 1615
rect 31096 1609 31098 1615
rect 31042 1597 31098 1609
rect 31042 1559 31044 1597
rect 31044 1559 31096 1597
rect 31096 1559 31098 1597
rect 31042 1533 31098 1535
rect 31042 1481 31044 1533
rect 31044 1481 31096 1533
rect 31096 1481 31098 1533
rect 31042 1479 31098 1481
rect 31042 1417 31044 1455
rect 31044 1417 31096 1455
rect 31096 1417 31098 1455
rect 31042 1405 31098 1417
rect 31042 1399 31044 1405
rect 31044 1399 31096 1405
rect 31096 1399 31098 1405
rect 31042 1353 31044 1375
rect 31044 1353 31096 1375
rect 31096 1353 31098 1375
rect 31042 1341 31098 1353
rect 31042 1319 31044 1341
rect 31044 1319 31096 1341
rect 31096 1319 31098 1341
rect 31042 1289 31044 1295
rect 31044 1289 31096 1295
rect 31096 1289 31098 1295
rect 31042 1277 31098 1289
rect 31042 1239 31044 1277
rect 31044 1239 31096 1277
rect 31096 1239 31098 1277
rect 31042 1213 31098 1215
rect 31042 1161 31044 1213
rect 31044 1161 31096 1213
rect 31096 1161 31098 1213
rect 31042 1159 31098 1161
rect 31234 3133 31290 3135
rect 31234 3081 31236 3133
rect 31236 3081 31288 3133
rect 31288 3081 31290 3133
rect 31234 3079 31290 3081
rect 31234 3017 31236 3055
rect 31236 3017 31288 3055
rect 31288 3017 31290 3055
rect 31234 3005 31290 3017
rect 31234 2999 31236 3005
rect 31236 2999 31288 3005
rect 31288 2999 31290 3005
rect 31234 2953 31236 2975
rect 31236 2953 31288 2975
rect 31288 2953 31290 2975
rect 31234 2941 31290 2953
rect 31234 2919 31236 2941
rect 31236 2919 31288 2941
rect 31288 2919 31290 2941
rect 31234 2889 31236 2895
rect 31236 2889 31288 2895
rect 31288 2889 31290 2895
rect 31234 2877 31290 2889
rect 31234 2839 31236 2877
rect 31236 2839 31288 2877
rect 31288 2839 31290 2877
rect 31234 2813 31290 2815
rect 31234 2761 31236 2813
rect 31236 2761 31288 2813
rect 31288 2761 31290 2813
rect 31234 2759 31290 2761
rect 31234 2697 31236 2735
rect 31236 2697 31288 2735
rect 31288 2697 31290 2735
rect 31234 2685 31290 2697
rect 31234 2679 31236 2685
rect 31236 2679 31288 2685
rect 31288 2679 31290 2685
rect 31234 2633 31236 2655
rect 31236 2633 31288 2655
rect 31288 2633 31290 2655
rect 31234 2621 31290 2633
rect 31234 2599 31236 2621
rect 31236 2599 31288 2621
rect 31288 2599 31290 2621
rect 31234 2569 31236 2575
rect 31236 2569 31288 2575
rect 31288 2569 31290 2575
rect 31234 2557 31290 2569
rect 31234 2519 31236 2557
rect 31236 2519 31288 2557
rect 31288 2519 31290 2557
rect 31234 2493 31290 2495
rect 31234 2441 31236 2493
rect 31236 2441 31288 2493
rect 31288 2441 31290 2493
rect 31234 2439 31290 2441
rect 31234 2377 31236 2415
rect 31236 2377 31288 2415
rect 31288 2377 31290 2415
rect 31234 2365 31290 2377
rect 31234 2359 31236 2365
rect 31236 2359 31288 2365
rect 31288 2359 31290 2365
rect 31234 2313 31236 2335
rect 31236 2313 31288 2335
rect 31288 2313 31290 2335
rect 31234 2301 31290 2313
rect 31234 2279 31236 2301
rect 31236 2279 31288 2301
rect 31288 2279 31290 2301
rect 31234 2249 31236 2255
rect 31236 2249 31288 2255
rect 31288 2249 31290 2255
rect 31234 2237 31290 2249
rect 31234 2199 31236 2237
rect 31236 2199 31288 2237
rect 31288 2199 31290 2237
rect 31234 2173 31290 2175
rect 31234 2121 31236 2173
rect 31236 2121 31288 2173
rect 31288 2121 31290 2173
rect 31234 2119 31290 2121
rect 31234 2057 31236 2095
rect 31236 2057 31288 2095
rect 31288 2057 31290 2095
rect 31234 2045 31290 2057
rect 31234 2039 31236 2045
rect 31236 2039 31288 2045
rect 31288 2039 31290 2045
rect 31234 1993 31236 2015
rect 31236 1993 31288 2015
rect 31288 1993 31290 2015
rect 31234 1981 31290 1993
rect 31234 1959 31236 1981
rect 31236 1959 31288 1981
rect 31288 1959 31290 1981
rect 31234 1929 31236 1935
rect 31236 1929 31288 1935
rect 31288 1929 31290 1935
rect 31234 1917 31290 1929
rect 31234 1879 31236 1917
rect 31236 1879 31288 1917
rect 31288 1879 31290 1917
rect 31234 1853 31290 1855
rect 31234 1801 31236 1853
rect 31236 1801 31288 1853
rect 31288 1801 31290 1853
rect 31234 1799 31290 1801
rect 31234 1737 31236 1775
rect 31236 1737 31288 1775
rect 31288 1737 31290 1775
rect 31234 1725 31290 1737
rect 31234 1719 31236 1725
rect 31236 1719 31288 1725
rect 31288 1719 31290 1725
rect 31234 1673 31236 1695
rect 31236 1673 31288 1695
rect 31288 1673 31290 1695
rect 31234 1661 31290 1673
rect 31234 1639 31236 1661
rect 31236 1639 31288 1661
rect 31288 1639 31290 1661
rect 31234 1609 31236 1615
rect 31236 1609 31288 1615
rect 31288 1609 31290 1615
rect 31234 1597 31290 1609
rect 31234 1559 31236 1597
rect 31236 1559 31288 1597
rect 31288 1559 31290 1597
rect 31234 1533 31290 1535
rect 31234 1481 31236 1533
rect 31236 1481 31288 1533
rect 31288 1481 31290 1533
rect 31234 1479 31290 1481
rect 31234 1417 31236 1455
rect 31236 1417 31288 1455
rect 31288 1417 31290 1455
rect 31234 1405 31290 1417
rect 31234 1399 31236 1405
rect 31236 1399 31288 1405
rect 31288 1399 31290 1405
rect 31234 1353 31236 1375
rect 31236 1353 31288 1375
rect 31288 1353 31290 1375
rect 31234 1341 31290 1353
rect 31234 1319 31236 1341
rect 31236 1319 31288 1341
rect 31288 1319 31290 1341
rect 31234 1289 31236 1295
rect 31236 1289 31288 1295
rect 31288 1289 31290 1295
rect 31234 1277 31290 1289
rect 31234 1239 31236 1277
rect 31236 1239 31288 1277
rect 31288 1239 31290 1277
rect 31234 1213 31290 1215
rect 31234 1161 31236 1213
rect 31236 1161 31288 1213
rect 31288 1161 31290 1213
rect 31234 1159 31290 1161
rect 31426 3133 31482 3135
rect 31426 3081 31428 3133
rect 31428 3081 31480 3133
rect 31480 3081 31482 3133
rect 31426 3079 31482 3081
rect 31426 3017 31428 3055
rect 31428 3017 31480 3055
rect 31480 3017 31482 3055
rect 31426 3005 31482 3017
rect 31426 2999 31428 3005
rect 31428 2999 31480 3005
rect 31480 2999 31482 3005
rect 31426 2953 31428 2975
rect 31428 2953 31480 2975
rect 31480 2953 31482 2975
rect 31426 2941 31482 2953
rect 31426 2919 31428 2941
rect 31428 2919 31480 2941
rect 31480 2919 31482 2941
rect 31426 2889 31428 2895
rect 31428 2889 31480 2895
rect 31480 2889 31482 2895
rect 31426 2877 31482 2889
rect 31426 2839 31428 2877
rect 31428 2839 31480 2877
rect 31480 2839 31482 2877
rect 31426 2813 31482 2815
rect 31426 2761 31428 2813
rect 31428 2761 31480 2813
rect 31480 2761 31482 2813
rect 31426 2759 31482 2761
rect 31426 2697 31428 2735
rect 31428 2697 31480 2735
rect 31480 2697 31482 2735
rect 31426 2685 31482 2697
rect 31426 2679 31428 2685
rect 31428 2679 31480 2685
rect 31480 2679 31482 2685
rect 31426 2633 31428 2655
rect 31428 2633 31480 2655
rect 31480 2633 31482 2655
rect 31426 2621 31482 2633
rect 31426 2599 31428 2621
rect 31428 2599 31480 2621
rect 31480 2599 31482 2621
rect 31426 2569 31428 2575
rect 31428 2569 31480 2575
rect 31480 2569 31482 2575
rect 31426 2557 31482 2569
rect 31426 2519 31428 2557
rect 31428 2519 31480 2557
rect 31480 2519 31482 2557
rect 31426 2493 31482 2495
rect 31426 2441 31428 2493
rect 31428 2441 31480 2493
rect 31480 2441 31482 2493
rect 31426 2439 31482 2441
rect 31426 2377 31428 2415
rect 31428 2377 31480 2415
rect 31480 2377 31482 2415
rect 31426 2365 31482 2377
rect 31426 2359 31428 2365
rect 31428 2359 31480 2365
rect 31480 2359 31482 2365
rect 31426 2313 31428 2335
rect 31428 2313 31480 2335
rect 31480 2313 31482 2335
rect 31426 2301 31482 2313
rect 31426 2279 31428 2301
rect 31428 2279 31480 2301
rect 31480 2279 31482 2301
rect 31426 2249 31428 2255
rect 31428 2249 31480 2255
rect 31480 2249 31482 2255
rect 31426 2237 31482 2249
rect 31426 2199 31428 2237
rect 31428 2199 31480 2237
rect 31480 2199 31482 2237
rect 31426 2173 31482 2175
rect 31426 2121 31428 2173
rect 31428 2121 31480 2173
rect 31480 2121 31482 2173
rect 31426 2119 31482 2121
rect 31426 2057 31428 2095
rect 31428 2057 31480 2095
rect 31480 2057 31482 2095
rect 31426 2045 31482 2057
rect 31426 2039 31428 2045
rect 31428 2039 31480 2045
rect 31480 2039 31482 2045
rect 31426 1993 31428 2015
rect 31428 1993 31480 2015
rect 31480 1993 31482 2015
rect 31426 1981 31482 1993
rect 31426 1959 31428 1981
rect 31428 1959 31480 1981
rect 31480 1959 31482 1981
rect 31426 1929 31428 1935
rect 31428 1929 31480 1935
rect 31480 1929 31482 1935
rect 31426 1917 31482 1929
rect 31426 1879 31428 1917
rect 31428 1879 31480 1917
rect 31480 1879 31482 1917
rect 31426 1853 31482 1855
rect 31426 1801 31428 1853
rect 31428 1801 31480 1853
rect 31480 1801 31482 1853
rect 31426 1799 31482 1801
rect 31426 1737 31428 1775
rect 31428 1737 31480 1775
rect 31480 1737 31482 1775
rect 31426 1725 31482 1737
rect 31426 1719 31428 1725
rect 31428 1719 31480 1725
rect 31480 1719 31482 1725
rect 31426 1673 31428 1695
rect 31428 1673 31480 1695
rect 31480 1673 31482 1695
rect 31426 1661 31482 1673
rect 31426 1639 31428 1661
rect 31428 1639 31480 1661
rect 31480 1639 31482 1661
rect 31426 1609 31428 1615
rect 31428 1609 31480 1615
rect 31480 1609 31482 1615
rect 31426 1597 31482 1609
rect 31426 1559 31428 1597
rect 31428 1559 31480 1597
rect 31480 1559 31482 1597
rect 31426 1533 31482 1535
rect 31426 1481 31428 1533
rect 31428 1481 31480 1533
rect 31480 1481 31482 1533
rect 31426 1479 31482 1481
rect 31426 1417 31428 1455
rect 31428 1417 31480 1455
rect 31480 1417 31482 1455
rect 31426 1405 31482 1417
rect 31426 1399 31428 1405
rect 31428 1399 31480 1405
rect 31480 1399 31482 1405
rect 31426 1353 31428 1375
rect 31428 1353 31480 1375
rect 31480 1353 31482 1375
rect 31426 1341 31482 1353
rect 31426 1319 31428 1341
rect 31428 1319 31480 1341
rect 31480 1319 31482 1341
rect 31426 1289 31428 1295
rect 31428 1289 31480 1295
rect 31480 1289 31482 1295
rect 31426 1277 31482 1289
rect 31426 1239 31428 1277
rect 31428 1239 31480 1277
rect 31480 1239 31482 1277
rect 31426 1213 31482 1215
rect 31426 1161 31428 1213
rect 31428 1161 31480 1213
rect 31480 1161 31482 1213
rect 31426 1159 31482 1161
rect 31618 3133 31674 3135
rect 31618 3081 31620 3133
rect 31620 3081 31672 3133
rect 31672 3081 31674 3133
rect 31618 3079 31674 3081
rect 31618 3017 31620 3055
rect 31620 3017 31672 3055
rect 31672 3017 31674 3055
rect 31618 3005 31674 3017
rect 31618 2999 31620 3005
rect 31620 2999 31672 3005
rect 31672 2999 31674 3005
rect 31618 2953 31620 2975
rect 31620 2953 31672 2975
rect 31672 2953 31674 2975
rect 31618 2941 31674 2953
rect 31618 2919 31620 2941
rect 31620 2919 31672 2941
rect 31672 2919 31674 2941
rect 31618 2889 31620 2895
rect 31620 2889 31672 2895
rect 31672 2889 31674 2895
rect 31618 2877 31674 2889
rect 31618 2839 31620 2877
rect 31620 2839 31672 2877
rect 31672 2839 31674 2877
rect 31618 2813 31674 2815
rect 31618 2761 31620 2813
rect 31620 2761 31672 2813
rect 31672 2761 31674 2813
rect 31618 2759 31674 2761
rect 31618 2697 31620 2735
rect 31620 2697 31672 2735
rect 31672 2697 31674 2735
rect 31618 2685 31674 2697
rect 31618 2679 31620 2685
rect 31620 2679 31672 2685
rect 31672 2679 31674 2685
rect 31618 2633 31620 2655
rect 31620 2633 31672 2655
rect 31672 2633 31674 2655
rect 31618 2621 31674 2633
rect 31618 2599 31620 2621
rect 31620 2599 31672 2621
rect 31672 2599 31674 2621
rect 31618 2569 31620 2575
rect 31620 2569 31672 2575
rect 31672 2569 31674 2575
rect 31618 2557 31674 2569
rect 31618 2519 31620 2557
rect 31620 2519 31672 2557
rect 31672 2519 31674 2557
rect 31618 2493 31674 2495
rect 31618 2441 31620 2493
rect 31620 2441 31672 2493
rect 31672 2441 31674 2493
rect 31618 2439 31674 2441
rect 31618 2377 31620 2415
rect 31620 2377 31672 2415
rect 31672 2377 31674 2415
rect 31618 2365 31674 2377
rect 31618 2359 31620 2365
rect 31620 2359 31672 2365
rect 31672 2359 31674 2365
rect 31618 2313 31620 2335
rect 31620 2313 31672 2335
rect 31672 2313 31674 2335
rect 31618 2301 31674 2313
rect 31618 2279 31620 2301
rect 31620 2279 31672 2301
rect 31672 2279 31674 2301
rect 31618 2249 31620 2255
rect 31620 2249 31672 2255
rect 31672 2249 31674 2255
rect 31618 2237 31674 2249
rect 31618 2199 31620 2237
rect 31620 2199 31672 2237
rect 31672 2199 31674 2237
rect 31618 2173 31674 2175
rect 31618 2121 31620 2173
rect 31620 2121 31672 2173
rect 31672 2121 31674 2173
rect 31618 2119 31674 2121
rect 31618 2057 31620 2095
rect 31620 2057 31672 2095
rect 31672 2057 31674 2095
rect 31618 2045 31674 2057
rect 31618 2039 31620 2045
rect 31620 2039 31672 2045
rect 31672 2039 31674 2045
rect 31618 1993 31620 2015
rect 31620 1993 31672 2015
rect 31672 1993 31674 2015
rect 31618 1981 31674 1993
rect 31618 1959 31620 1981
rect 31620 1959 31672 1981
rect 31672 1959 31674 1981
rect 31618 1929 31620 1935
rect 31620 1929 31672 1935
rect 31672 1929 31674 1935
rect 31618 1917 31674 1929
rect 31618 1879 31620 1917
rect 31620 1879 31672 1917
rect 31672 1879 31674 1917
rect 31618 1853 31674 1855
rect 31618 1801 31620 1853
rect 31620 1801 31672 1853
rect 31672 1801 31674 1853
rect 31618 1799 31674 1801
rect 31618 1737 31620 1775
rect 31620 1737 31672 1775
rect 31672 1737 31674 1775
rect 31618 1725 31674 1737
rect 31618 1719 31620 1725
rect 31620 1719 31672 1725
rect 31672 1719 31674 1725
rect 31618 1673 31620 1695
rect 31620 1673 31672 1695
rect 31672 1673 31674 1695
rect 31618 1661 31674 1673
rect 31618 1639 31620 1661
rect 31620 1639 31672 1661
rect 31672 1639 31674 1661
rect 31618 1609 31620 1615
rect 31620 1609 31672 1615
rect 31672 1609 31674 1615
rect 31618 1597 31674 1609
rect 31618 1559 31620 1597
rect 31620 1559 31672 1597
rect 31672 1559 31674 1597
rect 31618 1533 31674 1535
rect 31618 1481 31620 1533
rect 31620 1481 31672 1533
rect 31672 1481 31674 1533
rect 31618 1479 31674 1481
rect 31618 1417 31620 1455
rect 31620 1417 31672 1455
rect 31672 1417 31674 1455
rect 31618 1405 31674 1417
rect 31618 1399 31620 1405
rect 31620 1399 31672 1405
rect 31672 1399 31674 1405
rect 31618 1353 31620 1375
rect 31620 1353 31672 1375
rect 31672 1353 31674 1375
rect 31618 1341 31674 1353
rect 31618 1319 31620 1341
rect 31620 1319 31672 1341
rect 31672 1319 31674 1341
rect 31618 1289 31620 1295
rect 31620 1289 31672 1295
rect 31672 1289 31674 1295
rect 31618 1277 31674 1289
rect 31618 1239 31620 1277
rect 31620 1239 31672 1277
rect 31672 1239 31674 1277
rect 31618 1213 31674 1215
rect 31618 1161 31620 1213
rect 31620 1161 31672 1213
rect 31672 1161 31674 1213
rect 31618 1159 31674 1161
rect 31810 3133 31866 3135
rect 31810 3081 31812 3133
rect 31812 3081 31864 3133
rect 31864 3081 31866 3133
rect 31810 3079 31866 3081
rect 31810 3017 31812 3055
rect 31812 3017 31864 3055
rect 31864 3017 31866 3055
rect 31810 3005 31866 3017
rect 31810 2999 31812 3005
rect 31812 2999 31864 3005
rect 31864 2999 31866 3005
rect 31810 2953 31812 2975
rect 31812 2953 31864 2975
rect 31864 2953 31866 2975
rect 31810 2941 31866 2953
rect 31810 2919 31812 2941
rect 31812 2919 31864 2941
rect 31864 2919 31866 2941
rect 31810 2889 31812 2895
rect 31812 2889 31864 2895
rect 31864 2889 31866 2895
rect 31810 2877 31866 2889
rect 31810 2839 31812 2877
rect 31812 2839 31864 2877
rect 31864 2839 31866 2877
rect 31810 2813 31866 2815
rect 31810 2761 31812 2813
rect 31812 2761 31864 2813
rect 31864 2761 31866 2813
rect 31810 2759 31866 2761
rect 31810 2697 31812 2735
rect 31812 2697 31864 2735
rect 31864 2697 31866 2735
rect 31810 2685 31866 2697
rect 31810 2679 31812 2685
rect 31812 2679 31864 2685
rect 31864 2679 31866 2685
rect 31810 2633 31812 2655
rect 31812 2633 31864 2655
rect 31864 2633 31866 2655
rect 31810 2621 31866 2633
rect 31810 2599 31812 2621
rect 31812 2599 31864 2621
rect 31864 2599 31866 2621
rect 31810 2569 31812 2575
rect 31812 2569 31864 2575
rect 31864 2569 31866 2575
rect 31810 2557 31866 2569
rect 31810 2519 31812 2557
rect 31812 2519 31864 2557
rect 31864 2519 31866 2557
rect 31810 2493 31866 2495
rect 31810 2441 31812 2493
rect 31812 2441 31864 2493
rect 31864 2441 31866 2493
rect 31810 2439 31866 2441
rect 31810 2377 31812 2415
rect 31812 2377 31864 2415
rect 31864 2377 31866 2415
rect 31810 2365 31866 2377
rect 31810 2359 31812 2365
rect 31812 2359 31864 2365
rect 31864 2359 31866 2365
rect 31810 2313 31812 2335
rect 31812 2313 31864 2335
rect 31864 2313 31866 2335
rect 31810 2301 31866 2313
rect 31810 2279 31812 2301
rect 31812 2279 31864 2301
rect 31864 2279 31866 2301
rect 31810 2249 31812 2255
rect 31812 2249 31864 2255
rect 31864 2249 31866 2255
rect 31810 2237 31866 2249
rect 31810 2199 31812 2237
rect 31812 2199 31864 2237
rect 31864 2199 31866 2237
rect 31810 2173 31866 2175
rect 31810 2121 31812 2173
rect 31812 2121 31864 2173
rect 31864 2121 31866 2173
rect 31810 2119 31866 2121
rect 31810 2057 31812 2095
rect 31812 2057 31864 2095
rect 31864 2057 31866 2095
rect 31810 2045 31866 2057
rect 31810 2039 31812 2045
rect 31812 2039 31864 2045
rect 31864 2039 31866 2045
rect 31810 1993 31812 2015
rect 31812 1993 31864 2015
rect 31864 1993 31866 2015
rect 31810 1981 31866 1993
rect 31810 1959 31812 1981
rect 31812 1959 31864 1981
rect 31864 1959 31866 1981
rect 31810 1929 31812 1935
rect 31812 1929 31864 1935
rect 31864 1929 31866 1935
rect 31810 1917 31866 1929
rect 31810 1879 31812 1917
rect 31812 1879 31864 1917
rect 31864 1879 31866 1917
rect 31810 1853 31866 1855
rect 31810 1801 31812 1853
rect 31812 1801 31864 1853
rect 31864 1801 31866 1853
rect 31810 1799 31866 1801
rect 31810 1737 31812 1775
rect 31812 1737 31864 1775
rect 31864 1737 31866 1775
rect 31810 1725 31866 1737
rect 31810 1719 31812 1725
rect 31812 1719 31864 1725
rect 31864 1719 31866 1725
rect 31810 1673 31812 1695
rect 31812 1673 31864 1695
rect 31864 1673 31866 1695
rect 31810 1661 31866 1673
rect 31810 1639 31812 1661
rect 31812 1639 31864 1661
rect 31864 1639 31866 1661
rect 31810 1609 31812 1615
rect 31812 1609 31864 1615
rect 31864 1609 31866 1615
rect 31810 1597 31866 1609
rect 31810 1559 31812 1597
rect 31812 1559 31864 1597
rect 31864 1559 31866 1597
rect 31810 1533 31866 1535
rect 31810 1481 31812 1533
rect 31812 1481 31864 1533
rect 31864 1481 31866 1533
rect 31810 1479 31866 1481
rect 31810 1417 31812 1455
rect 31812 1417 31864 1455
rect 31864 1417 31866 1455
rect 31810 1405 31866 1417
rect 31810 1399 31812 1405
rect 31812 1399 31864 1405
rect 31864 1399 31866 1405
rect 31810 1353 31812 1375
rect 31812 1353 31864 1375
rect 31864 1353 31866 1375
rect 31810 1341 31866 1353
rect 31810 1319 31812 1341
rect 31812 1319 31864 1341
rect 31864 1319 31866 1341
rect 31810 1289 31812 1295
rect 31812 1289 31864 1295
rect 31864 1289 31866 1295
rect 31810 1277 31866 1289
rect 31810 1239 31812 1277
rect 31812 1239 31864 1277
rect 31864 1239 31866 1277
rect 31810 1213 31866 1215
rect 31810 1161 31812 1213
rect 31812 1161 31864 1213
rect 31864 1161 31866 1213
rect 31810 1159 31866 1161
rect 32002 3133 32058 3135
rect 32002 3081 32004 3133
rect 32004 3081 32056 3133
rect 32056 3081 32058 3133
rect 32002 3079 32058 3081
rect 32002 3017 32004 3055
rect 32004 3017 32056 3055
rect 32056 3017 32058 3055
rect 32002 3005 32058 3017
rect 32002 2999 32004 3005
rect 32004 2999 32056 3005
rect 32056 2999 32058 3005
rect 32002 2953 32004 2975
rect 32004 2953 32056 2975
rect 32056 2953 32058 2975
rect 32002 2941 32058 2953
rect 32002 2919 32004 2941
rect 32004 2919 32056 2941
rect 32056 2919 32058 2941
rect 32002 2889 32004 2895
rect 32004 2889 32056 2895
rect 32056 2889 32058 2895
rect 32002 2877 32058 2889
rect 32002 2839 32004 2877
rect 32004 2839 32056 2877
rect 32056 2839 32058 2877
rect 32002 2813 32058 2815
rect 32002 2761 32004 2813
rect 32004 2761 32056 2813
rect 32056 2761 32058 2813
rect 32002 2759 32058 2761
rect 32002 2697 32004 2735
rect 32004 2697 32056 2735
rect 32056 2697 32058 2735
rect 32002 2685 32058 2697
rect 32002 2679 32004 2685
rect 32004 2679 32056 2685
rect 32056 2679 32058 2685
rect 32002 2633 32004 2655
rect 32004 2633 32056 2655
rect 32056 2633 32058 2655
rect 32002 2621 32058 2633
rect 32002 2599 32004 2621
rect 32004 2599 32056 2621
rect 32056 2599 32058 2621
rect 32002 2569 32004 2575
rect 32004 2569 32056 2575
rect 32056 2569 32058 2575
rect 32002 2557 32058 2569
rect 32002 2519 32004 2557
rect 32004 2519 32056 2557
rect 32056 2519 32058 2557
rect 32002 2493 32058 2495
rect 32002 2441 32004 2493
rect 32004 2441 32056 2493
rect 32056 2441 32058 2493
rect 32002 2439 32058 2441
rect 32002 2377 32004 2415
rect 32004 2377 32056 2415
rect 32056 2377 32058 2415
rect 32002 2365 32058 2377
rect 32002 2359 32004 2365
rect 32004 2359 32056 2365
rect 32056 2359 32058 2365
rect 32002 2313 32004 2335
rect 32004 2313 32056 2335
rect 32056 2313 32058 2335
rect 32002 2301 32058 2313
rect 32002 2279 32004 2301
rect 32004 2279 32056 2301
rect 32056 2279 32058 2301
rect 32002 2249 32004 2255
rect 32004 2249 32056 2255
rect 32056 2249 32058 2255
rect 32002 2237 32058 2249
rect 32002 2199 32004 2237
rect 32004 2199 32056 2237
rect 32056 2199 32058 2237
rect 32002 2173 32058 2175
rect 32002 2121 32004 2173
rect 32004 2121 32056 2173
rect 32056 2121 32058 2173
rect 32002 2119 32058 2121
rect 32002 2057 32004 2095
rect 32004 2057 32056 2095
rect 32056 2057 32058 2095
rect 32002 2045 32058 2057
rect 32002 2039 32004 2045
rect 32004 2039 32056 2045
rect 32056 2039 32058 2045
rect 32002 1993 32004 2015
rect 32004 1993 32056 2015
rect 32056 1993 32058 2015
rect 32002 1981 32058 1993
rect 32002 1959 32004 1981
rect 32004 1959 32056 1981
rect 32056 1959 32058 1981
rect 32002 1929 32004 1935
rect 32004 1929 32056 1935
rect 32056 1929 32058 1935
rect 32002 1917 32058 1929
rect 32002 1879 32004 1917
rect 32004 1879 32056 1917
rect 32056 1879 32058 1917
rect 32002 1853 32058 1855
rect 32002 1801 32004 1853
rect 32004 1801 32056 1853
rect 32056 1801 32058 1853
rect 32002 1799 32058 1801
rect 32002 1737 32004 1775
rect 32004 1737 32056 1775
rect 32056 1737 32058 1775
rect 32002 1725 32058 1737
rect 32002 1719 32004 1725
rect 32004 1719 32056 1725
rect 32056 1719 32058 1725
rect 32002 1673 32004 1695
rect 32004 1673 32056 1695
rect 32056 1673 32058 1695
rect 32002 1661 32058 1673
rect 32002 1639 32004 1661
rect 32004 1639 32056 1661
rect 32056 1639 32058 1661
rect 32002 1609 32004 1615
rect 32004 1609 32056 1615
rect 32056 1609 32058 1615
rect 32002 1597 32058 1609
rect 32002 1559 32004 1597
rect 32004 1559 32056 1597
rect 32056 1559 32058 1597
rect 32002 1533 32058 1535
rect 32002 1481 32004 1533
rect 32004 1481 32056 1533
rect 32056 1481 32058 1533
rect 32002 1479 32058 1481
rect 32002 1417 32004 1455
rect 32004 1417 32056 1455
rect 32056 1417 32058 1455
rect 32002 1405 32058 1417
rect 32002 1399 32004 1405
rect 32004 1399 32056 1405
rect 32056 1399 32058 1405
rect 32002 1353 32004 1375
rect 32004 1353 32056 1375
rect 32056 1353 32058 1375
rect 32002 1341 32058 1353
rect 32002 1319 32004 1341
rect 32004 1319 32056 1341
rect 32056 1319 32058 1341
rect 32002 1289 32004 1295
rect 32004 1289 32056 1295
rect 32056 1289 32058 1295
rect 32002 1277 32058 1289
rect 32002 1239 32004 1277
rect 32004 1239 32056 1277
rect 32056 1239 32058 1277
rect 32002 1213 32058 1215
rect 32002 1161 32004 1213
rect 32004 1161 32056 1213
rect 32056 1161 32058 1213
rect 32002 1159 32058 1161
rect 32194 3133 32250 3135
rect 32194 3081 32196 3133
rect 32196 3081 32248 3133
rect 32248 3081 32250 3133
rect 32194 3079 32250 3081
rect 32194 3017 32196 3055
rect 32196 3017 32248 3055
rect 32248 3017 32250 3055
rect 32194 3005 32250 3017
rect 32194 2999 32196 3005
rect 32196 2999 32248 3005
rect 32248 2999 32250 3005
rect 32194 2953 32196 2975
rect 32196 2953 32248 2975
rect 32248 2953 32250 2975
rect 32194 2941 32250 2953
rect 32194 2919 32196 2941
rect 32196 2919 32248 2941
rect 32248 2919 32250 2941
rect 32194 2889 32196 2895
rect 32196 2889 32248 2895
rect 32248 2889 32250 2895
rect 32194 2877 32250 2889
rect 32194 2839 32196 2877
rect 32196 2839 32248 2877
rect 32248 2839 32250 2877
rect 32194 2813 32250 2815
rect 32194 2761 32196 2813
rect 32196 2761 32248 2813
rect 32248 2761 32250 2813
rect 32194 2759 32250 2761
rect 32194 2697 32196 2735
rect 32196 2697 32248 2735
rect 32248 2697 32250 2735
rect 32194 2685 32250 2697
rect 32194 2679 32196 2685
rect 32196 2679 32248 2685
rect 32248 2679 32250 2685
rect 32194 2633 32196 2655
rect 32196 2633 32248 2655
rect 32248 2633 32250 2655
rect 32194 2621 32250 2633
rect 32194 2599 32196 2621
rect 32196 2599 32248 2621
rect 32248 2599 32250 2621
rect 32194 2569 32196 2575
rect 32196 2569 32248 2575
rect 32248 2569 32250 2575
rect 32194 2557 32250 2569
rect 32194 2519 32196 2557
rect 32196 2519 32248 2557
rect 32248 2519 32250 2557
rect 32194 2493 32250 2495
rect 32194 2441 32196 2493
rect 32196 2441 32248 2493
rect 32248 2441 32250 2493
rect 32194 2439 32250 2441
rect 32194 2377 32196 2415
rect 32196 2377 32248 2415
rect 32248 2377 32250 2415
rect 32194 2365 32250 2377
rect 32194 2359 32196 2365
rect 32196 2359 32248 2365
rect 32248 2359 32250 2365
rect 32194 2313 32196 2335
rect 32196 2313 32248 2335
rect 32248 2313 32250 2335
rect 32194 2301 32250 2313
rect 32194 2279 32196 2301
rect 32196 2279 32248 2301
rect 32248 2279 32250 2301
rect 32194 2249 32196 2255
rect 32196 2249 32248 2255
rect 32248 2249 32250 2255
rect 32194 2237 32250 2249
rect 32194 2199 32196 2237
rect 32196 2199 32248 2237
rect 32248 2199 32250 2237
rect 32194 2173 32250 2175
rect 32194 2121 32196 2173
rect 32196 2121 32248 2173
rect 32248 2121 32250 2173
rect 32194 2119 32250 2121
rect 32194 2057 32196 2095
rect 32196 2057 32248 2095
rect 32248 2057 32250 2095
rect 32194 2045 32250 2057
rect 32194 2039 32196 2045
rect 32196 2039 32248 2045
rect 32248 2039 32250 2045
rect 32194 1993 32196 2015
rect 32196 1993 32248 2015
rect 32248 1993 32250 2015
rect 32194 1981 32250 1993
rect 32194 1959 32196 1981
rect 32196 1959 32248 1981
rect 32248 1959 32250 1981
rect 32194 1929 32196 1935
rect 32196 1929 32248 1935
rect 32248 1929 32250 1935
rect 32194 1917 32250 1929
rect 32194 1879 32196 1917
rect 32196 1879 32248 1917
rect 32248 1879 32250 1917
rect 32194 1853 32250 1855
rect 32194 1801 32196 1853
rect 32196 1801 32248 1853
rect 32248 1801 32250 1853
rect 32194 1799 32250 1801
rect 32194 1737 32196 1775
rect 32196 1737 32248 1775
rect 32248 1737 32250 1775
rect 32194 1725 32250 1737
rect 32194 1719 32196 1725
rect 32196 1719 32248 1725
rect 32248 1719 32250 1725
rect 32194 1673 32196 1695
rect 32196 1673 32248 1695
rect 32248 1673 32250 1695
rect 32194 1661 32250 1673
rect 32194 1639 32196 1661
rect 32196 1639 32248 1661
rect 32248 1639 32250 1661
rect 32194 1609 32196 1615
rect 32196 1609 32248 1615
rect 32248 1609 32250 1615
rect 32194 1597 32250 1609
rect 32194 1559 32196 1597
rect 32196 1559 32248 1597
rect 32248 1559 32250 1597
rect 32194 1533 32250 1535
rect 32194 1481 32196 1533
rect 32196 1481 32248 1533
rect 32248 1481 32250 1533
rect 32194 1479 32250 1481
rect 32194 1417 32196 1455
rect 32196 1417 32248 1455
rect 32248 1417 32250 1455
rect 32194 1405 32250 1417
rect 32194 1399 32196 1405
rect 32196 1399 32248 1405
rect 32248 1399 32250 1405
rect 32194 1353 32196 1375
rect 32196 1353 32248 1375
rect 32248 1353 32250 1375
rect 32194 1341 32250 1353
rect 32194 1319 32196 1341
rect 32196 1319 32248 1341
rect 32248 1319 32250 1341
rect 32194 1289 32196 1295
rect 32196 1289 32248 1295
rect 32248 1289 32250 1295
rect 32194 1277 32250 1289
rect 32194 1239 32196 1277
rect 32196 1239 32248 1277
rect 32248 1239 32250 1277
rect 32194 1213 32250 1215
rect 32194 1161 32196 1213
rect 32196 1161 32248 1213
rect 32248 1161 32250 1213
rect 32194 1159 32250 1161
rect 32386 3133 32442 3135
rect 32386 3081 32388 3133
rect 32388 3081 32440 3133
rect 32440 3081 32442 3133
rect 32386 3079 32442 3081
rect 32386 3017 32388 3055
rect 32388 3017 32440 3055
rect 32440 3017 32442 3055
rect 32386 3005 32442 3017
rect 32386 2999 32388 3005
rect 32388 2999 32440 3005
rect 32440 2999 32442 3005
rect 32386 2953 32388 2975
rect 32388 2953 32440 2975
rect 32440 2953 32442 2975
rect 32386 2941 32442 2953
rect 32386 2919 32388 2941
rect 32388 2919 32440 2941
rect 32440 2919 32442 2941
rect 32386 2889 32388 2895
rect 32388 2889 32440 2895
rect 32440 2889 32442 2895
rect 32386 2877 32442 2889
rect 32386 2839 32388 2877
rect 32388 2839 32440 2877
rect 32440 2839 32442 2877
rect 32386 2813 32442 2815
rect 32386 2761 32388 2813
rect 32388 2761 32440 2813
rect 32440 2761 32442 2813
rect 32386 2759 32442 2761
rect 32386 2697 32388 2735
rect 32388 2697 32440 2735
rect 32440 2697 32442 2735
rect 32386 2685 32442 2697
rect 32386 2679 32388 2685
rect 32388 2679 32440 2685
rect 32440 2679 32442 2685
rect 32386 2633 32388 2655
rect 32388 2633 32440 2655
rect 32440 2633 32442 2655
rect 32386 2621 32442 2633
rect 32386 2599 32388 2621
rect 32388 2599 32440 2621
rect 32440 2599 32442 2621
rect 32386 2569 32388 2575
rect 32388 2569 32440 2575
rect 32440 2569 32442 2575
rect 32386 2557 32442 2569
rect 32386 2519 32388 2557
rect 32388 2519 32440 2557
rect 32440 2519 32442 2557
rect 32386 2493 32442 2495
rect 32386 2441 32388 2493
rect 32388 2441 32440 2493
rect 32440 2441 32442 2493
rect 32386 2439 32442 2441
rect 32386 2377 32388 2415
rect 32388 2377 32440 2415
rect 32440 2377 32442 2415
rect 32386 2365 32442 2377
rect 32386 2359 32388 2365
rect 32388 2359 32440 2365
rect 32440 2359 32442 2365
rect 32386 2313 32388 2335
rect 32388 2313 32440 2335
rect 32440 2313 32442 2335
rect 32386 2301 32442 2313
rect 32386 2279 32388 2301
rect 32388 2279 32440 2301
rect 32440 2279 32442 2301
rect 32386 2249 32388 2255
rect 32388 2249 32440 2255
rect 32440 2249 32442 2255
rect 32386 2237 32442 2249
rect 32386 2199 32388 2237
rect 32388 2199 32440 2237
rect 32440 2199 32442 2237
rect 32386 2173 32442 2175
rect 32386 2121 32388 2173
rect 32388 2121 32440 2173
rect 32440 2121 32442 2173
rect 32386 2119 32442 2121
rect 32386 2057 32388 2095
rect 32388 2057 32440 2095
rect 32440 2057 32442 2095
rect 32386 2045 32442 2057
rect 32386 2039 32388 2045
rect 32388 2039 32440 2045
rect 32440 2039 32442 2045
rect 32386 1993 32388 2015
rect 32388 1993 32440 2015
rect 32440 1993 32442 2015
rect 32386 1981 32442 1993
rect 32386 1959 32388 1981
rect 32388 1959 32440 1981
rect 32440 1959 32442 1981
rect 32386 1929 32388 1935
rect 32388 1929 32440 1935
rect 32440 1929 32442 1935
rect 32386 1917 32442 1929
rect 32386 1879 32388 1917
rect 32388 1879 32440 1917
rect 32440 1879 32442 1917
rect 32386 1853 32442 1855
rect 32386 1801 32388 1853
rect 32388 1801 32440 1853
rect 32440 1801 32442 1853
rect 32386 1799 32442 1801
rect 32386 1737 32388 1775
rect 32388 1737 32440 1775
rect 32440 1737 32442 1775
rect 32386 1725 32442 1737
rect 32386 1719 32388 1725
rect 32388 1719 32440 1725
rect 32440 1719 32442 1725
rect 32386 1673 32388 1695
rect 32388 1673 32440 1695
rect 32440 1673 32442 1695
rect 32386 1661 32442 1673
rect 32386 1639 32388 1661
rect 32388 1639 32440 1661
rect 32440 1639 32442 1661
rect 32386 1609 32388 1615
rect 32388 1609 32440 1615
rect 32440 1609 32442 1615
rect 32386 1597 32442 1609
rect 32386 1559 32388 1597
rect 32388 1559 32440 1597
rect 32440 1559 32442 1597
rect 32386 1533 32442 1535
rect 32386 1481 32388 1533
rect 32388 1481 32440 1533
rect 32440 1481 32442 1533
rect 32386 1479 32442 1481
rect 32386 1417 32388 1455
rect 32388 1417 32440 1455
rect 32440 1417 32442 1455
rect 32386 1405 32442 1417
rect 32386 1399 32388 1405
rect 32388 1399 32440 1405
rect 32440 1399 32442 1405
rect 32386 1353 32388 1375
rect 32388 1353 32440 1375
rect 32440 1353 32442 1375
rect 32386 1341 32442 1353
rect 32386 1319 32388 1341
rect 32388 1319 32440 1341
rect 32440 1319 32442 1341
rect 32386 1289 32388 1295
rect 32388 1289 32440 1295
rect 32440 1289 32442 1295
rect 32386 1277 32442 1289
rect 32386 1239 32388 1277
rect 32388 1239 32440 1277
rect 32440 1239 32442 1277
rect 32386 1213 32442 1215
rect 32386 1161 32388 1213
rect 32388 1161 32440 1213
rect 32440 1161 32442 1213
rect 32386 1159 32442 1161
rect 32578 3133 32634 3135
rect 32578 3081 32580 3133
rect 32580 3081 32632 3133
rect 32632 3081 32634 3133
rect 32578 3079 32634 3081
rect 32578 3017 32580 3055
rect 32580 3017 32632 3055
rect 32632 3017 32634 3055
rect 32578 3005 32634 3017
rect 32578 2999 32580 3005
rect 32580 2999 32632 3005
rect 32632 2999 32634 3005
rect 32578 2953 32580 2975
rect 32580 2953 32632 2975
rect 32632 2953 32634 2975
rect 32578 2941 32634 2953
rect 32578 2919 32580 2941
rect 32580 2919 32632 2941
rect 32632 2919 32634 2941
rect 32578 2889 32580 2895
rect 32580 2889 32632 2895
rect 32632 2889 32634 2895
rect 32578 2877 32634 2889
rect 32578 2839 32580 2877
rect 32580 2839 32632 2877
rect 32632 2839 32634 2877
rect 32578 2813 32634 2815
rect 32578 2761 32580 2813
rect 32580 2761 32632 2813
rect 32632 2761 32634 2813
rect 32578 2759 32634 2761
rect 32578 2697 32580 2735
rect 32580 2697 32632 2735
rect 32632 2697 32634 2735
rect 32578 2685 32634 2697
rect 32578 2679 32580 2685
rect 32580 2679 32632 2685
rect 32632 2679 32634 2685
rect 32578 2633 32580 2655
rect 32580 2633 32632 2655
rect 32632 2633 32634 2655
rect 32578 2621 32634 2633
rect 32578 2599 32580 2621
rect 32580 2599 32632 2621
rect 32632 2599 32634 2621
rect 32578 2569 32580 2575
rect 32580 2569 32632 2575
rect 32632 2569 32634 2575
rect 32578 2557 32634 2569
rect 32578 2519 32580 2557
rect 32580 2519 32632 2557
rect 32632 2519 32634 2557
rect 32578 2493 32634 2495
rect 32578 2441 32580 2493
rect 32580 2441 32632 2493
rect 32632 2441 32634 2493
rect 32578 2439 32634 2441
rect 32578 2377 32580 2415
rect 32580 2377 32632 2415
rect 32632 2377 32634 2415
rect 32578 2365 32634 2377
rect 32578 2359 32580 2365
rect 32580 2359 32632 2365
rect 32632 2359 32634 2365
rect 32578 2313 32580 2335
rect 32580 2313 32632 2335
rect 32632 2313 32634 2335
rect 32578 2301 32634 2313
rect 32578 2279 32580 2301
rect 32580 2279 32632 2301
rect 32632 2279 32634 2301
rect 32578 2249 32580 2255
rect 32580 2249 32632 2255
rect 32632 2249 32634 2255
rect 32578 2237 32634 2249
rect 32578 2199 32580 2237
rect 32580 2199 32632 2237
rect 32632 2199 32634 2237
rect 32578 2173 32634 2175
rect 32578 2121 32580 2173
rect 32580 2121 32632 2173
rect 32632 2121 32634 2173
rect 32578 2119 32634 2121
rect 32578 2057 32580 2095
rect 32580 2057 32632 2095
rect 32632 2057 32634 2095
rect 32578 2045 32634 2057
rect 32578 2039 32580 2045
rect 32580 2039 32632 2045
rect 32632 2039 32634 2045
rect 32578 1993 32580 2015
rect 32580 1993 32632 2015
rect 32632 1993 32634 2015
rect 32578 1981 32634 1993
rect 32578 1959 32580 1981
rect 32580 1959 32632 1981
rect 32632 1959 32634 1981
rect 32578 1929 32580 1935
rect 32580 1929 32632 1935
rect 32632 1929 32634 1935
rect 32578 1917 32634 1929
rect 32578 1879 32580 1917
rect 32580 1879 32632 1917
rect 32632 1879 32634 1917
rect 32578 1853 32634 1855
rect 32578 1801 32580 1853
rect 32580 1801 32632 1853
rect 32632 1801 32634 1853
rect 32578 1799 32634 1801
rect 32578 1737 32580 1775
rect 32580 1737 32632 1775
rect 32632 1737 32634 1775
rect 32578 1725 32634 1737
rect 32578 1719 32580 1725
rect 32580 1719 32632 1725
rect 32632 1719 32634 1725
rect 32578 1673 32580 1695
rect 32580 1673 32632 1695
rect 32632 1673 32634 1695
rect 32578 1661 32634 1673
rect 32578 1639 32580 1661
rect 32580 1639 32632 1661
rect 32632 1639 32634 1661
rect 32578 1609 32580 1615
rect 32580 1609 32632 1615
rect 32632 1609 32634 1615
rect 32578 1597 32634 1609
rect 32578 1559 32580 1597
rect 32580 1559 32632 1597
rect 32632 1559 32634 1597
rect 32578 1533 32634 1535
rect 32578 1481 32580 1533
rect 32580 1481 32632 1533
rect 32632 1481 32634 1533
rect 32578 1479 32634 1481
rect 32578 1417 32580 1455
rect 32580 1417 32632 1455
rect 32632 1417 32634 1455
rect 32578 1405 32634 1417
rect 32578 1399 32580 1405
rect 32580 1399 32632 1405
rect 32632 1399 32634 1405
rect 32578 1353 32580 1375
rect 32580 1353 32632 1375
rect 32632 1353 32634 1375
rect 32578 1341 32634 1353
rect 32578 1319 32580 1341
rect 32580 1319 32632 1341
rect 32632 1319 32634 1341
rect 32578 1289 32580 1295
rect 32580 1289 32632 1295
rect 32632 1289 32634 1295
rect 32578 1277 32634 1289
rect 32578 1239 32580 1277
rect 32580 1239 32632 1277
rect 32632 1239 32634 1277
rect 32578 1213 32634 1215
rect 32578 1161 32580 1213
rect 32580 1161 32632 1213
rect 32632 1161 32634 1213
rect 32578 1159 32634 1161
rect 32770 3133 32826 3135
rect 32770 3081 32772 3133
rect 32772 3081 32824 3133
rect 32824 3081 32826 3133
rect 32770 3079 32826 3081
rect 32770 3017 32772 3055
rect 32772 3017 32824 3055
rect 32824 3017 32826 3055
rect 32770 3005 32826 3017
rect 32770 2999 32772 3005
rect 32772 2999 32824 3005
rect 32824 2999 32826 3005
rect 32770 2953 32772 2975
rect 32772 2953 32824 2975
rect 32824 2953 32826 2975
rect 32770 2941 32826 2953
rect 32770 2919 32772 2941
rect 32772 2919 32824 2941
rect 32824 2919 32826 2941
rect 32770 2889 32772 2895
rect 32772 2889 32824 2895
rect 32824 2889 32826 2895
rect 32770 2877 32826 2889
rect 32770 2839 32772 2877
rect 32772 2839 32824 2877
rect 32824 2839 32826 2877
rect 32770 2813 32826 2815
rect 32770 2761 32772 2813
rect 32772 2761 32824 2813
rect 32824 2761 32826 2813
rect 32770 2759 32826 2761
rect 32770 2697 32772 2735
rect 32772 2697 32824 2735
rect 32824 2697 32826 2735
rect 32770 2685 32826 2697
rect 32770 2679 32772 2685
rect 32772 2679 32824 2685
rect 32824 2679 32826 2685
rect 32770 2633 32772 2655
rect 32772 2633 32824 2655
rect 32824 2633 32826 2655
rect 32770 2621 32826 2633
rect 32770 2599 32772 2621
rect 32772 2599 32824 2621
rect 32824 2599 32826 2621
rect 32770 2569 32772 2575
rect 32772 2569 32824 2575
rect 32824 2569 32826 2575
rect 32770 2557 32826 2569
rect 32770 2519 32772 2557
rect 32772 2519 32824 2557
rect 32824 2519 32826 2557
rect 32770 2493 32826 2495
rect 32770 2441 32772 2493
rect 32772 2441 32824 2493
rect 32824 2441 32826 2493
rect 32770 2439 32826 2441
rect 32770 2377 32772 2415
rect 32772 2377 32824 2415
rect 32824 2377 32826 2415
rect 32770 2365 32826 2377
rect 32770 2359 32772 2365
rect 32772 2359 32824 2365
rect 32824 2359 32826 2365
rect 32770 2313 32772 2335
rect 32772 2313 32824 2335
rect 32824 2313 32826 2335
rect 32770 2301 32826 2313
rect 32770 2279 32772 2301
rect 32772 2279 32824 2301
rect 32824 2279 32826 2301
rect 32770 2249 32772 2255
rect 32772 2249 32824 2255
rect 32824 2249 32826 2255
rect 32770 2237 32826 2249
rect 32770 2199 32772 2237
rect 32772 2199 32824 2237
rect 32824 2199 32826 2237
rect 32770 2173 32826 2175
rect 32770 2121 32772 2173
rect 32772 2121 32824 2173
rect 32824 2121 32826 2173
rect 32770 2119 32826 2121
rect 32770 2057 32772 2095
rect 32772 2057 32824 2095
rect 32824 2057 32826 2095
rect 32770 2045 32826 2057
rect 32770 2039 32772 2045
rect 32772 2039 32824 2045
rect 32824 2039 32826 2045
rect 32770 1993 32772 2015
rect 32772 1993 32824 2015
rect 32824 1993 32826 2015
rect 32770 1981 32826 1993
rect 32770 1959 32772 1981
rect 32772 1959 32824 1981
rect 32824 1959 32826 1981
rect 32770 1929 32772 1935
rect 32772 1929 32824 1935
rect 32824 1929 32826 1935
rect 32770 1917 32826 1929
rect 32770 1879 32772 1917
rect 32772 1879 32824 1917
rect 32824 1879 32826 1917
rect 32770 1853 32826 1855
rect 32770 1801 32772 1853
rect 32772 1801 32824 1853
rect 32824 1801 32826 1853
rect 32770 1799 32826 1801
rect 32770 1737 32772 1775
rect 32772 1737 32824 1775
rect 32824 1737 32826 1775
rect 32770 1725 32826 1737
rect 32770 1719 32772 1725
rect 32772 1719 32824 1725
rect 32824 1719 32826 1725
rect 32770 1673 32772 1695
rect 32772 1673 32824 1695
rect 32824 1673 32826 1695
rect 32770 1661 32826 1673
rect 32770 1639 32772 1661
rect 32772 1639 32824 1661
rect 32824 1639 32826 1661
rect 32770 1609 32772 1615
rect 32772 1609 32824 1615
rect 32824 1609 32826 1615
rect 32770 1597 32826 1609
rect 32770 1559 32772 1597
rect 32772 1559 32824 1597
rect 32824 1559 32826 1597
rect 32770 1533 32826 1535
rect 32770 1481 32772 1533
rect 32772 1481 32824 1533
rect 32824 1481 32826 1533
rect 32770 1479 32826 1481
rect 32770 1417 32772 1455
rect 32772 1417 32824 1455
rect 32824 1417 32826 1455
rect 32770 1405 32826 1417
rect 32770 1399 32772 1405
rect 32772 1399 32824 1405
rect 32824 1399 32826 1405
rect 32770 1353 32772 1375
rect 32772 1353 32824 1375
rect 32824 1353 32826 1375
rect 32770 1341 32826 1353
rect 32770 1319 32772 1341
rect 32772 1319 32824 1341
rect 32824 1319 32826 1341
rect 32770 1289 32772 1295
rect 32772 1289 32824 1295
rect 32824 1289 32826 1295
rect 32770 1277 32826 1289
rect 32770 1239 32772 1277
rect 32772 1239 32824 1277
rect 32824 1239 32826 1277
rect 32770 1213 32826 1215
rect 32770 1161 32772 1213
rect 32772 1161 32824 1213
rect 32824 1161 32826 1213
rect 32770 1159 32826 1161
rect 32962 3133 33018 3135
rect 32962 3081 32964 3133
rect 32964 3081 33016 3133
rect 33016 3081 33018 3133
rect 32962 3079 33018 3081
rect 32962 3017 32964 3055
rect 32964 3017 33016 3055
rect 33016 3017 33018 3055
rect 32962 3005 33018 3017
rect 32962 2999 32964 3005
rect 32964 2999 33016 3005
rect 33016 2999 33018 3005
rect 32962 2953 32964 2975
rect 32964 2953 33016 2975
rect 33016 2953 33018 2975
rect 32962 2941 33018 2953
rect 32962 2919 32964 2941
rect 32964 2919 33016 2941
rect 33016 2919 33018 2941
rect 32962 2889 32964 2895
rect 32964 2889 33016 2895
rect 33016 2889 33018 2895
rect 32962 2877 33018 2889
rect 32962 2839 32964 2877
rect 32964 2839 33016 2877
rect 33016 2839 33018 2877
rect 32962 2813 33018 2815
rect 32962 2761 32964 2813
rect 32964 2761 33016 2813
rect 33016 2761 33018 2813
rect 32962 2759 33018 2761
rect 32962 2697 32964 2735
rect 32964 2697 33016 2735
rect 33016 2697 33018 2735
rect 32962 2685 33018 2697
rect 32962 2679 32964 2685
rect 32964 2679 33016 2685
rect 33016 2679 33018 2685
rect 32962 2633 32964 2655
rect 32964 2633 33016 2655
rect 33016 2633 33018 2655
rect 32962 2621 33018 2633
rect 32962 2599 32964 2621
rect 32964 2599 33016 2621
rect 33016 2599 33018 2621
rect 32962 2569 32964 2575
rect 32964 2569 33016 2575
rect 33016 2569 33018 2575
rect 32962 2557 33018 2569
rect 32962 2519 32964 2557
rect 32964 2519 33016 2557
rect 33016 2519 33018 2557
rect 32962 2493 33018 2495
rect 32962 2441 32964 2493
rect 32964 2441 33016 2493
rect 33016 2441 33018 2493
rect 32962 2439 33018 2441
rect 32962 2377 32964 2415
rect 32964 2377 33016 2415
rect 33016 2377 33018 2415
rect 32962 2365 33018 2377
rect 32962 2359 32964 2365
rect 32964 2359 33016 2365
rect 33016 2359 33018 2365
rect 32962 2313 32964 2335
rect 32964 2313 33016 2335
rect 33016 2313 33018 2335
rect 32962 2301 33018 2313
rect 32962 2279 32964 2301
rect 32964 2279 33016 2301
rect 33016 2279 33018 2301
rect 32962 2249 32964 2255
rect 32964 2249 33016 2255
rect 33016 2249 33018 2255
rect 32962 2237 33018 2249
rect 32962 2199 32964 2237
rect 32964 2199 33016 2237
rect 33016 2199 33018 2237
rect 32962 2173 33018 2175
rect 32962 2121 32964 2173
rect 32964 2121 33016 2173
rect 33016 2121 33018 2173
rect 32962 2119 33018 2121
rect 32962 2057 32964 2095
rect 32964 2057 33016 2095
rect 33016 2057 33018 2095
rect 32962 2045 33018 2057
rect 32962 2039 32964 2045
rect 32964 2039 33016 2045
rect 33016 2039 33018 2045
rect 32962 1993 32964 2015
rect 32964 1993 33016 2015
rect 33016 1993 33018 2015
rect 32962 1981 33018 1993
rect 32962 1959 32964 1981
rect 32964 1959 33016 1981
rect 33016 1959 33018 1981
rect 32962 1929 32964 1935
rect 32964 1929 33016 1935
rect 33016 1929 33018 1935
rect 32962 1917 33018 1929
rect 32962 1879 32964 1917
rect 32964 1879 33016 1917
rect 33016 1879 33018 1917
rect 32962 1853 33018 1855
rect 32962 1801 32964 1853
rect 32964 1801 33016 1853
rect 33016 1801 33018 1853
rect 32962 1799 33018 1801
rect 32962 1737 32964 1775
rect 32964 1737 33016 1775
rect 33016 1737 33018 1775
rect 32962 1725 33018 1737
rect 32962 1719 32964 1725
rect 32964 1719 33016 1725
rect 33016 1719 33018 1725
rect 32962 1673 32964 1695
rect 32964 1673 33016 1695
rect 33016 1673 33018 1695
rect 32962 1661 33018 1673
rect 32962 1639 32964 1661
rect 32964 1639 33016 1661
rect 33016 1639 33018 1661
rect 32962 1609 32964 1615
rect 32964 1609 33016 1615
rect 33016 1609 33018 1615
rect 32962 1597 33018 1609
rect 32962 1559 32964 1597
rect 32964 1559 33016 1597
rect 33016 1559 33018 1597
rect 32962 1533 33018 1535
rect 32962 1481 32964 1533
rect 32964 1481 33016 1533
rect 33016 1481 33018 1533
rect 32962 1479 33018 1481
rect 32962 1417 32964 1455
rect 32964 1417 33016 1455
rect 33016 1417 33018 1455
rect 32962 1405 33018 1417
rect 32962 1399 32964 1405
rect 32964 1399 33016 1405
rect 33016 1399 33018 1405
rect 32962 1353 32964 1375
rect 32964 1353 33016 1375
rect 33016 1353 33018 1375
rect 32962 1341 33018 1353
rect 32962 1319 32964 1341
rect 32964 1319 33016 1341
rect 33016 1319 33018 1341
rect 32962 1289 32964 1295
rect 32964 1289 33016 1295
rect 33016 1289 33018 1295
rect 32962 1277 33018 1289
rect 32962 1239 32964 1277
rect 32964 1239 33016 1277
rect 33016 1239 33018 1277
rect 32962 1213 33018 1215
rect 32962 1161 32964 1213
rect 32964 1161 33016 1213
rect 33016 1161 33018 1213
rect 32962 1159 33018 1161
rect 33154 3133 33210 3135
rect 33154 3081 33156 3133
rect 33156 3081 33208 3133
rect 33208 3081 33210 3133
rect 33154 3079 33210 3081
rect 33154 3017 33156 3055
rect 33156 3017 33208 3055
rect 33208 3017 33210 3055
rect 33154 3005 33210 3017
rect 33154 2999 33156 3005
rect 33156 2999 33208 3005
rect 33208 2999 33210 3005
rect 33154 2953 33156 2975
rect 33156 2953 33208 2975
rect 33208 2953 33210 2975
rect 33154 2941 33210 2953
rect 33154 2919 33156 2941
rect 33156 2919 33208 2941
rect 33208 2919 33210 2941
rect 33154 2889 33156 2895
rect 33156 2889 33208 2895
rect 33208 2889 33210 2895
rect 33154 2877 33210 2889
rect 33154 2839 33156 2877
rect 33156 2839 33208 2877
rect 33208 2839 33210 2877
rect 33154 2813 33210 2815
rect 33154 2761 33156 2813
rect 33156 2761 33208 2813
rect 33208 2761 33210 2813
rect 33154 2759 33210 2761
rect 33154 2697 33156 2735
rect 33156 2697 33208 2735
rect 33208 2697 33210 2735
rect 33154 2685 33210 2697
rect 33154 2679 33156 2685
rect 33156 2679 33208 2685
rect 33208 2679 33210 2685
rect 33154 2633 33156 2655
rect 33156 2633 33208 2655
rect 33208 2633 33210 2655
rect 33154 2621 33210 2633
rect 33154 2599 33156 2621
rect 33156 2599 33208 2621
rect 33208 2599 33210 2621
rect 33154 2569 33156 2575
rect 33156 2569 33208 2575
rect 33208 2569 33210 2575
rect 33154 2557 33210 2569
rect 33154 2519 33156 2557
rect 33156 2519 33208 2557
rect 33208 2519 33210 2557
rect 33154 2493 33210 2495
rect 33154 2441 33156 2493
rect 33156 2441 33208 2493
rect 33208 2441 33210 2493
rect 33154 2439 33210 2441
rect 33154 2377 33156 2415
rect 33156 2377 33208 2415
rect 33208 2377 33210 2415
rect 33154 2365 33210 2377
rect 33154 2359 33156 2365
rect 33156 2359 33208 2365
rect 33208 2359 33210 2365
rect 33154 2313 33156 2335
rect 33156 2313 33208 2335
rect 33208 2313 33210 2335
rect 33154 2301 33210 2313
rect 33154 2279 33156 2301
rect 33156 2279 33208 2301
rect 33208 2279 33210 2301
rect 33154 2249 33156 2255
rect 33156 2249 33208 2255
rect 33208 2249 33210 2255
rect 33154 2237 33210 2249
rect 33154 2199 33156 2237
rect 33156 2199 33208 2237
rect 33208 2199 33210 2237
rect 33154 2173 33210 2175
rect 33154 2121 33156 2173
rect 33156 2121 33208 2173
rect 33208 2121 33210 2173
rect 33154 2119 33210 2121
rect 33154 2057 33156 2095
rect 33156 2057 33208 2095
rect 33208 2057 33210 2095
rect 33154 2045 33210 2057
rect 33154 2039 33156 2045
rect 33156 2039 33208 2045
rect 33208 2039 33210 2045
rect 33154 1993 33156 2015
rect 33156 1993 33208 2015
rect 33208 1993 33210 2015
rect 33154 1981 33210 1993
rect 33154 1959 33156 1981
rect 33156 1959 33208 1981
rect 33208 1959 33210 1981
rect 33154 1929 33156 1935
rect 33156 1929 33208 1935
rect 33208 1929 33210 1935
rect 33154 1917 33210 1929
rect 33154 1879 33156 1917
rect 33156 1879 33208 1917
rect 33208 1879 33210 1917
rect 33154 1853 33210 1855
rect 33154 1801 33156 1853
rect 33156 1801 33208 1853
rect 33208 1801 33210 1853
rect 33154 1799 33210 1801
rect 33154 1737 33156 1775
rect 33156 1737 33208 1775
rect 33208 1737 33210 1775
rect 33154 1725 33210 1737
rect 33154 1719 33156 1725
rect 33156 1719 33208 1725
rect 33208 1719 33210 1725
rect 33154 1673 33156 1695
rect 33156 1673 33208 1695
rect 33208 1673 33210 1695
rect 33154 1661 33210 1673
rect 33154 1639 33156 1661
rect 33156 1639 33208 1661
rect 33208 1639 33210 1661
rect 33154 1609 33156 1615
rect 33156 1609 33208 1615
rect 33208 1609 33210 1615
rect 33154 1597 33210 1609
rect 33154 1559 33156 1597
rect 33156 1559 33208 1597
rect 33208 1559 33210 1597
rect 33154 1533 33210 1535
rect 33154 1481 33156 1533
rect 33156 1481 33208 1533
rect 33208 1481 33210 1533
rect 33154 1479 33210 1481
rect 33154 1417 33156 1455
rect 33156 1417 33208 1455
rect 33208 1417 33210 1455
rect 33154 1405 33210 1417
rect 33154 1399 33156 1405
rect 33156 1399 33208 1405
rect 33208 1399 33210 1405
rect 33154 1353 33156 1375
rect 33156 1353 33208 1375
rect 33208 1353 33210 1375
rect 33154 1341 33210 1353
rect 33154 1319 33156 1341
rect 33156 1319 33208 1341
rect 33208 1319 33210 1341
rect 33154 1289 33156 1295
rect 33156 1289 33208 1295
rect 33208 1289 33210 1295
rect 33154 1277 33210 1289
rect 33154 1239 33156 1277
rect 33156 1239 33208 1277
rect 33208 1239 33210 1277
rect 33154 1213 33210 1215
rect 33154 1161 33156 1213
rect 33156 1161 33208 1213
rect 33208 1161 33210 1213
rect 33154 1159 33210 1161
rect 33346 3133 33402 3135
rect 33346 3081 33348 3133
rect 33348 3081 33400 3133
rect 33400 3081 33402 3133
rect 33346 3079 33402 3081
rect 33346 3017 33348 3055
rect 33348 3017 33400 3055
rect 33400 3017 33402 3055
rect 33346 3005 33402 3017
rect 33346 2999 33348 3005
rect 33348 2999 33400 3005
rect 33400 2999 33402 3005
rect 33346 2953 33348 2975
rect 33348 2953 33400 2975
rect 33400 2953 33402 2975
rect 33346 2941 33402 2953
rect 33346 2919 33348 2941
rect 33348 2919 33400 2941
rect 33400 2919 33402 2941
rect 33346 2889 33348 2895
rect 33348 2889 33400 2895
rect 33400 2889 33402 2895
rect 33346 2877 33402 2889
rect 33346 2839 33348 2877
rect 33348 2839 33400 2877
rect 33400 2839 33402 2877
rect 33346 2813 33402 2815
rect 33346 2761 33348 2813
rect 33348 2761 33400 2813
rect 33400 2761 33402 2813
rect 33346 2759 33402 2761
rect 33346 2697 33348 2735
rect 33348 2697 33400 2735
rect 33400 2697 33402 2735
rect 33346 2685 33402 2697
rect 33346 2679 33348 2685
rect 33348 2679 33400 2685
rect 33400 2679 33402 2685
rect 33346 2633 33348 2655
rect 33348 2633 33400 2655
rect 33400 2633 33402 2655
rect 33346 2621 33402 2633
rect 33346 2599 33348 2621
rect 33348 2599 33400 2621
rect 33400 2599 33402 2621
rect 33346 2569 33348 2575
rect 33348 2569 33400 2575
rect 33400 2569 33402 2575
rect 33346 2557 33402 2569
rect 33346 2519 33348 2557
rect 33348 2519 33400 2557
rect 33400 2519 33402 2557
rect 33346 2493 33402 2495
rect 33346 2441 33348 2493
rect 33348 2441 33400 2493
rect 33400 2441 33402 2493
rect 33346 2439 33402 2441
rect 33346 2377 33348 2415
rect 33348 2377 33400 2415
rect 33400 2377 33402 2415
rect 33346 2365 33402 2377
rect 33346 2359 33348 2365
rect 33348 2359 33400 2365
rect 33400 2359 33402 2365
rect 33346 2313 33348 2335
rect 33348 2313 33400 2335
rect 33400 2313 33402 2335
rect 33346 2301 33402 2313
rect 33346 2279 33348 2301
rect 33348 2279 33400 2301
rect 33400 2279 33402 2301
rect 33346 2249 33348 2255
rect 33348 2249 33400 2255
rect 33400 2249 33402 2255
rect 33346 2237 33402 2249
rect 33346 2199 33348 2237
rect 33348 2199 33400 2237
rect 33400 2199 33402 2237
rect 33346 2173 33402 2175
rect 33346 2121 33348 2173
rect 33348 2121 33400 2173
rect 33400 2121 33402 2173
rect 33346 2119 33402 2121
rect 33346 2057 33348 2095
rect 33348 2057 33400 2095
rect 33400 2057 33402 2095
rect 33346 2045 33402 2057
rect 33346 2039 33348 2045
rect 33348 2039 33400 2045
rect 33400 2039 33402 2045
rect 33346 1993 33348 2015
rect 33348 1993 33400 2015
rect 33400 1993 33402 2015
rect 33346 1981 33402 1993
rect 33346 1959 33348 1981
rect 33348 1959 33400 1981
rect 33400 1959 33402 1981
rect 33346 1929 33348 1935
rect 33348 1929 33400 1935
rect 33400 1929 33402 1935
rect 33346 1917 33402 1929
rect 33346 1879 33348 1917
rect 33348 1879 33400 1917
rect 33400 1879 33402 1917
rect 33346 1853 33402 1855
rect 33346 1801 33348 1853
rect 33348 1801 33400 1853
rect 33400 1801 33402 1853
rect 33346 1799 33402 1801
rect 33346 1737 33348 1775
rect 33348 1737 33400 1775
rect 33400 1737 33402 1775
rect 33346 1725 33402 1737
rect 33346 1719 33348 1725
rect 33348 1719 33400 1725
rect 33400 1719 33402 1725
rect 33346 1673 33348 1695
rect 33348 1673 33400 1695
rect 33400 1673 33402 1695
rect 33346 1661 33402 1673
rect 33346 1639 33348 1661
rect 33348 1639 33400 1661
rect 33400 1639 33402 1661
rect 33346 1609 33348 1615
rect 33348 1609 33400 1615
rect 33400 1609 33402 1615
rect 33346 1597 33402 1609
rect 33346 1559 33348 1597
rect 33348 1559 33400 1597
rect 33400 1559 33402 1597
rect 33346 1533 33402 1535
rect 33346 1481 33348 1533
rect 33348 1481 33400 1533
rect 33400 1481 33402 1533
rect 33346 1479 33402 1481
rect 33346 1417 33348 1455
rect 33348 1417 33400 1455
rect 33400 1417 33402 1455
rect 33346 1405 33402 1417
rect 33346 1399 33348 1405
rect 33348 1399 33400 1405
rect 33400 1399 33402 1405
rect 33346 1353 33348 1375
rect 33348 1353 33400 1375
rect 33400 1353 33402 1375
rect 33346 1341 33402 1353
rect 33346 1319 33348 1341
rect 33348 1319 33400 1341
rect 33400 1319 33402 1341
rect 33346 1289 33348 1295
rect 33348 1289 33400 1295
rect 33400 1289 33402 1295
rect 33346 1277 33402 1289
rect 33346 1239 33348 1277
rect 33348 1239 33400 1277
rect 33400 1239 33402 1277
rect 33346 1213 33402 1215
rect 33346 1161 33348 1213
rect 33348 1161 33400 1213
rect 33400 1161 33402 1213
rect 33346 1159 33402 1161
rect 33538 3133 33594 3135
rect 33538 3081 33540 3133
rect 33540 3081 33592 3133
rect 33592 3081 33594 3133
rect 33538 3079 33594 3081
rect 33538 3017 33540 3055
rect 33540 3017 33592 3055
rect 33592 3017 33594 3055
rect 33538 3005 33594 3017
rect 33538 2999 33540 3005
rect 33540 2999 33592 3005
rect 33592 2999 33594 3005
rect 33538 2953 33540 2975
rect 33540 2953 33592 2975
rect 33592 2953 33594 2975
rect 33538 2941 33594 2953
rect 33538 2919 33540 2941
rect 33540 2919 33592 2941
rect 33592 2919 33594 2941
rect 33538 2889 33540 2895
rect 33540 2889 33592 2895
rect 33592 2889 33594 2895
rect 33538 2877 33594 2889
rect 33538 2839 33540 2877
rect 33540 2839 33592 2877
rect 33592 2839 33594 2877
rect 33538 2813 33594 2815
rect 33538 2761 33540 2813
rect 33540 2761 33592 2813
rect 33592 2761 33594 2813
rect 33538 2759 33594 2761
rect 33538 2697 33540 2735
rect 33540 2697 33592 2735
rect 33592 2697 33594 2735
rect 33538 2685 33594 2697
rect 33538 2679 33540 2685
rect 33540 2679 33592 2685
rect 33592 2679 33594 2685
rect 33538 2633 33540 2655
rect 33540 2633 33592 2655
rect 33592 2633 33594 2655
rect 33538 2621 33594 2633
rect 33538 2599 33540 2621
rect 33540 2599 33592 2621
rect 33592 2599 33594 2621
rect 33538 2569 33540 2575
rect 33540 2569 33592 2575
rect 33592 2569 33594 2575
rect 33538 2557 33594 2569
rect 33538 2519 33540 2557
rect 33540 2519 33592 2557
rect 33592 2519 33594 2557
rect 33538 2493 33594 2495
rect 33538 2441 33540 2493
rect 33540 2441 33592 2493
rect 33592 2441 33594 2493
rect 33538 2439 33594 2441
rect 33538 2377 33540 2415
rect 33540 2377 33592 2415
rect 33592 2377 33594 2415
rect 33538 2365 33594 2377
rect 33538 2359 33540 2365
rect 33540 2359 33592 2365
rect 33592 2359 33594 2365
rect 33538 2313 33540 2335
rect 33540 2313 33592 2335
rect 33592 2313 33594 2335
rect 33538 2301 33594 2313
rect 33538 2279 33540 2301
rect 33540 2279 33592 2301
rect 33592 2279 33594 2301
rect 33538 2249 33540 2255
rect 33540 2249 33592 2255
rect 33592 2249 33594 2255
rect 33538 2237 33594 2249
rect 33538 2199 33540 2237
rect 33540 2199 33592 2237
rect 33592 2199 33594 2237
rect 33538 2173 33594 2175
rect 33538 2121 33540 2173
rect 33540 2121 33592 2173
rect 33592 2121 33594 2173
rect 33538 2119 33594 2121
rect 33538 2057 33540 2095
rect 33540 2057 33592 2095
rect 33592 2057 33594 2095
rect 33538 2045 33594 2057
rect 33538 2039 33540 2045
rect 33540 2039 33592 2045
rect 33592 2039 33594 2045
rect 33538 1993 33540 2015
rect 33540 1993 33592 2015
rect 33592 1993 33594 2015
rect 33538 1981 33594 1993
rect 33538 1959 33540 1981
rect 33540 1959 33592 1981
rect 33592 1959 33594 1981
rect 33538 1929 33540 1935
rect 33540 1929 33592 1935
rect 33592 1929 33594 1935
rect 33538 1917 33594 1929
rect 33538 1879 33540 1917
rect 33540 1879 33592 1917
rect 33592 1879 33594 1917
rect 33538 1853 33594 1855
rect 33538 1801 33540 1853
rect 33540 1801 33592 1853
rect 33592 1801 33594 1853
rect 33538 1799 33594 1801
rect 33538 1737 33540 1775
rect 33540 1737 33592 1775
rect 33592 1737 33594 1775
rect 33538 1725 33594 1737
rect 33538 1719 33540 1725
rect 33540 1719 33592 1725
rect 33592 1719 33594 1725
rect 33538 1673 33540 1695
rect 33540 1673 33592 1695
rect 33592 1673 33594 1695
rect 33538 1661 33594 1673
rect 33538 1639 33540 1661
rect 33540 1639 33592 1661
rect 33592 1639 33594 1661
rect 33538 1609 33540 1615
rect 33540 1609 33592 1615
rect 33592 1609 33594 1615
rect 33538 1597 33594 1609
rect 33538 1559 33540 1597
rect 33540 1559 33592 1597
rect 33592 1559 33594 1597
rect 33538 1533 33594 1535
rect 33538 1481 33540 1533
rect 33540 1481 33592 1533
rect 33592 1481 33594 1533
rect 33538 1479 33594 1481
rect 33538 1417 33540 1455
rect 33540 1417 33592 1455
rect 33592 1417 33594 1455
rect 33538 1405 33594 1417
rect 33538 1399 33540 1405
rect 33540 1399 33592 1405
rect 33592 1399 33594 1405
rect 33538 1353 33540 1375
rect 33540 1353 33592 1375
rect 33592 1353 33594 1375
rect 33538 1341 33594 1353
rect 33538 1319 33540 1341
rect 33540 1319 33592 1341
rect 33592 1319 33594 1341
rect 33538 1289 33540 1295
rect 33540 1289 33592 1295
rect 33592 1289 33594 1295
rect 33538 1277 33594 1289
rect 33538 1239 33540 1277
rect 33540 1239 33592 1277
rect 33592 1239 33594 1277
rect 33538 1213 33594 1215
rect 33538 1161 33540 1213
rect 33540 1161 33592 1213
rect 33592 1161 33594 1213
rect 33538 1159 33594 1161
rect 33730 3133 33786 3135
rect 33730 3081 33732 3133
rect 33732 3081 33784 3133
rect 33784 3081 33786 3133
rect 33730 3079 33786 3081
rect 33730 3017 33732 3055
rect 33732 3017 33784 3055
rect 33784 3017 33786 3055
rect 33730 3005 33786 3017
rect 33730 2999 33732 3005
rect 33732 2999 33784 3005
rect 33784 2999 33786 3005
rect 33730 2953 33732 2975
rect 33732 2953 33784 2975
rect 33784 2953 33786 2975
rect 33730 2941 33786 2953
rect 33730 2919 33732 2941
rect 33732 2919 33784 2941
rect 33784 2919 33786 2941
rect 33730 2889 33732 2895
rect 33732 2889 33784 2895
rect 33784 2889 33786 2895
rect 33730 2877 33786 2889
rect 33730 2839 33732 2877
rect 33732 2839 33784 2877
rect 33784 2839 33786 2877
rect 33730 2813 33786 2815
rect 33730 2761 33732 2813
rect 33732 2761 33784 2813
rect 33784 2761 33786 2813
rect 33730 2759 33786 2761
rect 33730 2697 33732 2735
rect 33732 2697 33784 2735
rect 33784 2697 33786 2735
rect 33730 2685 33786 2697
rect 33730 2679 33732 2685
rect 33732 2679 33784 2685
rect 33784 2679 33786 2685
rect 33730 2633 33732 2655
rect 33732 2633 33784 2655
rect 33784 2633 33786 2655
rect 33730 2621 33786 2633
rect 33730 2599 33732 2621
rect 33732 2599 33784 2621
rect 33784 2599 33786 2621
rect 33730 2569 33732 2575
rect 33732 2569 33784 2575
rect 33784 2569 33786 2575
rect 33730 2557 33786 2569
rect 33730 2519 33732 2557
rect 33732 2519 33784 2557
rect 33784 2519 33786 2557
rect 33730 2493 33786 2495
rect 33730 2441 33732 2493
rect 33732 2441 33784 2493
rect 33784 2441 33786 2493
rect 33730 2439 33786 2441
rect 33730 2377 33732 2415
rect 33732 2377 33784 2415
rect 33784 2377 33786 2415
rect 33730 2365 33786 2377
rect 33730 2359 33732 2365
rect 33732 2359 33784 2365
rect 33784 2359 33786 2365
rect 33730 2313 33732 2335
rect 33732 2313 33784 2335
rect 33784 2313 33786 2335
rect 33730 2301 33786 2313
rect 33730 2279 33732 2301
rect 33732 2279 33784 2301
rect 33784 2279 33786 2301
rect 33730 2249 33732 2255
rect 33732 2249 33784 2255
rect 33784 2249 33786 2255
rect 33730 2237 33786 2249
rect 33730 2199 33732 2237
rect 33732 2199 33784 2237
rect 33784 2199 33786 2237
rect 33730 2173 33786 2175
rect 33730 2121 33732 2173
rect 33732 2121 33784 2173
rect 33784 2121 33786 2173
rect 33730 2119 33786 2121
rect 33730 2057 33732 2095
rect 33732 2057 33784 2095
rect 33784 2057 33786 2095
rect 33730 2045 33786 2057
rect 33730 2039 33732 2045
rect 33732 2039 33784 2045
rect 33784 2039 33786 2045
rect 33730 1993 33732 2015
rect 33732 1993 33784 2015
rect 33784 1993 33786 2015
rect 33730 1981 33786 1993
rect 33730 1959 33732 1981
rect 33732 1959 33784 1981
rect 33784 1959 33786 1981
rect 33730 1929 33732 1935
rect 33732 1929 33784 1935
rect 33784 1929 33786 1935
rect 33730 1917 33786 1929
rect 33730 1879 33732 1917
rect 33732 1879 33784 1917
rect 33784 1879 33786 1917
rect 33730 1853 33786 1855
rect 33730 1801 33732 1853
rect 33732 1801 33784 1853
rect 33784 1801 33786 1853
rect 33730 1799 33786 1801
rect 33730 1737 33732 1775
rect 33732 1737 33784 1775
rect 33784 1737 33786 1775
rect 33730 1725 33786 1737
rect 33730 1719 33732 1725
rect 33732 1719 33784 1725
rect 33784 1719 33786 1725
rect 33730 1673 33732 1695
rect 33732 1673 33784 1695
rect 33784 1673 33786 1695
rect 33730 1661 33786 1673
rect 33730 1639 33732 1661
rect 33732 1639 33784 1661
rect 33784 1639 33786 1661
rect 33730 1609 33732 1615
rect 33732 1609 33784 1615
rect 33784 1609 33786 1615
rect 33730 1597 33786 1609
rect 33730 1559 33732 1597
rect 33732 1559 33784 1597
rect 33784 1559 33786 1597
rect 33730 1533 33786 1535
rect 33730 1481 33732 1533
rect 33732 1481 33784 1533
rect 33784 1481 33786 1533
rect 33730 1479 33786 1481
rect 33730 1417 33732 1455
rect 33732 1417 33784 1455
rect 33784 1417 33786 1455
rect 33730 1405 33786 1417
rect 33730 1399 33732 1405
rect 33732 1399 33784 1405
rect 33784 1399 33786 1405
rect 33730 1353 33732 1375
rect 33732 1353 33784 1375
rect 33784 1353 33786 1375
rect 33730 1341 33786 1353
rect 33730 1319 33732 1341
rect 33732 1319 33784 1341
rect 33784 1319 33786 1341
rect 33730 1289 33732 1295
rect 33732 1289 33784 1295
rect 33784 1289 33786 1295
rect 33730 1277 33786 1289
rect 33730 1239 33732 1277
rect 33732 1239 33784 1277
rect 33784 1239 33786 1277
rect 33730 1213 33786 1215
rect 33730 1161 33732 1213
rect 33732 1161 33784 1213
rect 33784 1161 33786 1213
rect 33730 1159 33786 1161
rect 33922 3133 33978 3135
rect 33922 3081 33924 3133
rect 33924 3081 33976 3133
rect 33976 3081 33978 3133
rect 33922 3079 33978 3081
rect 33922 3017 33924 3055
rect 33924 3017 33976 3055
rect 33976 3017 33978 3055
rect 33922 3005 33978 3017
rect 33922 2999 33924 3005
rect 33924 2999 33976 3005
rect 33976 2999 33978 3005
rect 33922 2953 33924 2975
rect 33924 2953 33976 2975
rect 33976 2953 33978 2975
rect 33922 2941 33978 2953
rect 33922 2919 33924 2941
rect 33924 2919 33976 2941
rect 33976 2919 33978 2941
rect 33922 2889 33924 2895
rect 33924 2889 33976 2895
rect 33976 2889 33978 2895
rect 33922 2877 33978 2889
rect 33922 2839 33924 2877
rect 33924 2839 33976 2877
rect 33976 2839 33978 2877
rect 33922 2813 33978 2815
rect 33922 2761 33924 2813
rect 33924 2761 33976 2813
rect 33976 2761 33978 2813
rect 33922 2759 33978 2761
rect 33922 2697 33924 2735
rect 33924 2697 33976 2735
rect 33976 2697 33978 2735
rect 33922 2685 33978 2697
rect 33922 2679 33924 2685
rect 33924 2679 33976 2685
rect 33976 2679 33978 2685
rect 33922 2633 33924 2655
rect 33924 2633 33976 2655
rect 33976 2633 33978 2655
rect 33922 2621 33978 2633
rect 33922 2599 33924 2621
rect 33924 2599 33976 2621
rect 33976 2599 33978 2621
rect 33922 2569 33924 2575
rect 33924 2569 33976 2575
rect 33976 2569 33978 2575
rect 33922 2557 33978 2569
rect 33922 2519 33924 2557
rect 33924 2519 33976 2557
rect 33976 2519 33978 2557
rect 33922 2493 33978 2495
rect 33922 2441 33924 2493
rect 33924 2441 33976 2493
rect 33976 2441 33978 2493
rect 33922 2439 33978 2441
rect 33922 2377 33924 2415
rect 33924 2377 33976 2415
rect 33976 2377 33978 2415
rect 33922 2365 33978 2377
rect 33922 2359 33924 2365
rect 33924 2359 33976 2365
rect 33976 2359 33978 2365
rect 33922 2313 33924 2335
rect 33924 2313 33976 2335
rect 33976 2313 33978 2335
rect 33922 2301 33978 2313
rect 33922 2279 33924 2301
rect 33924 2279 33976 2301
rect 33976 2279 33978 2301
rect 33922 2249 33924 2255
rect 33924 2249 33976 2255
rect 33976 2249 33978 2255
rect 33922 2237 33978 2249
rect 33922 2199 33924 2237
rect 33924 2199 33976 2237
rect 33976 2199 33978 2237
rect 33922 2173 33978 2175
rect 33922 2121 33924 2173
rect 33924 2121 33976 2173
rect 33976 2121 33978 2173
rect 33922 2119 33978 2121
rect 33922 2057 33924 2095
rect 33924 2057 33976 2095
rect 33976 2057 33978 2095
rect 33922 2045 33978 2057
rect 33922 2039 33924 2045
rect 33924 2039 33976 2045
rect 33976 2039 33978 2045
rect 33922 1993 33924 2015
rect 33924 1993 33976 2015
rect 33976 1993 33978 2015
rect 33922 1981 33978 1993
rect 33922 1959 33924 1981
rect 33924 1959 33976 1981
rect 33976 1959 33978 1981
rect 33922 1929 33924 1935
rect 33924 1929 33976 1935
rect 33976 1929 33978 1935
rect 33922 1917 33978 1929
rect 33922 1879 33924 1917
rect 33924 1879 33976 1917
rect 33976 1879 33978 1917
rect 33922 1853 33978 1855
rect 33922 1801 33924 1853
rect 33924 1801 33976 1853
rect 33976 1801 33978 1853
rect 33922 1799 33978 1801
rect 33922 1737 33924 1775
rect 33924 1737 33976 1775
rect 33976 1737 33978 1775
rect 33922 1725 33978 1737
rect 33922 1719 33924 1725
rect 33924 1719 33976 1725
rect 33976 1719 33978 1725
rect 33922 1673 33924 1695
rect 33924 1673 33976 1695
rect 33976 1673 33978 1695
rect 33922 1661 33978 1673
rect 33922 1639 33924 1661
rect 33924 1639 33976 1661
rect 33976 1639 33978 1661
rect 33922 1609 33924 1615
rect 33924 1609 33976 1615
rect 33976 1609 33978 1615
rect 33922 1597 33978 1609
rect 33922 1559 33924 1597
rect 33924 1559 33976 1597
rect 33976 1559 33978 1597
rect 33922 1533 33978 1535
rect 33922 1481 33924 1533
rect 33924 1481 33976 1533
rect 33976 1481 33978 1533
rect 33922 1479 33978 1481
rect 33922 1417 33924 1455
rect 33924 1417 33976 1455
rect 33976 1417 33978 1455
rect 33922 1405 33978 1417
rect 33922 1399 33924 1405
rect 33924 1399 33976 1405
rect 33976 1399 33978 1405
rect 33922 1353 33924 1375
rect 33924 1353 33976 1375
rect 33976 1353 33978 1375
rect 33922 1341 33978 1353
rect 33922 1319 33924 1341
rect 33924 1319 33976 1341
rect 33976 1319 33978 1341
rect 33922 1289 33924 1295
rect 33924 1289 33976 1295
rect 33976 1289 33978 1295
rect 33922 1277 33978 1289
rect 33922 1239 33924 1277
rect 33924 1239 33976 1277
rect 33976 1239 33978 1277
rect 33922 1213 33978 1215
rect 33922 1161 33924 1213
rect 33924 1161 33976 1213
rect 33976 1161 33978 1213
rect 33922 1159 33978 1161
rect 34114 3133 34170 3135
rect 34114 3081 34116 3133
rect 34116 3081 34168 3133
rect 34168 3081 34170 3133
rect 34114 3079 34170 3081
rect 34114 3017 34116 3055
rect 34116 3017 34168 3055
rect 34168 3017 34170 3055
rect 34114 3005 34170 3017
rect 34114 2999 34116 3005
rect 34116 2999 34168 3005
rect 34168 2999 34170 3005
rect 34114 2953 34116 2975
rect 34116 2953 34168 2975
rect 34168 2953 34170 2975
rect 34114 2941 34170 2953
rect 34114 2919 34116 2941
rect 34116 2919 34168 2941
rect 34168 2919 34170 2941
rect 34114 2889 34116 2895
rect 34116 2889 34168 2895
rect 34168 2889 34170 2895
rect 34114 2877 34170 2889
rect 34114 2839 34116 2877
rect 34116 2839 34168 2877
rect 34168 2839 34170 2877
rect 34114 2813 34170 2815
rect 34114 2761 34116 2813
rect 34116 2761 34168 2813
rect 34168 2761 34170 2813
rect 34114 2759 34170 2761
rect 34114 2697 34116 2735
rect 34116 2697 34168 2735
rect 34168 2697 34170 2735
rect 34114 2685 34170 2697
rect 34114 2679 34116 2685
rect 34116 2679 34168 2685
rect 34168 2679 34170 2685
rect 34114 2633 34116 2655
rect 34116 2633 34168 2655
rect 34168 2633 34170 2655
rect 34114 2621 34170 2633
rect 34114 2599 34116 2621
rect 34116 2599 34168 2621
rect 34168 2599 34170 2621
rect 34114 2569 34116 2575
rect 34116 2569 34168 2575
rect 34168 2569 34170 2575
rect 34114 2557 34170 2569
rect 34114 2519 34116 2557
rect 34116 2519 34168 2557
rect 34168 2519 34170 2557
rect 34114 2493 34170 2495
rect 34114 2441 34116 2493
rect 34116 2441 34168 2493
rect 34168 2441 34170 2493
rect 34114 2439 34170 2441
rect 34114 2377 34116 2415
rect 34116 2377 34168 2415
rect 34168 2377 34170 2415
rect 34114 2365 34170 2377
rect 34114 2359 34116 2365
rect 34116 2359 34168 2365
rect 34168 2359 34170 2365
rect 34114 2313 34116 2335
rect 34116 2313 34168 2335
rect 34168 2313 34170 2335
rect 34114 2301 34170 2313
rect 34114 2279 34116 2301
rect 34116 2279 34168 2301
rect 34168 2279 34170 2301
rect 34114 2249 34116 2255
rect 34116 2249 34168 2255
rect 34168 2249 34170 2255
rect 34114 2237 34170 2249
rect 34114 2199 34116 2237
rect 34116 2199 34168 2237
rect 34168 2199 34170 2237
rect 34114 2173 34170 2175
rect 34114 2121 34116 2173
rect 34116 2121 34168 2173
rect 34168 2121 34170 2173
rect 34114 2119 34170 2121
rect 34114 2057 34116 2095
rect 34116 2057 34168 2095
rect 34168 2057 34170 2095
rect 34114 2045 34170 2057
rect 34114 2039 34116 2045
rect 34116 2039 34168 2045
rect 34168 2039 34170 2045
rect 34114 1993 34116 2015
rect 34116 1993 34168 2015
rect 34168 1993 34170 2015
rect 34114 1981 34170 1993
rect 34114 1959 34116 1981
rect 34116 1959 34168 1981
rect 34168 1959 34170 1981
rect 34114 1929 34116 1935
rect 34116 1929 34168 1935
rect 34168 1929 34170 1935
rect 34114 1917 34170 1929
rect 34114 1879 34116 1917
rect 34116 1879 34168 1917
rect 34168 1879 34170 1917
rect 34114 1853 34170 1855
rect 34114 1801 34116 1853
rect 34116 1801 34168 1853
rect 34168 1801 34170 1853
rect 34114 1799 34170 1801
rect 34114 1737 34116 1775
rect 34116 1737 34168 1775
rect 34168 1737 34170 1775
rect 34114 1725 34170 1737
rect 34114 1719 34116 1725
rect 34116 1719 34168 1725
rect 34168 1719 34170 1725
rect 34114 1673 34116 1695
rect 34116 1673 34168 1695
rect 34168 1673 34170 1695
rect 34114 1661 34170 1673
rect 34114 1639 34116 1661
rect 34116 1639 34168 1661
rect 34168 1639 34170 1661
rect 34114 1609 34116 1615
rect 34116 1609 34168 1615
rect 34168 1609 34170 1615
rect 34114 1597 34170 1609
rect 34114 1559 34116 1597
rect 34116 1559 34168 1597
rect 34168 1559 34170 1597
rect 34114 1533 34170 1535
rect 34114 1481 34116 1533
rect 34116 1481 34168 1533
rect 34168 1481 34170 1533
rect 34114 1479 34170 1481
rect 34114 1417 34116 1455
rect 34116 1417 34168 1455
rect 34168 1417 34170 1455
rect 34114 1405 34170 1417
rect 34114 1399 34116 1405
rect 34116 1399 34168 1405
rect 34168 1399 34170 1405
rect 34114 1353 34116 1375
rect 34116 1353 34168 1375
rect 34168 1353 34170 1375
rect 34114 1341 34170 1353
rect 34114 1319 34116 1341
rect 34116 1319 34168 1341
rect 34168 1319 34170 1341
rect 34114 1289 34116 1295
rect 34116 1289 34168 1295
rect 34168 1289 34170 1295
rect 34114 1277 34170 1289
rect 34114 1239 34116 1277
rect 34116 1239 34168 1277
rect 34168 1239 34170 1277
rect 34114 1213 34170 1215
rect 34114 1161 34116 1213
rect 34116 1161 34168 1213
rect 34168 1161 34170 1213
rect 34114 1159 34170 1161
rect 34306 3133 34362 3135
rect 34306 3081 34308 3133
rect 34308 3081 34360 3133
rect 34360 3081 34362 3133
rect 34306 3079 34362 3081
rect 34306 3017 34308 3055
rect 34308 3017 34360 3055
rect 34360 3017 34362 3055
rect 34306 3005 34362 3017
rect 34306 2999 34308 3005
rect 34308 2999 34360 3005
rect 34360 2999 34362 3005
rect 34306 2953 34308 2975
rect 34308 2953 34360 2975
rect 34360 2953 34362 2975
rect 34306 2941 34362 2953
rect 34306 2919 34308 2941
rect 34308 2919 34360 2941
rect 34360 2919 34362 2941
rect 34306 2889 34308 2895
rect 34308 2889 34360 2895
rect 34360 2889 34362 2895
rect 34306 2877 34362 2889
rect 34306 2839 34308 2877
rect 34308 2839 34360 2877
rect 34360 2839 34362 2877
rect 34306 2813 34362 2815
rect 34306 2761 34308 2813
rect 34308 2761 34360 2813
rect 34360 2761 34362 2813
rect 34306 2759 34362 2761
rect 34306 2697 34308 2735
rect 34308 2697 34360 2735
rect 34360 2697 34362 2735
rect 34306 2685 34362 2697
rect 34306 2679 34308 2685
rect 34308 2679 34360 2685
rect 34360 2679 34362 2685
rect 34306 2633 34308 2655
rect 34308 2633 34360 2655
rect 34360 2633 34362 2655
rect 34306 2621 34362 2633
rect 34306 2599 34308 2621
rect 34308 2599 34360 2621
rect 34360 2599 34362 2621
rect 34306 2569 34308 2575
rect 34308 2569 34360 2575
rect 34360 2569 34362 2575
rect 34306 2557 34362 2569
rect 34306 2519 34308 2557
rect 34308 2519 34360 2557
rect 34360 2519 34362 2557
rect 34306 2493 34362 2495
rect 34306 2441 34308 2493
rect 34308 2441 34360 2493
rect 34360 2441 34362 2493
rect 34306 2439 34362 2441
rect 34306 2377 34308 2415
rect 34308 2377 34360 2415
rect 34360 2377 34362 2415
rect 34306 2365 34362 2377
rect 34306 2359 34308 2365
rect 34308 2359 34360 2365
rect 34360 2359 34362 2365
rect 34306 2313 34308 2335
rect 34308 2313 34360 2335
rect 34360 2313 34362 2335
rect 34306 2301 34362 2313
rect 34306 2279 34308 2301
rect 34308 2279 34360 2301
rect 34360 2279 34362 2301
rect 34306 2249 34308 2255
rect 34308 2249 34360 2255
rect 34360 2249 34362 2255
rect 34306 2237 34362 2249
rect 34306 2199 34308 2237
rect 34308 2199 34360 2237
rect 34360 2199 34362 2237
rect 34306 2173 34362 2175
rect 34306 2121 34308 2173
rect 34308 2121 34360 2173
rect 34360 2121 34362 2173
rect 34306 2119 34362 2121
rect 34306 2057 34308 2095
rect 34308 2057 34360 2095
rect 34360 2057 34362 2095
rect 34306 2045 34362 2057
rect 34306 2039 34308 2045
rect 34308 2039 34360 2045
rect 34360 2039 34362 2045
rect 34306 1993 34308 2015
rect 34308 1993 34360 2015
rect 34360 1993 34362 2015
rect 34306 1981 34362 1993
rect 34306 1959 34308 1981
rect 34308 1959 34360 1981
rect 34360 1959 34362 1981
rect 34306 1929 34308 1935
rect 34308 1929 34360 1935
rect 34360 1929 34362 1935
rect 34306 1917 34362 1929
rect 34306 1879 34308 1917
rect 34308 1879 34360 1917
rect 34360 1879 34362 1917
rect 34306 1853 34362 1855
rect 34306 1801 34308 1853
rect 34308 1801 34360 1853
rect 34360 1801 34362 1853
rect 34306 1799 34362 1801
rect 34306 1737 34308 1775
rect 34308 1737 34360 1775
rect 34360 1737 34362 1775
rect 34306 1725 34362 1737
rect 34306 1719 34308 1725
rect 34308 1719 34360 1725
rect 34360 1719 34362 1725
rect 34306 1673 34308 1695
rect 34308 1673 34360 1695
rect 34360 1673 34362 1695
rect 34306 1661 34362 1673
rect 34306 1639 34308 1661
rect 34308 1639 34360 1661
rect 34360 1639 34362 1661
rect 34306 1609 34308 1615
rect 34308 1609 34360 1615
rect 34360 1609 34362 1615
rect 34306 1597 34362 1609
rect 34306 1559 34308 1597
rect 34308 1559 34360 1597
rect 34360 1559 34362 1597
rect 34306 1533 34362 1535
rect 34306 1481 34308 1533
rect 34308 1481 34360 1533
rect 34360 1481 34362 1533
rect 34306 1479 34362 1481
rect 34306 1417 34308 1455
rect 34308 1417 34360 1455
rect 34360 1417 34362 1455
rect 34306 1405 34362 1417
rect 34306 1399 34308 1405
rect 34308 1399 34360 1405
rect 34360 1399 34362 1405
rect 34306 1353 34308 1375
rect 34308 1353 34360 1375
rect 34360 1353 34362 1375
rect 34306 1341 34362 1353
rect 34306 1319 34308 1341
rect 34308 1319 34360 1341
rect 34360 1319 34362 1341
rect 34306 1289 34308 1295
rect 34308 1289 34360 1295
rect 34360 1289 34362 1295
rect 34306 1277 34362 1289
rect 34306 1239 34308 1277
rect 34308 1239 34360 1277
rect 34360 1239 34362 1277
rect 34306 1213 34362 1215
rect 34306 1161 34308 1213
rect 34308 1161 34360 1213
rect 34360 1161 34362 1213
rect 34306 1159 34362 1161
rect 34498 3133 34554 3135
rect 34498 3081 34500 3133
rect 34500 3081 34552 3133
rect 34552 3081 34554 3133
rect 34498 3079 34554 3081
rect 34498 3017 34500 3055
rect 34500 3017 34552 3055
rect 34552 3017 34554 3055
rect 34498 3005 34554 3017
rect 34498 2999 34500 3005
rect 34500 2999 34552 3005
rect 34552 2999 34554 3005
rect 34498 2953 34500 2975
rect 34500 2953 34552 2975
rect 34552 2953 34554 2975
rect 34498 2941 34554 2953
rect 34498 2919 34500 2941
rect 34500 2919 34552 2941
rect 34552 2919 34554 2941
rect 34498 2889 34500 2895
rect 34500 2889 34552 2895
rect 34552 2889 34554 2895
rect 34498 2877 34554 2889
rect 34498 2839 34500 2877
rect 34500 2839 34552 2877
rect 34552 2839 34554 2877
rect 34498 2813 34554 2815
rect 34498 2761 34500 2813
rect 34500 2761 34552 2813
rect 34552 2761 34554 2813
rect 34498 2759 34554 2761
rect 34498 2697 34500 2735
rect 34500 2697 34552 2735
rect 34552 2697 34554 2735
rect 34498 2685 34554 2697
rect 34498 2679 34500 2685
rect 34500 2679 34552 2685
rect 34552 2679 34554 2685
rect 34498 2633 34500 2655
rect 34500 2633 34552 2655
rect 34552 2633 34554 2655
rect 34498 2621 34554 2633
rect 34498 2599 34500 2621
rect 34500 2599 34552 2621
rect 34552 2599 34554 2621
rect 34498 2569 34500 2575
rect 34500 2569 34552 2575
rect 34552 2569 34554 2575
rect 34498 2557 34554 2569
rect 34498 2519 34500 2557
rect 34500 2519 34552 2557
rect 34552 2519 34554 2557
rect 34498 2493 34554 2495
rect 34498 2441 34500 2493
rect 34500 2441 34552 2493
rect 34552 2441 34554 2493
rect 34498 2439 34554 2441
rect 34498 2377 34500 2415
rect 34500 2377 34552 2415
rect 34552 2377 34554 2415
rect 34498 2365 34554 2377
rect 34498 2359 34500 2365
rect 34500 2359 34552 2365
rect 34552 2359 34554 2365
rect 34498 2313 34500 2335
rect 34500 2313 34552 2335
rect 34552 2313 34554 2335
rect 34498 2301 34554 2313
rect 34498 2279 34500 2301
rect 34500 2279 34552 2301
rect 34552 2279 34554 2301
rect 34498 2249 34500 2255
rect 34500 2249 34552 2255
rect 34552 2249 34554 2255
rect 34498 2237 34554 2249
rect 34498 2199 34500 2237
rect 34500 2199 34552 2237
rect 34552 2199 34554 2237
rect 34498 2173 34554 2175
rect 34498 2121 34500 2173
rect 34500 2121 34552 2173
rect 34552 2121 34554 2173
rect 34498 2119 34554 2121
rect 34498 2057 34500 2095
rect 34500 2057 34552 2095
rect 34552 2057 34554 2095
rect 34498 2045 34554 2057
rect 34498 2039 34500 2045
rect 34500 2039 34552 2045
rect 34552 2039 34554 2045
rect 34498 1993 34500 2015
rect 34500 1993 34552 2015
rect 34552 1993 34554 2015
rect 34498 1981 34554 1993
rect 34498 1959 34500 1981
rect 34500 1959 34552 1981
rect 34552 1959 34554 1981
rect 34498 1929 34500 1935
rect 34500 1929 34552 1935
rect 34552 1929 34554 1935
rect 34498 1917 34554 1929
rect 34498 1879 34500 1917
rect 34500 1879 34552 1917
rect 34552 1879 34554 1917
rect 34498 1853 34554 1855
rect 34498 1801 34500 1853
rect 34500 1801 34552 1853
rect 34552 1801 34554 1853
rect 34498 1799 34554 1801
rect 34498 1737 34500 1775
rect 34500 1737 34552 1775
rect 34552 1737 34554 1775
rect 34498 1725 34554 1737
rect 34498 1719 34500 1725
rect 34500 1719 34552 1725
rect 34552 1719 34554 1725
rect 34498 1673 34500 1695
rect 34500 1673 34552 1695
rect 34552 1673 34554 1695
rect 34498 1661 34554 1673
rect 34498 1639 34500 1661
rect 34500 1639 34552 1661
rect 34552 1639 34554 1661
rect 34498 1609 34500 1615
rect 34500 1609 34552 1615
rect 34552 1609 34554 1615
rect 34498 1597 34554 1609
rect 34498 1559 34500 1597
rect 34500 1559 34552 1597
rect 34552 1559 34554 1597
rect 34498 1533 34554 1535
rect 34498 1481 34500 1533
rect 34500 1481 34552 1533
rect 34552 1481 34554 1533
rect 34498 1479 34554 1481
rect 34498 1417 34500 1455
rect 34500 1417 34552 1455
rect 34552 1417 34554 1455
rect 34498 1405 34554 1417
rect 34498 1399 34500 1405
rect 34500 1399 34552 1405
rect 34552 1399 34554 1405
rect 34498 1353 34500 1375
rect 34500 1353 34552 1375
rect 34552 1353 34554 1375
rect 34498 1341 34554 1353
rect 34498 1319 34500 1341
rect 34500 1319 34552 1341
rect 34552 1319 34554 1341
rect 34498 1289 34500 1295
rect 34500 1289 34552 1295
rect 34552 1289 34554 1295
rect 34498 1277 34554 1289
rect 34498 1239 34500 1277
rect 34500 1239 34552 1277
rect 34552 1239 34554 1277
rect 34498 1213 34554 1215
rect 34498 1161 34500 1213
rect 34500 1161 34552 1213
rect 34552 1161 34554 1213
rect 34498 1159 34554 1161
rect 34690 3133 34746 3135
rect 34690 3081 34692 3133
rect 34692 3081 34744 3133
rect 34744 3081 34746 3133
rect 34690 3079 34746 3081
rect 34690 3017 34692 3055
rect 34692 3017 34744 3055
rect 34744 3017 34746 3055
rect 34690 3005 34746 3017
rect 34690 2999 34692 3005
rect 34692 2999 34744 3005
rect 34744 2999 34746 3005
rect 34690 2953 34692 2975
rect 34692 2953 34744 2975
rect 34744 2953 34746 2975
rect 34690 2941 34746 2953
rect 34690 2919 34692 2941
rect 34692 2919 34744 2941
rect 34744 2919 34746 2941
rect 34690 2889 34692 2895
rect 34692 2889 34744 2895
rect 34744 2889 34746 2895
rect 34690 2877 34746 2889
rect 34690 2839 34692 2877
rect 34692 2839 34744 2877
rect 34744 2839 34746 2877
rect 34690 2813 34746 2815
rect 34690 2761 34692 2813
rect 34692 2761 34744 2813
rect 34744 2761 34746 2813
rect 34690 2759 34746 2761
rect 34690 2697 34692 2735
rect 34692 2697 34744 2735
rect 34744 2697 34746 2735
rect 34690 2685 34746 2697
rect 34690 2679 34692 2685
rect 34692 2679 34744 2685
rect 34744 2679 34746 2685
rect 34690 2633 34692 2655
rect 34692 2633 34744 2655
rect 34744 2633 34746 2655
rect 34690 2621 34746 2633
rect 34690 2599 34692 2621
rect 34692 2599 34744 2621
rect 34744 2599 34746 2621
rect 34690 2569 34692 2575
rect 34692 2569 34744 2575
rect 34744 2569 34746 2575
rect 34690 2557 34746 2569
rect 34690 2519 34692 2557
rect 34692 2519 34744 2557
rect 34744 2519 34746 2557
rect 34690 2493 34746 2495
rect 34690 2441 34692 2493
rect 34692 2441 34744 2493
rect 34744 2441 34746 2493
rect 34690 2439 34746 2441
rect 34690 2377 34692 2415
rect 34692 2377 34744 2415
rect 34744 2377 34746 2415
rect 34690 2365 34746 2377
rect 34690 2359 34692 2365
rect 34692 2359 34744 2365
rect 34744 2359 34746 2365
rect 34690 2313 34692 2335
rect 34692 2313 34744 2335
rect 34744 2313 34746 2335
rect 34690 2301 34746 2313
rect 34690 2279 34692 2301
rect 34692 2279 34744 2301
rect 34744 2279 34746 2301
rect 34690 2249 34692 2255
rect 34692 2249 34744 2255
rect 34744 2249 34746 2255
rect 34690 2237 34746 2249
rect 34690 2199 34692 2237
rect 34692 2199 34744 2237
rect 34744 2199 34746 2237
rect 34690 2173 34746 2175
rect 34690 2121 34692 2173
rect 34692 2121 34744 2173
rect 34744 2121 34746 2173
rect 34690 2119 34746 2121
rect 34690 2057 34692 2095
rect 34692 2057 34744 2095
rect 34744 2057 34746 2095
rect 34690 2045 34746 2057
rect 34690 2039 34692 2045
rect 34692 2039 34744 2045
rect 34744 2039 34746 2045
rect 34690 1993 34692 2015
rect 34692 1993 34744 2015
rect 34744 1993 34746 2015
rect 34690 1981 34746 1993
rect 34690 1959 34692 1981
rect 34692 1959 34744 1981
rect 34744 1959 34746 1981
rect 34690 1929 34692 1935
rect 34692 1929 34744 1935
rect 34744 1929 34746 1935
rect 34690 1917 34746 1929
rect 34690 1879 34692 1917
rect 34692 1879 34744 1917
rect 34744 1879 34746 1917
rect 34690 1853 34746 1855
rect 34690 1801 34692 1853
rect 34692 1801 34744 1853
rect 34744 1801 34746 1853
rect 34690 1799 34746 1801
rect 34690 1737 34692 1775
rect 34692 1737 34744 1775
rect 34744 1737 34746 1775
rect 34690 1725 34746 1737
rect 34690 1719 34692 1725
rect 34692 1719 34744 1725
rect 34744 1719 34746 1725
rect 34690 1673 34692 1695
rect 34692 1673 34744 1695
rect 34744 1673 34746 1695
rect 34690 1661 34746 1673
rect 34690 1639 34692 1661
rect 34692 1639 34744 1661
rect 34744 1639 34746 1661
rect 34690 1609 34692 1615
rect 34692 1609 34744 1615
rect 34744 1609 34746 1615
rect 34690 1597 34746 1609
rect 34690 1559 34692 1597
rect 34692 1559 34744 1597
rect 34744 1559 34746 1597
rect 34690 1533 34746 1535
rect 34690 1481 34692 1533
rect 34692 1481 34744 1533
rect 34744 1481 34746 1533
rect 34690 1479 34746 1481
rect 34690 1417 34692 1455
rect 34692 1417 34744 1455
rect 34744 1417 34746 1455
rect 34690 1405 34746 1417
rect 34690 1399 34692 1405
rect 34692 1399 34744 1405
rect 34744 1399 34746 1405
rect 34690 1353 34692 1375
rect 34692 1353 34744 1375
rect 34744 1353 34746 1375
rect 34690 1341 34746 1353
rect 34690 1319 34692 1341
rect 34692 1319 34744 1341
rect 34744 1319 34746 1341
rect 34690 1289 34692 1295
rect 34692 1289 34744 1295
rect 34744 1289 34746 1295
rect 34690 1277 34746 1289
rect 34690 1239 34692 1277
rect 34692 1239 34744 1277
rect 34744 1239 34746 1277
rect 34690 1213 34746 1215
rect 34690 1161 34692 1213
rect 34692 1161 34744 1213
rect 34744 1161 34746 1213
rect 34690 1159 34746 1161
rect 34882 3133 34938 3135
rect 34882 3081 34884 3133
rect 34884 3081 34936 3133
rect 34936 3081 34938 3133
rect 34882 3079 34938 3081
rect 34882 3017 34884 3055
rect 34884 3017 34936 3055
rect 34936 3017 34938 3055
rect 34882 3005 34938 3017
rect 34882 2999 34884 3005
rect 34884 2999 34936 3005
rect 34936 2999 34938 3005
rect 34882 2953 34884 2975
rect 34884 2953 34936 2975
rect 34936 2953 34938 2975
rect 34882 2941 34938 2953
rect 34882 2919 34884 2941
rect 34884 2919 34936 2941
rect 34936 2919 34938 2941
rect 34882 2889 34884 2895
rect 34884 2889 34936 2895
rect 34936 2889 34938 2895
rect 34882 2877 34938 2889
rect 34882 2839 34884 2877
rect 34884 2839 34936 2877
rect 34936 2839 34938 2877
rect 34882 2813 34938 2815
rect 34882 2761 34884 2813
rect 34884 2761 34936 2813
rect 34936 2761 34938 2813
rect 34882 2759 34938 2761
rect 34882 2697 34884 2735
rect 34884 2697 34936 2735
rect 34936 2697 34938 2735
rect 34882 2685 34938 2697
rect 34882 2679 34884 2685
rect 34884 2679 34936 2685
rect 34936 2679 34938 2685
rect 34882 2633 34884 2655
rect 34884 2633 34936 2655
rect 34936 2633 34938 2655
rect 34882 2621 34938 2633
rect 34882 2599 34884 2621
rect 34884 2599 34936 2621
rect 34936 2599 34938 2621
rect 34882 2569 34884 2575
rect 34884 2569 34936 2575
rect 34936 2569 34938 2575
rect 34882 2557 34938 2569
rect 34882 2519 34884 2557
rect 34884 2519 34936 2557
rect 34936 2519 34938 2557
rect 34882 2493 34938 2495
rect 34882 2441 34884 2493
rect 34884 2441 34936 2493
rect 34936 2441 34938 2493
rect 34882 2439 34938 2441
rect 34882 2377 34884 2415
rect 34884 2377 34936 2415
rect 34936 2377 34938 2415
rect 34882 2365 34938 2377
rect 34882 2359 34884 2365
rect 34884 2359 34936 2365
rect 34936 2359 34938 2365
rect 34882 2313 34884 2335
rect 34884 2313 34936 2335
rect 34936 2313 34938 2335
rect 34882 2301 34938 2313
rect 34882 2279 34884 2301
rect 34884 2279 34936 2301
rect 34936 2279 34938 2301
rect 34882 2249 34884 2255
rect 34884 2249 34936 2255
rect 34936 2249 34938 2255
rect 34882 2237 34938 2249
rect 34882 2199 34884 2237
rect 34884 2199 34936 2237
rect 34936 2199 34938 2237
rect 34882 2173 34938 2175
rect 34882 2121 34884 2173
rect 34884 2121 34936 2173
rect 34936 2121 34938 2173
rect 34882 2119 34938 2121
rect 34882 2057 34884 2095
rect 34884 2057 34936 2095
rect 34936 2057 34938 2095
rect 34882 2045 34938 2057
rect 34882 2039 34884 2045
rect 34884 2039 34936 2045
rect 34936 2039 34938 2045
rect 34882 1993 34884 2015
rect 34884 1993 34936 2015
rect 34936 1993 34938 2015
rect 34882 1981 34938 1993
rect 34882 1959 34884 1981
rect 34884 1959 34936 1981
rect 34936 1959 34938 1981
rect 34882 1929 34884 1935
rect 34884 1929 34936 1935
rect 34936 1929 34938 1935
rect 34882 1917 34938 1929
rect 34882 1879 34884 1917
rect 34884 1879 34936 1917
rect 34936 1879 34938 1917
rect 34882 1853 34938 1855
rect 34882 1801 34884 1853
rect 34884 1801 34936 1853
rect 34936 1801 34938 1853
rect 34882 1799 34938 1801
rect 34882 1737 34884 1775
rect 34884 1737 34936 1775
rect 34936 1737 34938 1775
rect 34882 1725 34938 1737
rect 34882 1719 34884 1725
rect 34884 1719 34936 1725
rect 34936 1719 34938 1725
rect 34882 1673 34884 1695
rect 34884 1673 34936 1695
rect 34936 1673 34938 1695
rect 34882 1661 34938 1673
rect 34882 1639 34884 1661
rect 34884 1639 34936 1661
rect 34936 1639 34938 1661
rect 34882 1609 34884 1615
rect 34884 1609 34936 1615
rect 34936 1609 34938 1615
rect 34882 1597 34938 1609
rect 34882 1559 34884 1597
rect 34884 1559 34936 1597
rect 34936 1559 34938 1597
rect 34882 1533 34938 1535
rect 34882 1481 34884 1533
rect 34884 1481 34936 1533
rect 34936 1481 34938 1533
rect 34882 1479 34938 1481
rect 34882 1417 34884 1455
rect 34884 1417 34936 1455
rect 34936 1417 34938 1455
rect 34882 1405 34938 1417
rect 34882 1399 34884 1405
rect 34884 1399 34936 1405
rect 34936 1399 34938 1405
rect 34882 1353 34884 1375
rect 34884 1353 34936 1375
rect 34936 1353 34938 1375
rect 34882 1341 34938 1353
rect 34882 1319 34884 1341
rect 34884 1319 34936 1341
rect 34936 1319 34938 1341
rect 34882 1289 34884 1295
rect 34884 1289 34936 1295
rect 34936 1289 34938 1295
rect 34882 1277 34938 1289
rect 34882 1239 34884 1277
rect 34884 1239 34936 1277
rect 34936 1239 34938 1277
rect 34882 1213 34938 1215
rect 34882 1161 34884 1213
rect 34884 1161 34936 1213
rect 34936 1161 34938 1213
rect 34882 1159 34938 1161
rect 35074 3133 35130 3135
rect 35074 3081 35076 3133
rect 35076 3081 35128 3133
rect 35128 3081 35130 3133
rect 35074 3079 35130 3081
rect 35074 3017 35076 3055
rect 35076 3017 35128 3055
rect 35128 3017 35130 3055
rect 35074 3005 35130 3017
rect 35074 2999 35076 3005
rect 35076 2999 35128 3005
rect 35128 2999 35130 3005
rect 35074 2953 35076 2975
rect 35076 2953 35128 2975
rect 35128 2953 35130 2975
rect 35074 2941 35130 2953
rect 35074 2919 35076 2941
rect 35076 2919 35128 2941
rect 35128 2919 35130 2941
rect 35074 2889 35076 2895
rect 35076 2889 35128 2895
rect 35128 2889 35130 2895
rect 35074 2877 35130 2889
rect 35074 2839 35076 2877
rect 35076 2839 35128 2877
rect 35128 2839 35130 2877
rect 35074 2813 35130 2815
rect 35074 2761 35076 2813
rect 35076 2761 35128 2813
rect 35128 2761 35130 2813
rect 35074 2759 35130 2761
rect 35074 2697 35076 2735
rect 35076 2697 35128 2735
rect 35128 2697 35130 2735
rect 35074 2685 35130 2697
rect 35074 2679 35076 2685
rect 35076 2679 35128 2685
rect 35128 2679 35130 2685
rect 35074 2633 35076 2655
rect 35076 2633 35128 2655
rect 35128 2633 35130 2655
rect 35074 2621 35130 2633
rect 35074 2599 35076 2621
rect 35076 2599 35128 2621
rect 35128 2599 35130 2621
rect 35074 2569 35076 2575
rect 35076 2569 35128 2575
rect 35128 2569 35130 2575
rect 35074 2557 35130 2569
rect 35074 2519 35076 2557
rect 35076 2519 35128 2557
rect 35128 2519 35130 2557
rect 35074 2493 35130 2495
rect 35074 2441 35076 2493
rect 35076 2441 35128 2493
rect 35128 2441 35130 2493
rect 35074 2439 35130 2441
rect 35074 2377 35076 2415
rect 35076 2377 35128 2415
rect 35128 2377 35130 2415
rect 35074 2365 35130 2377
rect 35074 2359 35076 2365
rect 35076 2359 35128 2365
rect 35128 2359 35130 2365
rect 35074 2313 35076 2335
rect 35076 2313 35128 2335
rect 35128 2313 35130 2335
rect 35074 2301 35130 2313
rect 35074 2279 35076 2301
rect 35076 2279 35128 2301
rect 35128 2279 35130 2301
rect 35074 2249 35076 2255
rect 35076 2249 35128 2255
rect 35128 2249 35130 2255
rect 35074 2237 35130 2249
rect 35074 2199 35076 2237
rect 35076 2199 35128 2237
rect 35128 2199 35130 2237
rect 35074 2173 35130 2175
rect 35074 2121 35076 2173
rect 35076 2121 35128 2173
rect 35128 2121 35130 2173
rect 35074 2119 35130 2121
rect 35074 2057 35076 2095
rect 35076 2057 35128 2095
rect 35128 2057 35130 2095
rect 35074 2045 35130 2057
rect 35074 2039 35076 2045
rect 35076 2039 35128 2045
rect 35128 2039 35130 2045
rect 35074 1993 35076 2015
rect 35076 1993 35128 2015
rect 35128 1993 35130 2015
rect 35074 1981 35130 1993
rect 35074 1959 35076 1981
rect 35076 1959 35128 1981
rect 35128 1959 35130 1981
rect 35074 1929 35076 1935
rect 35076 1929 35128 1935
rect 35128 1929 35130 1935
rect 35074 1917 35130 1929
rect 35074 1879 35076 1917
rect 35076 1879 35128 1917
rect 35128 1879 35130 1917
rect 35074 1853 35130 1855
rect 35074 1801 35076 1853
rect 35076 1801 35128 1853
rect 35128 1801 35130 1853
rect 35074 1799 35130 1801
rect 35074 1737 35076 1775
rect 35076 1737 35128 1775
rect 35128 1737 35130 1775
rect 35074 1725 35130 1737
rect 35074 1719 35076 1725
rect 35076 1719 35128 1725
rect 35128 1719 35130 1725
rect 35074 1673 35076 1695
rect 35076 1673 35128 1695
rect 35128 1673 35130 1695
rect 35074 1661 35130 1673
rect 35074 1639 35076 1661
rect 35076 1639 35128 1661
rect 35128 1639 35130 1661
rect 35074 1609 35076 1615
rect 35076 1609 35128 1615
rect 35128 1609 35130 1615
rect 35074 1597 35130 1609
rect 35074 1559 35076 1597
rect 35076 1559 35128 1597
rect 35128 1559 35130 1597
rect 35074 1533 35130 1535
rect 35074 1481 35076 1533
rect 35076 1481 35128 1533
rect 35128 1481 35130 1533
rect 35074 1479 35130 1481
rect 35074 1417 35076 1455
rect 35076 1417 35128 1455
rect 35128 1417 35130 1455
rect 35074 1405 35130 1417
rect 35074 1399 35076 1405
rect 35076 1399 35128 1405
rect 35128 1399 35130 1405
rect 35074 1353 35076 1375
rect 35076 1353 35128 1375
rect 35128 1353 35130 1375
rect 35074 1341 35130 1353
rect 35074 1319 35076 1341
rect 35076 1319 35128 1341
rect 35128 1319 35130 1341
rect 35074 1289 35076 1295
rect 35076 1289 35128 1295
rect 35128 1289 35130 1295
rect 35074 1277 35130 1289
rect 35074 1239 35076 1277
rect 35076 1239 35128 1277
rect 35128 1239 35130 1277
rect 35074 1213 35130 1215
rect 35074 1161 35076 1213
rect 35076 1161 35128 1213
rect 35128 1161 35130 1213
rect 35074 1159 35130 1161
rect 35266 3133 35322 3135
rect 35266 3081 35268 3133
rect 35268 3081 35320 3133
rect 35320 3081 35322 3133
rect 35266 3079 35322 3081
rect 35266 3017 35268 3055
rect 35268 3017 35320 3055
rect 35320 3017 35322 3055
rect 35266 3005 35322 3017
rect 35266 2999 35268 3005
rect 35268 2999 35320 3005
rect 35320 2999 35322 3005
rect 35266 2953 35268 2975
rect 35268 2953 35320 2975
rect 35320 2953 35322 2975
rect 35266 2941 35322 2953
rect 35266 2919 35268 2941
rect 35268 2919 35320 2941
rect 35320 2919 35322 2941
rect 35266 2889 35268 2895
rect 35268 2889 35320 2895
rect 35320 2889 35322 2895
rect 35266 2877 35322 2889
rect 35266 2839 35268 2877
rect 35268 2839 35320 2877
rect 35320 2839 35322 2877
rect 35266 2813 35322 2815
rect 35266 2761 35268 2813
rect 35268 2761 35320 2813
rect 35320 2761 35322 2813
rect 35266 2759 35322 2761
rect 35266 2697 35268 2735
rect 35268 2697 35320 2735
rect 35320 2697 35322 2735
rect 35266 2685 35322 2697
rect 35266 2679 35268 2685
rect 35268 2679 35320 2685
rect 35320 2679 35322 2685
rect 35266 2633 35268 2655
rect 35268 2633 35320 2655
rect 35320 2633 35322 2655
rect 35266 2621 35322 2633
rect 35266 2599 35268 2621
rect 35268 2599 35320 2621
rect 35320 2599 35322 2621
rect 35266 2569 35268 2575
rect 35268 2569 35320 2575
rect 35320 2569 35322 2575
rect 35266 2557 35322 2569
rect 35266 2519 35268 2557
rect 35268 2519 35320 2557
rect 35320 2519 35322 2557
rect 35266 2493 35322 2495
rect 35266 2441 35268 2493
rect 35268 2441 35320 2493
rect 35320 2441 35322 2493
rect 35266 2439 35322 2441
rect 35266 2377 35268 2415
rect 35268 2377 35320 2415
rect 35320 2377 35322 2415
rect 35266 2365 35322 2377
rect 35266 2359 35268 2365
rect 35268 2359 35320 2365
rect 35320 2359 35322 2365
rect 35266 2313 35268 2335
rect 35268 2313 35320 2335
rect 35320 2313 35322 2335
rect 35266 2301 35322 2313
rect 35266 2279 35268 2301
rect 35268 2279 35320 2301
rect 35320 2279 35322 2301
rect 35266 2249 35268 2255
rect 35268 2249 35320 2255
rect 35320 2249 35322 2255
rect 35266 2237 35322 2249
rect 35266 2199 35268 2237
rect 35268 2199 35320 2237
rect 35320 2199 35322 2237
rect 35266 2173 35322 2175
rect 35266 2121 35268 2173
rect 35268 2121 35320 2173
rect 35320 2121 35322 2173
rect 35266 2119 35322 2121
rect 35266 2057 35268 2095
rect 35268 2057 35320 2095
rect 35320 2057 35322 2095
rect 35266 2045 35322 2057
rect 35266 2039 35268 2045
rect 35268 2039 35320 2045
rect 35320 2039 35322 2045
rect 35266 1993 35268 2015
rect 35268 1993 35320 2015
rect 35320 1993 35322 2015
rect 35266 1981 35322 1993
rect 35266 1959 35268 1981
rect 35268 1959 35320 1981
rect 35320 1959 35322 1981
rect 35266 1929 35268 1935
rect 35268 1929 35320 1935
rect 35320 1929 35322 1935
rect 35266 1917 35322 1929
rect 35266 1879 35268 1917
rect 35268 1879 35320 1917
rect 35320 1879 35322 1917
rect 35266 1853 35322 1855
rect 35266 1801 35268 1853
rect 35268 1801 35320 1853
rect 35320 1801 35322 1853
rect 35266 1799 35322 1801
rect 35266 1737 35268 1775
rect 35268 1737 35320 1775
rect 35320 1737 35322 1775
rect 35266 1725 35322 1737
rect 35266 1719 35268 1725
rect 35268 1719 35320 1725
rect 35320 1719 35322 1725
rect 35266 1673 35268 1695
rect 35268 1673 35320 1695
rect 35320 1673 35322 1695
rect 35266 1661 35322 1673
rect 35266 1639 35268 1661
rect 35268 1639 35320 1661
rect 35320 1639 35322 1661
rect 35266 1609 35268 1615
rect 35268 1609 35320 1615
rect 35320 1609 35322 1615
rect 35266 1597 35322 1609
rect 35266 1559 35268 1597
rect 35268 1559 35320 1597
rect 35320 1559 35322 1597
rect 35266 1533 35322 1535
rect 35266 1481 35268 1533
rect 35268 1481 35320 1533
rect 35320 1481 35322 1533
rect 35266 1479 35322 1481
rect 35266 1417 35268 1455
rect 35268 1417 35320 1455
rect 35320 1417 35322 1455
rect 35266 1405 35322 1417
rect 35266 1399 35268 1405
rect 35268 1399 35320 1405
rect 35320 1399 35322 1405
rect 35266 1353 35268 1375
rect 35268 1353 35320 1375
rect 35320 1353 35322 1375
rect 35266 1341 35322 1353
rect 35266 1319 35268 1341
rect 35268 1319 35320 1341
rect 35320 1319 35322 1341
rect 35266 1289 35268 1295
rect 35268 1289 35320 1295
rect 35320 1289 35322 1295
rect 35266 1277 35322 1289
rect 35266 1239 35268 1277
rect 35268 1239 35320 1277
rect 35320 1239 35322 1277
rect 35266 1213 35322 1215
rect 35266 1161 35268 1213
rect 35268 1161 35320 1213
rect 35320 1161 35322 1213
rect 35266 1159 35322 1161
rect 35458 3133 35514 3135
rect 35458 3081 35460 3133
rect 35460 3081 35512 3133
rect 35512 3081 35514 3133
rect 35458 3079 35514 3081
rect 35458 3017 35460 3055
rect 35460 3017 35512 3055
rect 35512 3017 35514 3055
rect 35458 3005 35514 3017
rect 35458 2999 35460 3005
rect 35460 2999 35512 3005
rect 35512 2999 35514 3005
rect 35458 2953 35460 2975
rect 35460 2953 35512 2975
rect 35512 2953 35514 2975
rect 35458 2941 35514 2953
rect 35458 2919 35460 2941
rect 35460 2919 35512 2941
rect 35512 2919 35514 2941
rect 35458 2889 35460 2895
rect 35460 2889 35512 2895
rect 35512 2889 35514 2895
rect 35458 2877 35514 2889
rect 35458 2839 35460 2877
rect 35460 2839 35512 2877
rect 35512 2839 35514 2877
rect 35458 2813 35514 2815
rect 35458 2761 35460 2813
rect 35460 2761 35512 2813
rect 35512 2761 35514 2813
rect 35458 2759 35514 2761
rect 35458 2697 35460 2735
rect 35460 2697 35512 2735
rect 35512 2697 35514 2735
rect 35458 2685 35514 2697
rect 35458 2679 35460 2685
rect 35460 2679 35512 2685
rect 35512 2679 35514 2685
rect 35458 2633 35460 2655
rect 35460 2633 35512 2655
rect 35512 2633 35514 2655
rect 35458 2621 35514 2633
rect 35458 2599 35460 2621
rect 35460 2599 35512 2621
rect 35512 2599 35514 2621
rect 35458 2569 35460 2575
rect 35460 2569 35512 2575
rect 35512 2569 35514 2575
rect 35458 2557 35514 2569
rect 35458 2519 35460 2557
rect 35460 2519 35512 2557
rect 35512 2519 35514 2557
rect 35458 2493 35514 2495
rect 35458 2441 35460 2493
rect 35460 2441 35512 2493
rect 35512 2441 35514 2493
rect 35458 2439 35514 2441
rect 35458 2377 35460 2415
rect 35460 2377 35512 2415
rect 35512 2377 35514 2415
rect 35458 2365 35514 2377
rect 35458 2359 35460 2365
rect 35460 2359 35512 2365
rect 35512 2359 35514 2365
rect 35458 2313 35460 2335
rect 35460 2313 35512 2335
rect 35512 2313 35514 2335
rect 35458 2301 35514 2313
rect 35458 2279 35460 2301
rect 35460 2279 35512 2301
rect 35512 2279 35514 2301
rect 35458 2249 35460 2255
rect 35460 2249 35512 2255
rect 35512 2249 35514 2255
rect 35458 2237 35514 2249
rect 35458 2199 35460 2237
rect 35460 2199 35512 2237
rect 35512 2199 35514 2237
rect 35458 2173 35514 2175
rect 35458 2121 35460 2173
rect 35460 2121 35512 2173
rect 35512 2121 35514 2173
rect 35458 2119 35514 2121
rect 35458 2057 35460 2095
rect 35460 2057 35512 2095
rect 35512 2057 35514 2095
rect 35458 2045 35514 2057
rect 35458 2039 35460 2045
rect 35460 2039 35512 2045
rect 35512 2039 35514 2045
rect 35458 1993 35460 2015
rect 35460 1993 35512 2015
rect 35512 1993 35514 2015
rect 35458 1981 35514 1993
rect 35458 1959 35460 1981
rect 35460 1959 35512 1981
rect 35512 1959 35514 1981
rect 35458 1929 35460 1935
rect 35460 1929 35512 1935
rect 35512 1929 35514 1935
rect 35458 1917 35514 1929
rect 35458 1879 35460 1917
rect 35460 1879 35512 1917
rect 35512 1879 35514 1917
rect 35458 1853 35514 1855
rect 35458 1801 35460 1853
rect 35460 1801 35512 1853
rect 35512 1801 35514 1853
rect 35458 1799 35514 1801
rect 35458 1737 35460 1775
rect 35460 1737 35512 1775
rect 35512 1737 35514 1775
rect 35458 1725 35514 1737
rect 35458 1719 35460 1725
rect 35460 1719 35512 1725
rect 35512 1719 35514 1725
rect 35458 1673 35460 1695
rect 35460 1673 35512 1695
rect 35512 1673 35514 1695
rect 35458 1661 35514 1673
rect 35458 1639 35460 1661
rect 35460 1639 35512 1661
rect 35512 1639 35514 1661
rect 35458 1609 35460 1615
rect 35460 1609 35512 1615
rect 35512 1609 35514 1615
rect 35458 1597 35514 1609
rect 35458 1559 35460 1597
rect 35460 1559 35512 1597
rect 35512 1559 35514 1597
rect 35458 1533 35514 1535
rect 35458 1481 35460 1533
rect 35460 1481 35512 1533
rect 35512 1481 35514 1533
rect 35458 1479 35514 1481
rect 35458 1417 35460 1455
rect 35460 1417 35512 1455
rect 35512 1417 35514 1455
rect 35458 1405 35514 1417
rect 35458 1399 35460 1405
rect 35460 1399 35512 1405
rect 35512 1399 35514 1405
rect 35458 1353 35460 1375
rect 35460 1353 35512 1375
rect 35512 1353 35514 1375
rect 35458 1341 35514 1353
rect 35458 1319 35460 1341
rect 35460 1319 35512 1341
rect 35512 1319 35514 1341
rect 35458 1289 35460 1295
rect 35460 1289 35512 1295
rect 35512 1289 35514 1295
rect 35458 1277 35514 1289
rect 35458 1239 35460 1277
rect 35460 1239 35512 1277
rect 35512 1239 35514 1277
rect 35458 1213 35514 1215
rect 35458 1161 35460 1213
rect 35460 1161 35512 1213
rect 35512 1161 35514 1213
rect 35458 1159 35514 1161
rect 35650 3133 35706 3135
rect 35650 3081 35652 3133
rect 35652 3081 35704 3133
rect 35704 3081 35706 3133
rect 35650 3079 35706 3081
rect 35650 3017 35652 3055
rect 35652 3017 35704 3055
rect 35704 3017 35706 3055
rect 35650 3005 35706 3017
rect 35650 2999 35652 3005
rect 35652 2999 35704 3005
rect 35704 2999 35706 3005
rect 35650 2953 35652 2975
rect 35652 2953 35704 2975
rect 35704 2953 35706 2975
rect 35650 2941 35706 2953
rect 35650 2919 35652 2941
rect 35652 2919 35704 2941
rect 35704 2919 35706 2941
rect 35650 2889 35652 2895
rect 35652 2889 35704 2895
rect 35704 2889 35706 2895
rect 35650 2877 35706 2889
rect 35650 2839 35652 2877
rect 35652 2839 35704 2877
rect 35704 2839 35706 2877
rect 35650 2813 35706 2815
rect 35650 2761 35652 2813
rect 35652 2761 35704 2813
rect 35704 2761 35706 2813
rect 35650 2759 35706 2761
rect 35650 2697 35652 2735
rect 35652 2697 35704 2735
rect 35704 2697 35706 2735
rect 35650 2685 35706 2697
rect 35650 2679 35652 2685
rect 35652 2679 35704 2685
rect 35704 2679 35706 2685
rect 35650 2633 35652 2655
rect 35652 2633 35704 2655
rect 35704 2633 35706 2655
rect 35650 2621 35706 2633
rect 35650 2599 35652 2621
rect 35652 2599 35704 2621
rect 35704 2599 35706 2621
rect 35650 2569 35652 2575
rect 35652 2569 35704 2575
rect 35704 2569 35706 2575
rect 35650 2557 35706 2569
rect 35650 2519 35652 2557
rect 35652 2519 35704 2557
rect 35704 2519 35706 2557
rect 35650 2493 35706 2495
rect 35650 2441 35652 2493
rect 35652 2441 35704 2493
rect 35704 2441 35706 2493
rect 35650 2439 35706 2441
rect 35650 2377 35652 2415
rect 35652 2377 35704 2415
rect 35704 2377 35706 2415
rect 35650 2365 35706 2377
rect 35650 2359 35652 2365
rect 35652 2359 35704 2365
rect 35704 2359 35706 2365
rect 35650 2313 35652 2335
rect 35652 2313 35704 2335
rect 35704 2313 35706 2335
rect 35650 2301 35706 2313
rect 35650 2279 35652 2301
rect 35652 2279 35704 2301
rect 35704 2279 35706 2301
rect 35650 2249 35652 2255
rect 35652 2249 35704 2255
rect 35704 2249 35706 2255
rect 35650 2237 35706 2249
rect 35650 2199 35652 2237
rect 35652 2199 35704 2237
rect 35704 2199 35706 2237
rect 35650 2173 35706 2175
rect 35650 2121 35652 2173
rect 35652 2121 35704 2173
rect 35704 2121 35706 2173
rect 35650 2119 35706 2121
rect 35650 2057 35652 2095
rect 35652 2057 35704 2095
rect 35704 2057 35706 2095
rect 35650 2045 35706 2057
rect 35650 2039 35652 2045
rect 35652 2039 35704 2045
rect 35704 2039 35706 2045
rect 35650 1993 35652 2015
rect 35652 1993 35704 2015
rect 35704 1993 35706 2015
rect 35650 1981 35706 1993
rect 35650 1959 35652 1981
rect 35652 1959 35704 1981
rect 35704 1959 35706 1981
rect 35650 1929 35652 1935
rect 35652 1929 35704 1935
rect 35704 1929 35706 1935
rect 35650 1917 35706 1929
rect 35650 1879 35652 1917
rect 35652 1879 35704 1917
rect 35704 1879 35706 1917
rect 35650 1853 35706 1855
rect 35650 1801 35652 1853
rect 35652 1801 35704 1853
rect 35704 1801 35706 1853
rect 35650 1799 35706 1801
rect 35650 1737 35652 1775
rect 35652 1737 35704 1775
rect 35704 1737 35706 1775
rect 35650 1725 35706 1737
rect 35650 1719 35652 1725
rect 35652 1719 35704 1725
rect 35704 1719 35706 1725
rect 35650 1673 35652 1695
rect 35652 1673 35704 1695
rect 35704 1673 35706 1695
rect 35650 1661 35706 1673
rect 35650 1639 35652 1661
rect 35652 1639 35704 1661
rect 35704 1639 35706 1661
rect 35650 1609 35652 1615
rect 35652 1609 35704 1615
rect 35704 1609 35706 1615
rect 35650 1597 35706 1609
rect 35650 1559 35652 1597
rect 35652 1559 35704 1597
rect 35704 1559 35706 1597
rect 35650 1533 35706 1535
rect 35650 1481 35652 1533
rect 35652 1481 35704 1533
rect 35704 1481 35706 1533
rect 35650 1479 35706 1481
rect 35650 1417 35652 1455
rect 35652 1417 35704 1455
rect 35704 1417 35706 1455
rect 35650 1405 35706 1417
rect 35650 1399 35652 1405
rect 35652 1399 35704 1405
rect 35704 1399 35706 1405
rect 35650 1353 35652 1375
rect 35652 1353 35704 1375
rect 35704 1353 35706 1375
rect 35650 1341 35706 1353
rect 35650 1319 35652 1341
rect 35652 1319 35704 1341
rect 35704 1319 35706 1341
rect 35650 1289 35652 1295
rect 35652 1289 35704 1295
rect 35704 1289 35706 1295
rect 35650 1277 35706 1289
rect 35650 1239 35652 1277
rect 35652 1239 35704 1277
rect 35704 1239 35706 1277
rect 35650 1213 35706 1215
rect 35650 1161 35652 1213
rect 35652 1161 35704 1213
rect 35704 1161 35706 1213
rect 35650 1159 35706 1161
rect 35842 3133 35898 3135
rect 35842 3081 35844 3133
rect 35844 3081 35896 3133
rect 35896 3081 35898 3133
rect 35842 3079 35898 3081
rect 35842 3017 35844 3055
rect 35844 3017 35896 3055
rect 35896 3017 35898 3055
rect 35842 3005 35898 3017
rect 35842 2999 35844 3005
rect 35844 2999 35896 3005
rect 35896 2999 35898 3005
rect 35842 2953 35844 2975
rect 35844 2953 35896 2975
rect 35896 2953 35898 2975
rect 35842 2941 35898 2953
rect 35842 2919 35844 2941
rect 35844 2919 35896 2941
rect 35896 2919 35898 2941
rect 35842 2889 35844 2895
rect 35844 2889 35896 2895
rect 35896 2889 35898 2895
rect 35842 2877 35898 2889
rect 35842 2839 35844 2877
rect 35844 2839 35896 2877
rect 35896 2839 35898 2877
rect 35842 2813 35898 2815
rect 35842 2761 35844 2813
rect 35844 2761 35896 2813
rect 35896 2761 35898 2813
rect 35842 2759 35898 2761
rect 35842 2697 35844 2735
rect 35844 2697 35896 2735
rect 35896 2697 35898 2735
rect 35842 2685 35898 2697
rect 35842 2679 35844 2685
rect 35844 2679 35896 2685
rect 35896 2679 35898 2685
rect 35842 2633 35844 2655
rect 35844 2633 35896 2655
rect 35896 2633 35898 2655
rect 35842 2621 35898 2633
rect 35842 2599 35844 2621
rect 35844 2599 35896 2621
rect 35896 2599 35898 2621
rect 35842 2569 35844 2575
rect 35844 2569 35896 2575
rect 35896 2569 35898 2575
rect 35842 2557 35898 2569
rect 35842 2519 35844 2557
rect 35844 2519 35896 2557
rect 35896 2519 35898 2557
rect 35842 2493 35898 2495
rect 35842 2441 35844 2493
rect 35844 2441 35896 2493
rect 35896 2441 35898 2493
rect 35842 2439 35898 2441
rect 35842 2377 35844 2415
rect 35844 2377 35896 2415
rect 35896 2377 35898 2415
rect 35842 2365 35898 2377
rect 35842 2359 35844 2365
rect 35844 2359 35896 2365
rect 35896 2359 35898 2365
rect 35842 2313 35844 2335
rect 35844 2313 35896 2335
rect 35896 2313 35898 2335
rect 35842 2301 35898 2313
rect 35842 2279 35844 2301
rect 35844 2279 35896 2301
rect 35896 2279 35898 2301
rect 35842 2249 35844 2255
rect 35844 2249 35896 2255
rect 35896 2249 35898 2255
rect 35842 2237 35898 2249
rect 35842 2199 35844 2237
rect 35844 2199 35896 2237
rect 35896 2199 35898 2237
rect 35842 2173 35898 2175
rect 35842 2121 35844 2173
rect 35844 2121 35896 2173
rect 35896 2121 35898 2173
rect 35842 2119 35898 2121
rect 35842 2057 35844 2095
rect 35844 2057 35896 2095
rect 35896 2057 35898 2095
rect 35842 2045 35898 2057
rect 35842 2039 35844 2045
rect 35844 2039 35896 2045
rect 35896 2039 35898 2045
rect 35842 1993 35844 2015
rect 35844 1993 35896 2015
rect 35896 1993 35898 2015
rect 35842 1981 35898 1993
rect 35842 1959 35844 1981
rect 35844 1959 35896 1981
rect 35896 1959 35898 1981
rect 35842 1929 35844 1935
rect 35844 1929 35896 1935
rect 35896 1929 35898 1935
rect 35842 1917 35898 1929
rect 35842 1879 35844 1917
rect 35844 1879 35896 1917
rect 35896 1879 35898 1917
rect 35842 1853 35898 1855
rect 35842 1801 35844 1853
rect 35844 1801 35896 1853
rect 35896 1801 35898 1853
rect 35842 1799 35898 1801
rect 35842 1737 35844 1775
rect 35844 1737 35896 1775
rect 35896 1737 35898 1775
rect 35842 1725 35898 1737
rect 35842 1719 35844 1725
rect 35844 1719 35896 1725
rect 35896 1719 35898 1725
rect 35842 1673 35844 1695
rect 35844 1673 35896 1695
rect 35896 1673 35898 1695
rect 35842 1661 35898 1673
rect 35842 1639 35844 1661
rect 35844 1639 35896 1661
rect 35896 1639 35898 1661
rect 35842 1609 35844 1615
rect 35844 1609 35896 1615
rect 35896 1609 35898 1615
rect 35842 1597 35898 1609
rect 35842 1559 35844 1597
rect 35844 1559 35896 1597
rect 35896 1559 35898 1597
rect 35842 1533 35898 1535
rect 35842 1481 35844 1533
rect 35844 1481 35896 1533
rect 35896 1481 35898 1533
rect 35842 1479 35898 1481
rect 35842 1417 35844 1455
rect 35844 1417 35896 1455
rect 35896 1417 35898 1455
rect 35842 1405 35898 1417
rect 35842 1399 35844 1405
rect 35844 1399 35896 1405
rect 35896 1399 35898 1405
rect 35842 1353 35844 1375
rect 35844 1353 35896 1375
rect 35896 1353 35898 1375
rect 35842 1341 35898 1353
rect 35842 1319 35844 1341
rect 35844 1319 35896 1341
rect 35896 1319 35898 1341
rect 35842 1289 35844 1295
rect 35844 1289 35896 1295
rect 35896 1289 35898 1295
rect 35842 1277 35898 1289
rect 35842 1239 35844 1277
rect 35844 1239 35896 1277
rect 35896 1239 35898 1277
rect 35842 1213 35898 1215
rect 35842 1161 35844 1213
rect 35844 1161 35896 1213
rect 35896 1161 35898 1213
rect 35842 1159 35898 1161
rect 36034 3133 36090 3135
rect 36034 3081 36036 3133
rect 36036 3081 36088 3133
rect 36088 3081 36090 3133
rect 36034 3079 36090 3081
rect 36034 3017 36036 3055
rect 36036 3017 36088 3055
rect 36088 3017 36090 3055
rect 36034 3005 36090 3017
rect 36034 2999 36036 3005
rect 36036 2999 36088 3005
rect 36088 2999 36090 3005
rect 36034 2953 36036 2975
rect 36036 2953 36088 2975
rect 36088 2953 36090 2975
rect 36034 2941 36090 2953
rect 36034 2919 36036 2941
rect 36036 2919 36088 2941
rect 36088 2919 36090 2941
rect 36034 2889 36036 2895
rect 36036 2889 36088 2895
rect 36088 2889 36090 2895
rect 36034 2877 36090 2889
rect 36034 2839 36036 2877
rect 36036 2839 36088 2877
rect 36088 2839 36090 2877
rect 36034 2813 36090 2815
rect 36034 2761 36036 2813
rect 36036 2761 36088 2813
rect 36088 2761 36090 2813
rect 36034 2759 36090 2761
rect 36034 2697 36036 2735
rect 36036 2697 36088 2735
rect 36088 2697 36090 2735
rect 36034 2685 36090 2697
rect 36034 2679 36036 2685
rect 36036 2679 36088 2685
rect 36088 2679 36090 2685
rect 36034 2633 36036 2655
rect 36036 2633 36088 2655
rect 36088 2633 36090 2655
rect 36034 2621 36090 2633
rect 36034 2599 36036 2621
rect 36036 2599 36088 2621
rect 36088 2599 36090 2621
rect 36034 2569 36036 2575
rect 36036 2569 36088 2575
rect 36088 2569 36090 2575
rect 36034 2557 36090 2569
rect 36034 2519 36036 2557
rect 36036 2519 36088 2557
rect 36088 2519 36090 2557
rect 36034 2493 36090 2495
rect 36034 2441 36036 2493
rect 36036 2441 36088 2493
rect 36088 2441 36090 2493
rect 36034 2439 36090 2441
rect 36034 2377 36036 2415
rect 36036 2377 36088 2415
rect 36088 2377 36090 2415
rect 36034 2365 36090 2377
rect 36034 2359 36036 2365
rect 36036 2359 36088 2365
rect 36088 2359 36090 2365
rect 36034 2313 36036 2335
rect 36036 2313 36088 2335
rect 36088 2313 36090 2335
rect 36034 2301 36090 2313
rect 36034 2279 36036 2301
rect 36036 2279 36088 2301
rect 36088 2279 36090 2301
rect 36034 2249 36036 2255
rect 36036 2249 36088 2255
rect 36088 2249 36090 2255
rect 36034 2237 36090 2249
rect 36034 2199 36036 2237
rect 36036 2199 36088 2237
rect 36088 2199 36090 2237
rect 36034 2173 36090 2175
rect 36034 2121 36036 2173
rect 36036 2121 36088 2173
rect 36088 2121 36090 2173
rect 36034 2119 36090 2121
rect 36034 2057 36036 2095
rect 36036 2057 36088 2095
rect 36088 2057 36090 2095
rect 36034 2045 36090 2057
rect 36034 2039 36036 2045
rect 36036 2039 36088 2045
rect 36088 2039 36090 2045
rect 36034 1993 36036 2015
rect 36036 1993 36088 2015
rect 36088 1993 36090 2015
rect 36034 1981 36090 1993
rect 36034 1959 36036 1981
rect 36036 1959 36088 1981
rect 36088 1959 36090 1981
rect 36034 1929 36036 1935
rect 36036 1929 36088 1935
rect 36088 1929 36090 1935
rect 36034 1917 36090 1929
rect 36034 1879 36036 1917
rect 36036 1879 36088 1917
rect 36088 1879 36090 1917
rect 36034 1853 36090 1855
rect 36034 1801 36036 1853
rect 36036 1801 36088 1853
rect 36088 1801 36090 1853
rect 36034 1799 36090 1801
rect 36034 1737 36036 1775
rect 36036 1737 36088 1775
rect 36088 1737 36090 1775
rect 36034 1725 36090 1737
rect 36034 1719 36036 1725
rect 36036 1719 36088 1725
rect 36088 1719 36090 1725
rect 36034 1673 36036 1695
rect 36036 1673 36088 1695
rect 36088 1673 36090 1695
rect 36034 1661 36090 1673
rect 36034 1639 36036 1661
rect 36036 1639 36088 1661
rect 36088 1639 36090 1661
rect 36034 1609 36036 1615
rect 36036 1609 36088 1615
rect 36088 1609 36090 1615
rect 36034 1597 36090 1609
rect 36034 1559 36036 1597
rect 36036 1559 36088 1597
rect 36088 1559 36090 1597
rect 36034 1533 36090 1535
rect 36034 1481 36036 1533
rect 36036 1481 36088 1533
rect 36088 1481 36090 1533
rect 36034 1479 36090 1481
rect 36034 1417 36036 1455
rect 36036 1417 36088 1455
rect 36088 1417 36090 1455
rect 36034 1405 36090 1417
rect 36034 1399 36036 1405
rect 36036 1399 36088 1405
rect 36088 1399 36090 1405
rect 36034 1353 36036 1375
rect 36036 1353 36088 1375
rect 36088 1353 36090 1375
rect 36034 1341 36090 1353
rect 36034 1319 36036 1341
rect 36036 1319 36088 1341
rect 36088 1319 36090 1341
rect 36034 1289 36036 1295
rect 36036 1289 36088 1295
rect 36088 1289 36090 1295
rect 36034 1277 36090 1289
rect 36034 1239 36036 1277
rect 36036 1239 36088 1277
rect 36088 1239 36090 1277
rect 36034 1213 36090 1215
rect 36034 1161 36036 1213
rect 36036 1161 36088 1213
rect 36088 1161 36090 1213
rect 36034 1159 36090 1161
rect 36226 3133 36282 3135
rect 36226 3081 36228 3133
rect 36228 3081 36280 3133
rect 36280 3081 36282 3133
rect 36226 3079 36282 3081
rect 36226 3017 36228 3055
rect 36228 3017 36280 3055
rect 36280 3017 36282 3055
rect 36226 3005 36282 3017
rect 36226 2999 36228 3005
rect 36228 2999 36280 3005
rect 36280 2999 36282 3005
rect 36226 2953 36228 2975
rect 36228 2953 36280 2975
rect 36280 2953 36282 2975
rect 36226 2941 36282 2953
rect 36226 2919 36228 2941
rect 36228 2919 36280 2941
rect 36280 2919 36282 2941
rect 36226 2889 36228 2895
rect 36228 2889 36280 2895
rect 36280 2889 36282 2895
rect 36226 2877 36282 2889
rect 36226 2839 36228 2877
rect 36228 2839 36280 2877
rect 36280 2839 36282 2877
rect 36226 2813 36282 2815
rect 36226 2761 36228 2813
rect 36228 2761 36280 2813
rect 36280 2761 36282 2813
rect 36226 2759 36282 2761
rect 36226 2697 36228 2735
rect 36228 2697 36280 2735
rect 36280 2697 36282 2735
rect 36226 2685 36282 2697
rect 36226 2679 36228 2685
rect 36228 2679 36280 2685
rect 36280 2679 36282 2685
rect 36226 2633 36228 2655
rect 36228 2633 36280 2655
rect 36280 2633 36282 2655
rect 36226 2621 36282 2633
rect 36226 2599 36228 2621
rect 36228 2599 36280 2621
rect 36280 2599 36282 2621
rect 36226 2569 36228 2575
rect 36228 2569 36280 2575
rect 36280 2569 36282 2575
rect 36226 2557 36282 2569
rect 36226 2519 36228 2557
rect 36228 2519 36280 2557
rect 36280 2519 36282 2557
rect 36226 2493 36282 2495
rect 36226 2441 36228 2493
rect 36228 2441 36280 2493
rect 36280 2441 36282 2493
rect 36226 2439 36282 2441
rect 36226 2377 36228 2415
rect 36228 2377 36280 2415
rect 36280 2377 36282 2415
rect 36226 2365 36282 2377
rect 36226 2359 36228 2365
rect 36228 2359 36280 2365
rect 36280 2359 36282 2365
rect 36226 2313 36228 2335
rect 36228 2313 36280 2335
rect 36280 2313 36282 2335
rect 36226 2301 36282 2313
rect 36226 2279 36228 2301
rect 36228 2279 36280 2301
rect 36280 2279 36282 2301
rect 36226 2249 36228 2255
rect 36228 2249 36280 2255
rect 36280 2249 36282 2255
rect 36226 2237 36282 2249
rect 36226 2199 36228 2237
rect 36228 2199 36280 2237
rect 36280 2199 36282 2237
rect 36226 2173 36282 2175
rect 36226 2121 36228 2173
rect 36228 2121 36280 2173
rect 36280 2121 36282 2173
rect 36226 2119 36282 2121
rect 36226 2057 36228 2095
rect 36228 2057 36280 2095
rect 36280 2057 36282 2095
rect 36226 2045 36282 2057
rect 36226 2039 36228 2045
rect 36228 2039 36280 2045
rect 36280 2039 36282 2045
rect 36226 1993 36228 2015
rect 36228 1993 36280 2015
rect 36280 1993 36282 2015
rect 36226 1981 36282 1993
rect 36226 1959 36228 1981
rect 36228 1959 36280 1981
rect 36280 1959 36282 1981
rect 36226 1929 36228 1935
rect 36228 1929 36280 1935
rect 36280 1929 36282 1935
rect 36226 1917 36282 1929
rect 36226 1879 36228 1917
rect 36228 1879 36280 1917
rect 36280 1879 36282 1917
rect 36226 1853 36282 1855
rect 36226 1801 36228 1853
rect 36228 1801 36280 1853
rect 36280 1801 36282 1853
rect 36226 1799 36282 1801
rect 36226 1737 36228 1775
rect 36228 1737 36280 1775
rect 36280 1737 36282 1775
rect 36226 1725 36282 1737
rect 36226 1719 36228 1725
rect 36228 1719 36280 1725
rect 36280 1719 36282 1725
rect 36226 1673 36228 1695
rect 36228 1673 36280 1695
rect 36280 1673 36282 1695
rect 36226 1661 36282 1673
rect 36226 1639 36228 1661
rect 36228 1639 36280 1661
rect 36280 1639 36282 1661
rect 36226 1609 36228 1615
rect 36228 1609 36280 1615
rect 36280 1609 36282 1615
rect 36226 1597 36282 1609
rect 36226 1559 36228 1597
rect 36228 1559 36280 1597
rect 36280 1559 36282 1597
rect 36226 1533 36282 1535
rect 36226 1481 36228 1533
rect 36228 1481 36280 1533
rect 36280 1481 36282 1533
rect 36226 1479 36282 1481
rect 36226 1417 36228 1455
rect 36228 1417 36280 1455
rect 36280 1417 36282 1455
rect 36226 1405 36282 1417
rect 36226 1399 36228 1405
rect 36228 1399 36280 1405
rect 36280 1399 36282 1405
rect 36226 1353 36228 1375
rect 36228 1353 36280 1375
rect 36280 1353 36282 1375
rect 36226 1341 36282 1353
rect 36226 1319 36228 1341
rect 36228 1319 36280 1341
rect 36280 1319 36282 1341
rect 36226 1289 36228 1295
rect 36228 1289 36280 1295
rect 36280 1289 36282 1295
rect 36226 1277 36282 1289
rect 36226 1239 36228 1277
rect 36228 1239 36280 1277
rect 36280 1239 36282 1277
rect 36226 1213 36282 1215
rect 36226 1161 36228 1213
rect 36228 1161 36280 1213
rect 36280 1161 36282 1213
rect 36226 1159 36282 1161
rect 36418 3133 36474 3135
rect 36418 3081 36420 3133
rect 36420 3081 36472 3133
rect 36472 3081 36474 3133
rect 36418 3079 36474 3081
rect 36418 3017 36420 3055
rect 36420 3017 36472 3055
rect 36472 3017 36474 3055
rect 36418 3005 36474 3017
rect 36418 2999 36420 3005
rect 36420 2999 36472 3005
rect 36472 2999 36474 3005
rect 36418 2953 36420 2975
rect 36420 2953 36472 2975
rect 36472 2953 36474 2975
rect 36418 2941 36474 2953
rect 36418 2919 36420 2941
rect 36420 2919 36472 2941
rect 36472 2919 36474 2941
rect 36418 2889 36420 2895
rect 36420 2889 36472 2895
rect 36472 2889 36474 2895
rect 36418 2877 36474 2889
rect 36418 2839 36420 2877
rect 36420 2839 36472 2877
rect 36472 2839 36474 2877
rect 36418 2813 36474 2815
rect 36418 2761 36420 2813
rect 36420 2761 36472 2813
rect 36472 2761 36474 2813
rect 36418 2759 36474 2761
rect 36418 2697 36420 2735
rect 36420 2697 36472 2735
rect 36472 2697 36474 2735
rect 36418 2685 36474 2697
rect 36418 2679 36420 2685
rect 36420 2679 36472 2685
rect 36472 2679 36474 2685
rect 36418 2633 36420 2655
rect 36420 2633 36472 2655
rect 36472 2633 36474 2655
rect 36418 2621 36474 2633
rect 36418 2599 36420 2621
rect 36420 2599 36472 2621
rect 36472 2599 36474 2621
rect 36418 2569 36420 2575
rect 36420 2569 36472 2575
rect 36472 2569 36474 2575
rect 36418 2557 36474 2569
rect 36418 2519 36420 2557
rect 36420 2519 36472 2557
rect 36472 2519 36474 2557
rect 36418 2493 36474 2495
rect 36418 2441 36420 2493
rect 36420 2441 36472 2493
rect 36472 2441 36474 2493
rect 36418 2439 36474 2441
rect 36418 2377 36420 2415
rect 36420 2377 36472 2415
rect 36472 2377 36474 2415
rect 36418 2365 36474 2377
rect 36418 2359 36420 2365
rect 36420 2359 36472 2365
rect 36472 2359 36474 2365
rect 36418 2313 36420 2335
rect 36420 2313 36472 2335
rect 36472 2313 36474 2335
rect 36418 2301 36474 2313
rect 36418 2279 36420 2301
rect 36420 2279 36472 2301
rect 36472 2279 36474 2301
rect 36418 2249 36420 2255
rect 36420 2249 36472 2255
rect 36472 2249 36474 2255
rect 36418 2237 36474 2249
rect 36418 2199 36420 2237
rect 36420 2199 36472 2237
rect 36472 2199 36474 2237
rect 36418 2173 36474 2175
rect 36418 2121 36420 2173
rect 36420 2121 36472 2173
rect 36472 2121 36474 2173
rect 36418 2119 36474 2121
rect 36418 2057 36420 2095
rect 36420 2057 36472 2095
rect 36472 2057 36474 2095
rect 36418 2045 36474 2057
rect 36418 2039 36420 2045
rect 36420 2039 36472 2045
rect 36472 2039 36474 2045
rect 36418 1993 36420 2015
rect 36420 1993 36472 2015
rect 36472 1993 36474 2015
rect 36418 1981 36474 1993
rect 36418 1959 36420 1981
rect 36420 1959 36472 1981
rect 36472 1959 36474 1981
rect 36418 1929 36420 1935
rect 36420 1929 36472 1935
rect 36472 1929 36474 1935
rect 36418 1917 36474 1929
rect 36418 1879 36420 1917
rect 36420 1879 36472 1917
rect 36472 1879 36474 1917
rect 36418 1853 36474 1855
rect 36418 1801 36420 1853
rect 36420 1801 36472 1853
rect 36472 1801 36474 1853
rect 36418 1799 36474 1801
rect 36418 1737 36420 1775
rect 36420 1737 36472 1775
rect 36472 1737 36474 1775
rect 36418 1725 36474 1737
rect 36418 1719 36420 1725
rect 36420 1719 36472 1725
rect 36472 1719 36474 1725
rect 36418 1673 36420 1695
rect 36420 1673 36472 1695
rect 36472 1673 36474 1695
rect 36418 1661 36474 1673
rect 36418 1639 36420 1661
rect 36420 1639 36472 1661
rect 36472 1639 36474 1661
rect 36418 1609 36420 1615
rect 36420 1609 36472 1615
rect 36472 1609 36474 1615
rect 36418 1597 36474 1609
rect 36418 1559 36420 1597
rect 36420 1559 36472 1597
rect 36472 1559 36474 1597
rect 36418 1533 36474 1535
rect 36418 1481 36420 1533
rect 36420 1481 36472 1533
rect 36472 1481 36474 1533
rect 36418 1479 36474 1481
rect 36418 1417 36420 1455
rect 36420 1417 36472 1455
rect 36472 1417 36474 1455
rect 36418 1405 36474 1417
rect 36418 1399 36420 1405
rect 36420 1399 36472 1405
rect 36472 1399 36474 1405
rect 36418 1353 36420 1375
rect 36420 1353 36472 1375
rect 36472 1353 36474 1375
rect 36418 1341 36474 1353
rect 36418 1319 36420 1341
rect 36420 1319 36472 1341
rect 36472 1319 36474 1341
rect 36418 1289 36420 1295
rect 36420 1289 36472 1295
rect 36472 1289 36474 1295
rect 36418 1277 36474 1289
rect 36418 1239 36420 1277
rect 36420 1239 36472 1277
rect 36472 1239 36474 1277
rect 36418 1213 36474 1215
rect 36418 1161 36420 1213
rect 36420 1161 36472 1213
rect 36472 1161 36474 1213
rect 36418 1159 36474 1161
rect 36610 3133 36666 3135
rect 36610 3081 36612 3133
rect 36612 3081 36664 3133
rect 36664 3081 36666 3133
rect 36610 3079 36666 3081
rect 36610 3017 36612 3055
rect 36612 3017 36664 3055
rect 36664 3017 36666 3055
rect 36610 3005 36666 3017
rect 36610 2999 36612 3005
rect 36612 2999 36664 3005
rect 36664 2999 36666 3005
rect 36610 2953 36612 2975
rect 36612 2953 36664 2975
rect 36664 2953 36666 2975
rect 36610 2941 36666 2953
rect 36610 2919 36612 2941
rect 36612 2919 36664 2941
rect 36664 2919 36666 2941
rect 36610 2889 36612 2895
rect 36612 2889 36664 2895
rect 36664 2889 36666 2895
rect 36610 2877 36666 2889
rect 36610 2839 36612 2877
rect 36612 2839 36664 2877
rect 36664 2839 36666 2877
rect 36610 2813 36666 2815
rect 36610 2761 36612 2813
rect 36612 2761 36664 2813
rect 36664 2761 36666 2813
rect 36610 2759 36666 2761
rect 36610 2697 36612 2735
rect 36612 2697 36664 2735
rect 36664 2697 36666 2735
rect 36610 2685 36666 2697
rect 36610 2679 36612 2685
rect 36612 2679 36664 2685
rect 36664 2679 36666 2685
rect 36610 2633 36612 2655
rect 36612 2633 36664 2655
rect 36664 2633 36666 2655
rect 36610 2621 36666 2633
rect 36610 2599 36612 2621
rect 36612 2599 36664 2621
rect 36664 2599 36666 2621
rect 36610 2569 36612 2575
rect 36612 2569 36664 2575
rect 36664 2569 36666 2575
rect 36610 2557 36666 2569
rect 36610 2519 36612 2557
rect 36612 2519 36664 2557
rect 36664 2519 36666 2557
rect 36610 2493 36666 2495
rect 36610 2441 36612 2493
rect 36612 2441 36664 2493
rect 36664 2441 36666 2493
rect 36610 2439 36666 2441
rect 36610 2377 36612 2415
rect 36612 2377 36664 2415
rect 36664 2377 36666 2415
rect 36610 2365 36666 2377
rect 36610 2359 36612 2365
rect 36612 2359 36664 2365
rect 36664 2359 36666 2365
rect 36610 2313 36612 2335
rect 36612 2313 36664 2335
rect 36664 2313 36666 2335
rect 36610 2301 36666 2313
rect 36610 2279 36612 2301
rect 36612 2279 36664 2301
rect 36664 2279 36666 2301
rect 36610 2249 36612 2255
rect 36612 2249 36664 2255
rect 36664 2249 36666 2255
rect 36610 2237 36666 2249
rect 36610 2199 36612 2237
rect 36612 2199 36664 2237
rect 36664 2199 36666 2237
rect 36610 2173 36666 2175
rect 36610 2121 36612 2173
rect 36612 2121 36664 2173
rect 36664 2121 36666 2173
rect 36610 2119 36666 2121
rect 36610 2057 36612 2095
rect 36612 2057 36664 2095
rect 36664 2057 36666 2095
rect 36610 2045 36666 2057
rect 36610 2039 36612 2045
rect 36612 2039 36664 2045
rect 36664 2039 36666 2045
rect 36610 1993 36612 2015
rect 36612 1993 36664 2015
rect 36664 1993 36666 2015
rect 36610 1981 36666 1993
rect 36610 1959 36612 1981
rect 36612 1959 36664 1981
rect 36664 1959 36666 1981
rect 36610 1929 36612 1935
rect 36612 1929 36664 1935
rect 36664 1929 36666 1935
rect 36610 1917 36666 1929
rect 36610 1879 36612 1917
rect 36612 1879 36664 1917
rect 36664 1879 36666 1917
rect 36610 1853 36666 1855
rect 36610 1801 36612 1853
rect 36612 1801 36664 1853
rect 36664 1801 36666 1853
rect 36610 1799 36666 1801
rect 36610 1737 36612 1775
rect 36612 1737 36664 1775
rect 36664 1737 36666 1775
rect 36610 1725 36666 1737
rect 36610 1719 36612 1725
rect 36612 1719 36664 1725
rect 36664 1719 36666 1725
rect 36610 1673 36612 1695
rect 36612 1673 36664 1695
rect 36664 1673 36666 1695
rect 36610 1661 36666 1673
rect 36610 1639 36612 1661
rect 36612 1639 36664 1661
rect 36664 1639 36666 1661
rect 36610 1609 36612 1615
rect 36612 1609 36664 1615
rect 36664 1609 36666 1615
rect 36610 1597 36666 1609
rect 36610 1559 36612 1597
rect 36612 1559 36664 1597
rect 36664 1559 36666 1597
rect 36610 1533 36666 1535
rect 36610 1481 36612 1533
rect 36612 1481 36664 1533
rect 36664 1481 36666 1533
rect 36610 1479 36666 1481
rect 36610 1417 36612 1455
rect 36612 1417 36664 1455
rect 36664 1417 36666 1455
rect 36610 1405 36666 1417
rect 36610 1399 36612 1405
rect 36612 1399 36664 1405
rect 36664 1399 36666 1405
rect 36610 1353 36612 1375
rect 36612 1353 36664 1375
rect 36664 1353 36666 1375
rect 36610 1341 36666 1353
rect 36610 1319 36612 1341
rect 36612 1319 36664 1341
rect 36664 1319 36666 1341
rect 36610 1289 36612 1295
rect 36612 1289 36664 1295
rect 36664 1289 36666 1295
rect 36610 1277 36666 1289
rect 36610 1239 36612 1277
rect 36612 1239 36664 1277
rect 36664 1239 36666 1277
rect 36610 1213 36666 1215
rect 36610 1161 36612 1213
rect 36612 1161 36664 1213
rect 36664 1161 36666 1213
rect 36610 1159 36666 1161
rect 36802 3133 36858 3135
rect 36802 3081 36804 3133
rect 36804 3081 36856 3133
rect 36856 3081 36858 3133
rect 36802 3079 36858 3081
rect 36802 3017 36804 3055
rect 36804 3017 36856 3055
rect 36856 3017 36858 3055
rect 36802 3005 36858 3017
rect 36802 2999 36804 3005
rect 36804 2999 36856 3005
rect 36856 2999 36858 3005
rect 36802 2953 36804 2975
rect 36804 2953 36856 2975
rect 36856 2953 36858 2975
rect 36802 2941 36858 2953
rect 36802 2919 36804 2941
rect 36804 2919 36856 2941
rect 36856 2919 36858 2941
rect 36802 2889 36804 2895
rect 36804 2889 36856 2895
rect 36856 2889 36858 2895
rect 36802 2877 36858 2889
rect 36802 2839 36804 2877
rect 36804 2839 36856 2877
rect 36856 2839 36858 2877
rect 36802 2813 36858 2815
rect 36802 2761 36804 2813
rect 36804 2761 36856 2813
rect 36856 2761 36858 2813
rect 36802 2759 36858 2761
rect 36802 2697 36804 2735
rect 36804 2697 36856 2735
rect 36856 2697 36858 2735
rect 36802 2685 36858 2697
rect 36802 2679 36804 2685
rect 36804 2679 36856 2685
rect 36856 2679 36858 2685
rect 36802 2633 36804 2655
rect 36804 2633 36856 2655
rect 36856 2633 36858 2655
rect 36802 2621 36858 2633
rect 36802 2599 36804 2621
rect 36804 2599 36856 2621
rect 36856 2599 36858 2621
rect 36802 2569 36804 2575
rect 36804 2569 36856 2575
rect 36856 2569 36858 2575
rect 36802 2557 36858 2569
rect 36802 2519 36804 2557
rect 36804 2519 36856 2557
rect 36856 2519 36858 2557
rect 36802 2493 36858 2495
rect 36802 2441 36804 2493
rect 36804 2441 36856 2493
rect 36856 2441 36858 2493
rect 36802 2439 36858 2441
rect 36802 2377 36804 2415
rect 36804 2377 36856 2415
rect 36856 2377 36858 2415
rect 36802 2365 36858 2377
rect 36802 2359 36804 2365
rect 36804 2359 36856 2365
rect 36856 2359 36858 2365
rect 36802 2313 36804 2335
rect 36804 2313 36856 2335
rect 36856 2313 36858 2335
rect 36802 2301 36858 2313
rect 36802 2279 36804 2301
rect 36804 2279 36856 2301
rect 36856 2279 36858 2301
rect 36802 2249 36804 2255
rect 36804 2249 36856 2255
rect 36856 2249 36858 2255
rect 36802 2237 36858 2249
rect 36802 2199 36804 2237
rect 36804 2199 36856 2237
rect 36856 2199 36858 2237
rect 36802 2173 36858 2175
rect 36802 2121 36804 2173
rect 36804 2121 36856 2173
rect 36856 2121 36858 2173
rect 36802 2119 36858 2121
rect 36802 2057 36804 2095
rect 36804 2057 36856 2095
rect 36856 2057 36858 2095
rect 36802 2045 36858 2057
rect 36802 2039 36804 2045
rect 36804 2039 36856 2045
rect 36856 2039 36858 2045
rect 36802 1993 36804 2015
rect 36804 1993 36856 2015
rect 36856 1993 36858 2015
rect 36802 1981 36858 1993
rect 36802 1959 36804 1981
rect 36804 1959 36856 1981
rect 36856 1959 36858 1981
rect 36802 1929 36804 1935
rect 36804 1929 36856 1935
rect 36856 1929 36858 1935
rect 36802 1917 36858 1929
rect 36802 1879 36804 1917
rect 36804 1879 36856 1917
rect 36856 1879 36858 1917
rect 36802 1853 36858 1855
rect 36802 1801 36804 1853
rect 36804 1801 36856 1853
rect 36856 1801 36858 1853
rect 36802 1799 36858 1801
rect 36802 1737 36804 1775
rect 36804 1737 36856 1775
rect 36856 1737 36858 1775
rect 36802 1725 36858 1737
rect 36802 1719 36804 1725
rect 36804 1719 36856 1725
rect 36856 1719 36858 1725
rect 36802 1673 36804 1695
rect 36804 1673 36856 1695
rect 36856 1673 36858 1695
rect 36802 1661 36858 1673
rect 36802 1639 36804 1661
rect 36804 1639 36856 1661
rect 36856 1639 36858 1661
rect 36802 1609 36804 1615
rect 36804 1609 36856 1615
rect 36856 1609 36858 1615
rect 36802 1597 36858 1609
rect 36802 1559 36804 1597
rect 36804 1559 36856 1597
rect 36856 1559 36858 1597
rect 36802 1533 36858 1535
rect 36802 1481 36804 1533
rect 36804 1481 36856 1533
rect 36856 1481 36858 1533
rect 36802 1479 36858 1481
rect 36802 1417 36804 1455
rect 36804 1417 36856 1455
rect 36856 1417 36858 1455
rect 36802 1405 36858 1417
rect 36802 1399 36804 1405
rect 36804 1399 36856 1405
rect 36856 1399 36858 1405
rect 36802 1353 36804 1375
rect 36804 1353 36856 1375
rect 36856 1353 36858 1375
rect 36802 1341 36858 1353
rect 36802 1319 36804 1341
rect 36804 1319 36856 1341
rect 36856 1319 36858 1341
rect 36802 1289 36804 1295
rect 36804 1289 36856 1295
rect 36856 1289 36858 1295
rect 36802 1277 36858 1289
rect 36802 1239 36804 1277
rect 36804 1239 36856 1277
rect 36856 1239 36858 1277
rect 36802 1213 36858 1215
rect 36802 1161 36804 1213
rect 36804 1161 36856 1213
rect 36856 1161 36858 1213
rect 36802 1159 36858 1161
rect 36994 3133 37050 3135
rect 36994 3081 36996 3133
rect 36996 3081 37048 3133
rect 37048 3081 37050 3133
rect 36994 3079 37050 3081
rect 36994 3017 36996 3055
rect 36996 3017 37048 3055
rect 37048 3017 37050 3055
rect 36994 3005 37050 3017
rect 36994 2999 36996 3005
rect 36996 2999 37048 3005
rect 37048 2999 37050 3005
rect 36994 2953 36996 2975
rect 36996 2953 37048 2975
rect 37048 2953 37050 2975
rect 36994 2941 37050 2953
rect 36994 2919 36996 2941
rect 36996 2919 37048 2941
rect 37048 2919 37050 2941
rect 36994 2889 36996 2895
rect 36996 2889 37048 2895
rect 37048 2889 37050 2895
rect 36994 2877 37050 2889
rect 36994 2839 36996 2877
rect 36996 2839 37048 2877
rect 37048 2839 37050 2877
rect 36994 2813 37050 2815
rect 36994 2761 36996 2813
rect 36996 2761 37048 2813
rect 37048 2761 37050 2813
rect 36994 2759 37050 2761
rect 36994 2697 36996 2735
rect 36996 2697 37048 2735
rect 37048 2697 37050 2735
rect 36994 2685 37050 2697
rect 36994 2679 36996 2685
rect 36996 2679 37048 2685
rect 37048 2679 37050 2685
rect 36994 2633 36996 2655
rect 36996 2633 37048 2655
rect 37048 2633 37050 2655
rect 36994 2621 37050 2633
rect 36994 2599 36996 2621
rect 36996 2599 37048 2621
rect 37048 2599 37050 2621
rect 36994 2569 36996 2575
rect 36996 2569 37048 2575
rect 37048 2569 37050 2575
rect 36994 2557 37050 2569
rect 36994 2519 36996 2557
rect 36996 2519 37048 2557
rect 37048 2519 37050 2557
rect 36994 2493 37050 2495
rect 36994 2441 36996 2493
rect 36996 2441 37048 2493
rect 37048 2441 37050 2493
rect 36994 2439 37050 2441
rect 36994 2377 36996 2415
rect 36996 2377 37048 2415
rect 37048 2377 37050 2415
rect 36994 2365 37050 2377
rect 36994 2359 36996 2365
rect 36996 2359 37048 2365
rect 37048 2359 37050 2365
rect 36994 2313 36996 2335
rect 36996 2313 37048 2335
rect 37048 2313 37050 2335
rect 36994 2301 37050 2313
rect 36994 2279 36996 2301
rect 36996 2279 37048 2301
rect 37048 2279 37050 2301
rect 36994 2249 36996 2255
rect 36996 2249 37048 2255
rect 37048 2249 37050 2255
rect 36994 2237 37050 2249
rect 36994 2199 36996 2237
rect 36996 2199 37048 2237
rect 37048 2199 37050 2237
rect 36994 2173 37050 2175
rect 36994 2121 36996 2173
rect 36996 2121 37048 2173
rect 37048 2121 37050 2173
rect 36994 2119 37050 2121
rect 36994 2057 36996 2095
rect 36996 2057 37048 2095
rect 37048 2057 37050 2095
rect 36994 2045 37050 2057
rect 36994 2039 36996 2045
rect 36996 2039 37048 2045
rect 37048 2039 37050 2045
rect 36994 1993 36996 2015
rect 36996 1993 37048 2015
rect 37048 1993 37050 2015
rect 36994 1981 37050 1993
rect 36994 1959 36996 1981
rect 36996 1959 37048 1981
rect 37048 1959 37050 1981
rect 36994 1929 36996 1935
rect 36996 1929 37048 1935
rect 37048 1929 37050 1935
rect 36994 1917 37050 1929
rect 36994 1879 36996 1917
rect 36996 1879 37048 1917
rect 37048 1879 37050 1917
rect 36994 1853 37050 1855
rect 36994 1801 36996 1853
rect 36996 1801 37048 1853
rect 37048 1801 37050 1853
rect 36994 1799 37050 1801
rect 36994 1737 36996 1775
rect 36996 1737 37048 1775
rect 37048 1737 37050 1775
rect 36994 1725 37050 1737
rect 36994 1719 36996 1725
rect 36996 1719 37048 1725
rect 37048 1719 37050 1725
rect 36994 1673 36996 1695
rect 36996 1673 37048 1695
rect 37048 1673 37050 1695
rect 36994 1661 37050 1673
rect 36994 1639 36996 1661
rect 36996 1639 37048 1661
rect 37048 1639 37050 1661
rect 36994 1609 36996 1615
rect 36996 1609 37048 1615
rect 37048 1609 37050 1615
rect 36994 1597 37050 1609
rect 36994 1559 36996 1597
rect 36996 1559 37048 1597
rect 37048 1559 37050 1597
rect 36994 1533 37050 1535
rect 36994 1481 36996 1533
rect 36996 1481 37048 1533
rect 37048 1481 37050 1533
rect 36994 1479 37050 1481
rect 36994 1417 36996 1455
rect 36996 1417 37048 1455
rect 37048 1417 37050 1455
rect 36994 1405 37050 1417
rect 36994 1399 36996 1405
rect 36996 1399 37048 1405
rect 37048 1399 37050 1405
rect 36994 1353 36996 1375
rect 36996 1353 37048 1375
rect 37048 1353 37050 1375
rect 36994 1341 37050 1353
rect 36994 1319 36996 1341
rect 36996 1319 37048 1341
rect 37048 1319 37050 1341
rect 36994 1289 36996 1295
rect 36996 1289 37048 1295
rect 37048 1289 37050 1295
rect 36994 1277 37050 1289
rect 36994 1239 36996 1277
rect 36996 1239 37048 1277
rect 37048 1239 37050 1277
rect 36994 1213 37050 1215
rect 36994 1161 36996 1213
rect 36996 1161 37048 1213
rect 37048 1161 37050 1213
rect 36994 1159 37050 1161
rect 37186 3133 37242 3135
rect 37186 3081 37188 3133
rect 37188 3081 37240 3133
rect 37240 3081 37242 3133
rect 37186 3079 37242 3081
rect 37186 3017 37188 3055
rect 37188 3017 37240 3055
rect 37240 3017 37242 3055
rect 37186 3005 37242 3017
rect 37186 2999 37188 3005
rect 37188 2999 37240 3005
rect 37240 2999 37242 3005
rect 37186 2953 37188 2975
rect 37188 2953 37240 2975
rect 37240 2953 37242 2975
rect 37186 2941 37242 2953
rect 37186 2919 37188 2941
rect 37188 2919 37240 2941
rect 37240 2919 37242 2941
rect 37186 2889 37188 2895
rect 37188 2889 37240 2895
rect 37240 2889 37242 2895
rect 37186 2877 37242 2889
rect 37186 2839 37188 2877
rect 37188 2839 37240 2877
rect 37240 2839 37242 2877
rect 37186 2813 37242 2815
rect 37186 2761 37188 2813
rect 37188 2761 37240 2813
rect 37240 2761 37242 2813
rect 37186 2759 37242 2761
rect 37186 2697 37188 2735
rect 37188 2697 37240 2735
rect 37240 2697 37242 2735
rect 37186 2685 37242 2697
rect 37186 2679 37188 2685
rect 37188 2679 37240 2685
rect 37240 2679 37242 2685
rect 37186 2633 37188 2655
rect 37188 2633 37240 2655
rect 37240 2633 37242 2655
rect 37186 2621 37242 2633
rect 37186 2599 37188 2621
rect 37188 2599 37240 2621
rect 37240 2599 37242 2621
rect 37186 2569 37188 2575
rect 37188 2569 37240 2575
rect 37240 2569 37242 2575
rect 37186 2557 37242 2569
rect 37186 2519 37188 2557
rect 37188 2519 37240 2557
rect 37240 2519 37242 2557
rect 37186 2493 37242 2495
rect 37186 2441 37188 2493
rect 37188 2441 37240 2493
rect 37240 2441 37242 2493
rect 37186 2439 37242 2441
rect 37186 2377 37188 2415
rect 37188 2377 37240 2415
rect 37240 2377 37242 2415
rect 37186 2365 37242 2377
rect 37186 2359 37188 2365
rect 37188 2359 37240 2365
rect 37240 2359 37242 2365
rect 37186 2313 37188 2335
rect 37188 2313 37240 2335
rect 37240 2313 37242 2335
rect 37186 2301 37242 2313
rect 37186 2279 37188 2301
rect 37188 2279 37240 2301
rect 37240 2279 37242 2301
rect 37186 2249 37188 2255
rect 37188 2249 37240 2255
rect 37240 2249 37242 2255
rect 37186 2237 37242 2249
rect 37186 2199 37188 2237
rect 37188 2199 37240 2237
rect 37240 2199 37242 2237
rect 37186 2173 37242 2175
rect 37186 2121 37188 2173
rect 37188 2121 37240 2173
rect 37240 2121 37242 2173
rect 37186 2119 37242 2121
rect 37186 2057 37188 2095
rect 37188 2057 37240 2095
rect 37240 2057 37242 2095
rect 37186 2045 37242 2057
rect 37186 2039 37188 2045
rect 37188 2039 37240 2045
rect 37240 2039 37242 2045
rect 37186 1993 37188 2015
rect 37188 1993 37240 2015
rect 37240 1993 37242 2015
rect 37186 1981 37242 1993
rect 37186 1959 37188 1981
rect 37188 1959 37240 1981
rect 37240 1959 37242 1981
rect 37186 1929 37188 1935
rect 37188 1929 37240 1935
rect 37240 1929 37242 1935
rect 37186 1917 37242 1929
rect 37186 1879 37188 1917
rect 37188 1879 37240 1917
rect 37240 1879 37242 1917
rect 37186 1853 37242 1855
rect 37186 1801 37188 1853
rect 37188 1801 37240 1853
rect 37240 1801 37242 1853
rect 37186 1799 37242 1801
rect 37186 1737 37188 1775
rect 37188 1737 37240 1775
rect 37240 1737 37242 1775
rect 37186 1725 37242 1737
rect 37186 1719 37188 1725
rect 37188 1719 37240 1725
rect 37240 1719 37242 1725
rect 37186 1673 37188 1695
rect 37188 1673 37240 1695
rect 37240 1673 37242 1695
rect 37186 1661 37242 1673
rect 37186 1639 37188 1661
rect 37188 1639 37240 1661
rect 37240 1639 37242 1661
rect 37186 1609 37188 1615
rect 37188 1609 37240 1615
rect 37240 1609 37242 1615
rect 37186 1597 37242 1609
rect 37186 1559 37188 1597
rect 37188 1559 37240 1597
rect 37240 1559 37242 1597
rect 37186 1533 37242 1535
rect 37186 1481 37188 1533
rect 37188 1481 37240 1533
rect 37240 1481 37242 1533
rect 37186 1479 37242 1481
rect 37186 1417 37188 1455
rect 37188 1417 37240 1455
rect 37240 1417 37242 1455
rect 37186 1405 37242 1417
rect 37186 1399 37188 1405
rect 37188 1399 37240 1405
rect 37240 1399 37242 1405
rect 37186 1353 37188 1375
rect 37188 1353 37240 1375
rect 37240 1353 37242 1375
rect 37186 1341 37242 1353
rect 37186 1319 37188 1341
rect 37188 1319 37240 1341
rect 37240 1319 37242 1341
rect 37186 1289 37188 1295
rect 37188 1289 37240 1295
rect 37240 1289 37242 1295
rect 37186 1277 37242 1289
rect 37186 1239 37188 1277
rect 37188 1239 37240 1277
rect 37240 1239 37242 1277
rect 37186 1213 37242 1215
rect 37186 1161 37188 1213
rect 37188 1161 37240 1213
rect 37240 1161 37242 1213
rect 37186 1159 37242 1161
rect 37378 3133 37434 3135
rect 37378 3081 37380 3133
rect 37380 3081 37432 3133
rect 37432 3081 37434 3133
rect 37378 3079 37434 3081
rect 37378 3017 37380 3055
rect 37380 3017 37432 3055
rect 37432 3017 37434 3055
rect 37378 3005 37434 3017
rect 37378 2999 37380 3005
rect 37380 2999 37432 3005
rect 37432 2999 37434 3005
rect 37378 2953 37380 2975
rect 37380 2953 37432 2975
rect 37432 2953 37434 2975
rect 37378 2941 37434 2953
rect 37378 2919 37380 2941
rect 37380 2919 37432 2941
rect 37432 2919 37434 2941
rect 37378 2889 37380 2895
rect 37380 2889 37432 2895
rect 37432 2889 37434 2895
rect 37378 2877 37434 2889
rect 37378 2839 37380 2877
rect 37380 2839 37432 2877
rect 37432 2839 37434 2877
rect 37378 2813 37434 2815
rect 37378 2761 37380 2813
rect 37380 2761 37432 2813
rect 37432 2761 37434 2813
rect 37378 2759 37434 2761
rect 37378 2697 37380 2735
rect 37380 2697 37432 2735
rect 37432 2697 37434 2735
rect 37378 2685 37434 2697
rect 37378 2679 37380 2685
rect 37380 2679 37432 2685
rect 37432 2679 37434 2685
rect 37378 2633 37380 2655
rect 37380 2633 37432 2655
rect 37432 2633 37434 2655
rect 37378 2621 37434 2633
rect 37378 2599 37380 2621
rect 37380 2599 37432 2621
rect 37432 2599 37434 2621
rect 37378 2569 37380 2575
rect 37380 2569 37432 2575
rect 37432 2569 37434 2575
rect 37378 2557 37434 2569
rect 37378 2519 37380 2557
rect 37380 2519 37432 2557
rect 37432 2519 37434 2557
rect 37378 2493 37434 2495
rect 37378 2441 37380 2493
rect 37380 2441 37432 2493
rect 37432 2441 37434 2493
rect 37378 2439 37434 2441
rect 37378 2377 37380 2415
rect 37380 2377 37432 2415
rect 37432 2377 37434 2415
rect 37378 2365 37434 2377
rect 37378 2359 37380 2365
rect 37380 2359 37432 2365
rect 37432 2359 37434 2365
rect 37378 2313 37380 2335
rect 37380 2313 37432 2335
rect 37432 2313 37434 2335
rect 37378 2301 37434 2313
rect 37378 2279 37380 2301
rect 37380 2279 37432 2301
rect 37432 2279 37434 2301
rect 37378 2249 37380 2255
rect 37380 2249 37432 2255
rect 37432 2249 37434 2255
rect 37378 2237 37434 2249
rect 37378 2199 37380 2237
rect 37380 2199 37432 2237
rect 37432 2199 37434 2237
rect 37378 2173 37434 2175
rect 37378 2121 37380 2173
rect 37380 2121 37432 2173
rect 37432 2121 37434 2173
rect 37378 2119 37434 2121
rect 37378 2057 37380 2095
rect 37380 2057 37432 2095
rect 37432 2057 37434 2095
rect 37378 2045 37434 2057
rect 37378 2039 37380 2045
rect 37380 2039 37432 2045
rect 37432 2039 37434 2045
rect 37378 1993 37380 2015
rect 37380 1993 37432 2015
rect 37432 1993 37434 2015
rect 37378 1981 37434 1993
rect 37378 1959 37380 1981
rect 37380 1959 37432 1981
rect 37432 1959 37434 1981
rect 37378 1929 37380 1935
rect 37380 1929 37432 1935
rect 37432 1929 37434 1935
rect 37378 1917 37434 1929
rect 37378 1879 37380 1917
rect 37380 1879 37432 1917
rect 37432 1879 37434 1917
rect 37378 1853 37434 1855
rect 37378 1801 37380 1853
rect 37380 1801 37432 1853
rect 37432 1801 37434 1853
rect 37378 1799 37434 1801
rect 37378 1737 37380 1775
rect 37380 1737 37432 1775
rect 37432 1737 37434 1775
rect 37378 1725 37434 1737
rect 37378 1719 37380 1725
rect 37380 1719 37432 1725
rect 37432 1719 37434 1725
rect 37378 1673 37380 1695
rect 37380 1673 37432 1695
rect 37432 1673 37434 1695
rect 37378 1661 37434 1673
rect 37378 1639 37380 1661
rect 37380 1639 37432 1661
rect 37432 1639 37434 1661
rect 37378 1609 37380 1615
rect 37380 1609 37432 1615
rect 37432 1609 37434 1615
rect 37378 1597 37434 1609
rect 37378 1559 37380 1597
rect 37380 1559 37432 1597
rect 37432 1559 37434 1597
rect 37378 1533 37434 1535
rect 37378 1481 37380 1533
rect 37380 1481 37432 1533
rect 37432 1481 37434 1533
rect 37378 1479 37434 1481
rect 37378 1417 37380 1455
rect 37380 1417 37432 1455
rect 37432 1417 37434 1455
rect 37378 1405 37434 1417
rect 37378 1399 37380 1405
rect 37380 1399 37432 1405
rect 37432 1399 37434 1405
rect 37378 1353 37380 1375
rect 37380 1353 37432 1375
rect 37432 1353 37434 1375
rect 37378 1341 37434 1353
rect 37378 1319 37380 1341
rect 37380 1319 37432 1341
rect 37432 1319 37434 1341
rect 37378 1289 37380 1295
rect 37380 1289 37432 1295
rect 37432 1289 37434 1295
rect 37378 1277 37434 1289
rect 37378 1239 37380 1277
rect 37380 1239 37432 1277
rect 37432 1239 37434 1277
rect 37378 1213 37434 1215
rect 37378 1161 37380 1213
rect 37380 1161 37432 1213
rect 37432 1161 37434 1213
rect 37378 1159 37434 1161
rect 37570 3133 37626 3135
rect 37570 3081 37572 3133
rect 37572 3081 37624 3133
rect 37624 3081 37626 3133
rect 37570 3079 37626 3081
rect 37570 3017 37572 3055
rect 37572 3017 37624 3055
rect 37624 3017 37626 3055
rect 37570 3005 37626 3017
rect 37570 2999 37572 3005
rect 37572 2999 37624 3005
rect 37624 2999 37626 3005
rect 37570 2953 37572 2975
rect 37572 2953 37624 2975
rect 37624 2953 37626 2975
rect 37570 2941 37626 2953
rect 37570 2919 37572 2941
rect 37572 2919 37624 2941
rect 37624 2919 37626 2941
rect 37570 2889 37572 2895
rect 37572 2889 37624 2895
rect 37624 2889 37626 2895
rect 37570 2877 37626 2889
rect 37570 2839 37572 2877
rect 37572 2839 37624 2877
rect 37624 2839 37626 2877
rect 37570 2813 37626 2815
rect 37570 2761 37572 2813
rect 37572 2761 37624 2813
rect 37624 2761 37626 2813
rect 37570 2759 37626 2761
rect 37570 2697 37572 2735
rect 37572 2697 37624 2735
rect 37624 2697 37626 2735
rect 37570 2685 37626 2697
rect 37570 2679 37572 2685
rect 37572 2679 37624 2685
rect 37624 2679 37626 2685
rect 37570 2633 37572 2655
rect 37572 2633 37624 2655
rect 37624 2633 37626 2655
rect 37570 2621 37626 2633
rect 37570 2599 37572 2621
rect 37572 2599 37624 2621
rect 37624 2599 37626 2621
rect 37570 2569 37572 2575
rect 37572 2569 37624 2575
rect 37624 2569 37626 2575
rect 37570 2557 37626 2569
rect 37570 2519 37572 2557
rect 37572 2519 37624 2557
rect 37624 2519 37626 2557
rect 37570 2493 37626 2495
rect 37570 2441 37572 2493
rect 37572 2441 37624 2493
rect 37624 2441 37626 2493
rect 37570 2439 37626 2441
rect 37570 2377 37572 2415
rect 37572 2377 37624 2415
rect 37624 2377 37626 2415
rect 37570 2365 37626 2377
rect 37570 2359 37572 2365
rect 37572 2359 37624 2365
rect 37624 2359 37626 2365
rect 37570 2313 37572 2335
rect 37572 2313 37624 2335
rect 37624 2313 37626 2335
rect 37570 2301 37626 2313
rect 37570 2279 37572 2301
rect 37572 2279 37624 2301
rect 37624 2279 37626 2301
rect 37570 2249 37572 2255
rect 37572 2249 37624 2255
rect 37624 2249 37626 2255
rect 37570 2237 37626 2249
rect 37570 2199 37572 2237
rect 37572 2199 37624 2237
rect 37624 2199 37626 2237
rect 37570 2173 37626 2175
rect 37570 2121 37572 2173
rect 37572 2121 37624 2173
rect 37624 2121 37626 2173
rect 37570 2119 37626 2121
rect 37570 2057 37572 2095
rect 37572 2057 37624 2095
rect 37624 2057 37626 2095
rect 37570 2045 37626 2057
rect 37570 2039 37572 2045
rect 37572 2039 37624 2045
rect 37624 2039 37626 2045
rect 37570 1993 37572 2015
rect 37572 1993 37624 2015
rect 37624 1993 37626 2015
rect 37570 1981 37626 1993
rect 37570 1959 37572 1981
rect 37572 1959 37624 1981
rect 37624 1959 37626 1981
rect 37570 1929 37572 1935
rect 37572 1929 37624 1935
rect 37624 1929 37626 1935
rect 37570 1917 37626 1929
rect 37570 1879 37572 1917
rect 37572 1879 37624 1917
rect 37624 1879 37626 1917
rect 37570 1853 37626 1855
rect 37570 1801 37572 1853
rect 37572 1801 37624 1853
rect 37624 1801 37626 1853
rect 37570 1799 37626 1801
rect 37570 1737 37572 1775
rect 37572 1737 37624 1775
rect 37624 1737 37626 1775
rect 37570 1725 37626 1737
rect 37570 1719 37572 1725
rect 37572 1719 37624 1725
rect 37624 1719 37626 1725
rect 37570 1673 37572 1695
rect 37572 1673 37624 1695
rect 37624 1673 37626 1695
rect 37570 1661 37626 1673
rect 37570 1639 37572 1661
rect 37572 1639 37624 1661
rect 37624 1639 37626 1661
rect 37570 1609 37572 1615
rect 37572 1609 37624 1615
rect 37624 1609 37626 1615
rect 37570 1597 37626 1609
rect 37570 1559 37572 1597
rect 37572 1559 37624 1597
rect 37624 1559 37626 1597
rect 37570 1533 37626 1535
rect 37570 1481 37572 1533
rect 37572 1481 37624 1533
rect 37624 1481 37626 1533
rect 37570 1479 37626 1481
rect 37570 1417 37572 1455
rect 37572 1417 37624 1455
rect 37624 1417 37626 1455
rect 37570 1405 37626 1417
rect 37570 1399 37572 1405
rect 37572 1399 37624 1405
rect 37624 1399 37626 1405
rect 37570 1353 37572 1375
rect 37572 1353 37624 1375
rect 37624 1353 37626 1375
rect 37570 1341 37626 1353
rect 37570 1319 37572 1341
rect 37572 1319 37624 1341
rect 37624 1319 37626 1341
rect 37570 1289 37572 1295
rect 37572 1289 37624 1295
rect 37624 1289 37626 1295
rect 37570 1277 37626 1289
rect 37570 1239 37572 1277
rect 37572 1239 37624 1277
rect 37624 1239 37626 1277
rect 37570 1213 37626 1215
rect 37570 1161 37572 1213
rect 37572 1161 37624 1213
rect 37624 1161 37626 1213
rect 37570 1159 37626 1161
rect 37762 3133 37818 3135
rect 37762 3081 37764 3133
rect 37764 3081 37816 3133
rect 37816 3081 37818 3133
rect 37762 3079 37818 3081
rect 37762 3017 37764 3055
rect 37764 3017 37816 3055
rect 37816 3017 37818 3055
rect 37762 3005 37818 3017
rect 37762 2999 37764 3005
rect 37764 2999 37816 3005
rect 37816 2999 37818 3005
rect 37762 2953 37764 2975
rect 37764 2953 37816 2975
rect 37816 2953 37818 2975
rect 37762 2941 37818 2953
rect 37762 2919 37764 2941
rect 37764 2919 37816 2941
rect 37816 2919 37818 2941
rect 37762 2889 37764 2895
rect 37764 2889 37816 2895
rect 37816 2889 37818 2895
rect 37762 2877 37818 2889
rect 37762 2839 37764 2877
rect 37764 2839 37816 2877
rect 37816 2839 37818 2877
rect 37762 2813 37818 2815
rect 37762 2761 37764 2813
rect 37764 2761 37816 2813
rect 37816 2761 37818 2813
rect 37762 2759 37818 2761
rect 37762 2697 37764 2735
rect 37764 2697 37816 2735
rect 37816 2697 37818 2735
rect 37762 2685 37818 2697
rect 37762 2679 37764 2685
rect 37764 2679 37816 2685
rect 37816 2679 37818 2685
rect 37762 2633 37764 2655
rect 37764 2633 37816 2655
rect 37816 2633 37818 2655
rect 37762 2621 37818 2633
rect 37762 2599 37764 2621
rect 37764 2599 37816 2621
rect 37816 2599 37818 2621
rect 37762 2569 37764 2575
rect 37764 2569 37816 2575
rect 37816 2569 37818 2575
rect 37762 2557 37818 2569
rect 37762 2519 37764 2557
rect 37764 2519 37816 2557
rect 37816 2519 37818 2557
rect 37762 2493 37818 2495
rect 37762 2441 37764 2493
rect 37764 2441 37816 2493
rect 37816 2441 37818 2493
rect 37762 2439 37818 2441
rect 37762 2377 37764 2415
rect 37764 2377 37816 2415
rect 37816 2377 37818 2415
rect 37762 2365 37818 2377
rect 37762 2359 37764 2365
rect 37764 2359 37816 2365
rect 37816 2359 37818 2365
rect 37762 2313 37764 2335
rect 37764 2313 37816 2335
rect 37816 2313 37818 2335
rect 37762 2301 37818 2313
rect 37762 2279 37764 2301
rect 37764 2279 37816 2301
rect 37816 2279 37818 2301
rect 37762 2249 37764 2255
rect 37764 2249 37816 2255
rect 37816 2249 37818 2255
rect 37762 2237 37818 2249
rect 37762 2199 37764 2237
rect 37764 2199 37816 2237
rect 37816 2199 37818 2237
rect 37762 2173 37818 2175
rect 37762 2121 37764 2173
rect 37764 2121 37816 2173
rect 37816 2121 37818 2173
rect 37762 2119 37818 2121
rect 37762 2057 37764 2095
rect 37764 2057 37816 2095
rect 37816 2057 37818 2095
rect 37762 2045 37818 2057
rect 37762 2039 37764 2045
rect 37764 2039 37816 2045
rect 37816 2039 37818 2045
rect 37762 1993 37764 2015
rect 37764 1993 37816 2015
rect 37816 1993 37818 2015
rect 37762 1981 37818 1993
rect 37762 1959 37764 1981
rect 37764 1959 37816 1981
rect 37816 1959 37818 1981
rect 37762 1929 37764 1935
rect 37764 1929 37816 1935
rect 37816 1929 37818 1935
rect 37762 1917 37818 1929
rect 37762 1879 37764 1917
rect 37764 1879 37816 1917
rect 37816 1879 37818 1917
rect 37762 1853 37818 1855
rect 37762 1801 37764 1853
rect 37764 1801 37816 1853
rect 37816 1801 37818 1853
rect 37762 1799 37818 1801
rect 37762 1737 37764 1775
rect 37764 1737 37816 1775
rect 37816 1737 37818 1775
rect 37762 1725 37818 1737
rect 37762 1719 37764 1725
rect 37764 1719 37816 1725
rect 37816 1719 37818 1725
rect 37762 1673 37764 1695
rect 37764 1673 37816 1695
rect 37816 1673 37818 1695
rect 37762 1661 37818 1673
rect 37762 1639 37764 1661
rect 37764 1639 37816 1661
rect 37816 1639 37818 1661
rect 37762 1609 37764 1615
rect 37764 1609 37816 1615
rect 37816 1609 37818 1615
rect 37762 1597 37818 1609
rect 37762 1559 37764 1597
rect 37764 1559 37816 1597
rect 37816 1559 37818 1597
rect 37762 1533 37818 1535
rect 37762 1481 37764 1533
rect 37764 1481 37816 1533
rect 37816 1481 37818 1533
rect 37762 1479 37818 1481
rect 37762 1417 37764 1455
rect 37764 1417 37816 1455
rect 37816 1417 37818 1455
rect 37762 1405 37818 1417
rect 37762 1399 37764 1405
rect 37764 1399 37816 1405
rect 37816 1399 37818 1405
rect 37762 1353 37764 1375
rect 37764 1353 37816 1375
rect 37816 1353 37818 1375
rect 37762 1341 37818 1353
rect 37762 1319 37764 1341
rect 37764 1319 37816 1341
rect 37816 1319 37818 1341
rect 37762 1289 37764 1295
rect 37764 1289 37816 1295
rect 37816 1289 37818 1295
rect 37762 1277 37818 1289
rect 37762 1239 37764 1277
rect 37764 1239 37816 1277
rect 37816 1239 37818 1277
rect 37762 1213 37818 1215
rect 37762 1161 37764 1213
rect 37764 1161 37816 1213
rect 37816 1161 37818 1213
rect 37762 1159 37818 1161
rect 37954 3133 38010 3135
rect 37954 3081 37956 3133
rect 37956 3081 38008 3133
rect 38008 3081 38010 3133
rect 37954 3079 38010 3081
rect 37954 3017 37956 3055
rect 37956 3017 38008 3055
rect 38008 3017 38010 3055
rect 37954 3005 38010 3017
rect 37954 2999 37956 3005
rect 37956 2999 38008 3005
rect 38008 2999 38010 3005
rect 37954 2953 37956 2975
rect 37956 2953 38008 2975
rect 38008 2953 38010 2975
rect 37954 2941 38010 2953
rect 37954 2919 37956 2941
rect 37956 2919 38008 2941
rect 38008 2919 38010 2941
rect 37954 2889 37956 2895
rect 37956 2889 38008 2895
rect 38008 2889 38010 2895
rect 37954 2877 38010 2889
rect 37954 2839 37956 2877
rect 37956 2839 38008 2877
rect 38008 2839 38010 2877
rect 37954 2813 38010 2815
rect 37954 2761 37956 2813
rect 37956 2761 38008 2813
rect 38008 2761 38010 2813
rect 37954 2759 38010 2761
rect 37954 2697 37956 2735
rect 37956 2697 38008 2735
rect 38008 2697 38010 2735
rect 37954 2685 38010 2697
rect 37954 2679 37956 2685
rect 37956 2679 38008 2685
rect 38008 2679 38010 2685
rect 37954 2633 37956 2655
rect 37956 2633 38008 2655
rect 38008 2633 38010 2655
rect 37954 2621 38010 2633
rect 37954 2599 37956 2621
rect 37956 2599 38008 2621
rect 38008 2599 38010 2621
rect 37954 2569 37956 2575
rect 37956 2569 38008 2575
rect 38008 2569 38010 2575
rect 37954 2557 38010 2569
rect 37954 2519 37956 2557
rect 37956 2519 38008 2557
rect 38008 2519 38010 2557
rect 37954 2493 38010 2495
rect 37954 2441 37956 2493
rect 37956 2441 38008 2493
rect 38008 2441 38010 2493
rect 37954 2439 38010 2441
rect 37954 2377 37956 2415
rect 37956 2377 38008 2415
rect 38008 2377 38010 2415
rect 37954 2365 38010 2377
rect 37954 2359 37956 2365
rect 37956 2359 38008 2365
rect 38008 2359 38010 2365
rect 37954 2313 37956 2335
rect 37956 2313 38008 2335
rect 38008 2313 38010 2335
rect 37954 2301 38010 2313
rect 37954 2279 37956 2301
rect 37956 2279 38008 2301
rect 38008 2279 38010 2301
rect 37954 2249 37956 2255
rect 37956 2249 38008 2255
rect 38008 2249 38010 2255
rect 37954 2237 38010 2249
rect 37954 2199 37956 2237
rect 37956 2199 38008 2237
rect 38008 2199 38010 2237
rect 37954 2173 38010 2175
rect 37954 2121 37956 2173
rect 37956 2121 38008 2173
rect 38008 2121 38010 2173
rect 37954 2119 38010 2121
rect 37954 2057 37956 2095
rect 37956 2057 38008 2095
rect 38008 2057 38010 2095
rect 37954 2045 38010 2057
rect 37954 2039 37956 2045
rect 37956 2039 38008 2045
rect 38008 2039 38010 2045
rect 37954 1993 37956 2015
rect 37956 1993 38008 2015
rect 38008 1993 38010 2015
rect 37954 1981 38010 1993
rect 37954 1959 37956 1981
rect 37956 1959 38008 1981
rect 38008 1959 38010 1981
rect 37954 1929 37956 1935
rect 37956 1929 38008 1935
rect 38008 1929 38010 1935
rect 37954 1917 38010 1929
rect 37954 1879 37956 1917
rect 37956 1879 38008 1917
rect 38008 1879 38010 1917
rect 37954 1853 38010 1855
rect 37954 1801 37956 1853
rect 37956 1801 38008 1853
rect 38008 1801 38010 1853
rect 37954 1799 38010 1801
rect 37954 1737 37956 1775
rect 37956 1737 38008 1775
rect 38008 1737 38010 1775
rect 37954 1725 38010 1737
rect 37954 1719 37956 1725
rect 37956 1719 38008 1725
rect 38008 1719 38010 1725
rect 37954 1673 37956 1695
rect 37956 1673 38008 1695
rect 38008 1673 38010 1695
rect 37954 1661 38010 1673
rect 37954 1639 37956 1661
rect 37956 1639 38008 1661
rect 38008 1639 38010 1661
rect 37954 1609 37956 1615
rect 37956 1609 38008 1615
rect 38008 1609 38010 1615
rect 37954 1597 38010 1609
rect 37954 1559 37956 1597
rect 37956 1559 38008 1597
rect 38008 1559 38010 1597
rect 37954 1533 38010 1535
rect 37954 1481 37956 1533
rect 37956 1481 38008 1533
rect 38008 1481 38010 1533
rect 37954 1479 38010 1481
rect 37954 1417 37956 1455
rect 37956 1417 38008 1455
rect 38008 1417 38010 1455
rect 37954 1405 38010 1417
rect 37954 1399 37956 1405
rect 37956 1399 38008 1405
rect 38008 1399 38010 1405
rect 37954 1353 37956 1375
rect 37956 1353 38008 1375
rect 38008 1353 38010 1375
rect 37954 1341 38010 1353
rect 37954 1319 37956 1341
rect 37956 1319 38008 1341
rect 38008 1319 38010 1341
rect 37954 1289 37956 1295
rect 37956 1289 38008 1295
rect 38008 1289 38010 1295
rect 37954 1277 38010 1289
rect 37954 1239 37956 1277
rect 37956 1239 38008 1277
rect 38008 1239 38010 1277
rect 37954 1213 38010 1215
rect 37954 1161 37956 1213
rect 37956 1161 38008 1213
rect 38008 1161 38010 1213
rect 37954 1159 38010 1161
rect 38146 3133 38202 3135
rect 38146 3081 38148 3133
rect 38148 3081 38200 3133
rect 38200 3081 38202 3133
rect 38146 3079 38202 3081
rect 38146 3017 38148 3055
rect 38148 3017 38200 3055
rect 38200 3017 38202 3055
rect 38146 3005 38202 3017
rect 38146 2999 38148 3005
rect 38148 2999 38200 3005
rect 38200 2999 38202 3005
rect 38146 2953 38148 2975
rect 38148 2953 38200 2975
rect 38200 2953 38202 2975
rect 38146 2941 38202 2953
rect 38146 2919 38148 2941
rect 38148 2919 38200 2941
rect 38200 2919 38202 2941
rect 38146 2889 38148 2895
rect 38148 2889 38200 2895
rect 38200 2889 38202 2895
rect 38146 2877 38202 2889
rect 38146 2839 38148 2877
rect 38148 2839 38200 2877
rect 38200 2839 38202 2877
rect 38146 2813 38202 2815
rect 38146 2761 38148 2813
rect 38148 2761 38200 2813
rect 38200 2761 38202 2813
rect 38146 2759 38202 2761
rect 38146 2697 38148 2735
rect 38148 2697 38200 2735
rect 38200 2697 38202 2735
rect 38146 2685 38202 2697
rect 38146 2679 38148 2685
rect 38148 2679 38200 2685
rect 38200 2679 38202 2685
rect 38146 2633 38148 2655
rect 38148 2633 38200 2655
rect 38200 2633 38202 2655
rect 38146 2621 38202 2633
rect 38146 2599 38148 2621
rect 38148 2599 38200 2621
rect 38200 2599 38202 2621
rect 38146 2569 38148 2575
rect 38148 2569 38200 2575
rect 38200 2569 38202 2575
rect 38146 2557 38202 2569
rect 38146 2519 38148 2557
rect 38148 2519 38200 2557
rect 38200 2519 38202 2557
rect 38146 2493 38202 2495
rect 38146 2441 38148 2493
rect 38148 2441 38200 2493
rect 38200 2441 38202 2493
rect 38146 2439 38202 2441
rect 38146 2377 38148 2415
rect 38148 2377 38200 2415
rect 38200 2377 38202 2415
rect 38146 2365 38202 2377
rect 38146 2359 38148 2365
rect 38148 2359 38200 2365
rect 38200 2359 38202 2365
rect 38146 2313 38148 2335
rect 38148 2313 38200 2335
rect 38200 2313 38202 2335
rect 38146 2301 38202 2313
rect 38146 2279 38148 2301
rect 38148 2279 38200 2301
rect 38200 2279 38202 2301
rect 38146 2249 38148 2255
rect 38148 2249 38200 2255
rect 38200 2249 38202 2255
rect 38146 2237 38202 2249
rect 38146 2199 38148 2237
rect 38148 2199 38200 2237
rect 38200 2199 38202 2237
rect 38146 2173 38202 2175
rect 38146 2121 38148 2173
rect 38148 2121 38200 2173
rect 38200 2121 38202 2173
rect 38146 2119 38202 2121
rect 38146 2057 38148 2095
rect 38148 2057 38200 2095
rect 38200 2057 38202 2095
rect 38146 2045 38202 2057
rect 38146 2039 38148 2045
rect 38148 2039 38200 2045
rect 38200 2039 38202 2045
rect 38146 1993 38148 2015
rect 38148 1993 38200 2015
rect 38200 1993 38202 2015
rect 38146 1981 38202 1993
rect 38146 1959 38148 1981
rect 38148 1959 38200 1981
rect 38200 1959 38202 1981
rect 38146 1929 38148 1935
rect 38148 1929 38200 1935
rect 38200 1929 38202 1935
rect 38146 1917 38202 1929
rect 38146 1879 38148 1917
rect 38148 1879 38200 1917
rect 38200 1879 38202 1917
rect 38146 1853 38202 1855
rect 38146 1801 38148 1853
rect 38148 1801 38200 1853
rect 38200 1801 38202 1853
rect 38146 1799 38202 1801
rect 38146 1737 38148 1775
rect 38148 1737 38200 1775
rect 38200 1737 38202 1775
rect 38146 1725 38202 1737
rect 38146 1719 38148 1725
rect 38148 1719 38200 1725
rect 38200 1719 38202 1725
rect 38146 1673 38148 1695
rect 38148 1673 38200 1695
rect 38200 1673 38202 1695
rect 38146 1661 38202 1673
rect 38146 1639 38148 1661
rect 38148 1639 38200 1661
rect 38200 1639 38202 1661
rect 38146 1609 38148 1615
rect 38148 1609 38200 1615
rect 38200 1609 38202 1615
rect 38146 1597 38202 1609
rect 38146 1559 38148 1597
rect 38148 1559 38200 1597
rect 38200 1559 38202 1597
rect 38146 1533 38202 1535
rect 38146 1481 38148 1533
rect 38148 1481 38200 1533
rect 38200 1481 38202 1533
rect 38146 1479 38202 1481
rect 38146 1417 38148 1455
rect 38148 1417 38200 1455
rect 38200 1417 38202 1455
rect 38146 1405 38202 1417
rect 38146 1399 38148 1405
rect 38148 1399 38200 1405
rect 38200 1399 38202 1405
rect 38146 1353 38148 1375
rect 38148 1353 38200 1375
rect 38200 1353 38202 1375
rect 38146 1341 38202 1353
rect 38146 1319 38148 1341
rect 38148 1319 38200 1341
rect 38200 1319 38202 1341
rect 38146 1289 38148 1295
rect 38148 1289 38200 1295
rect 38200 1289 38202 1295
rect 38146 1277 38202 1289
rect 38146 1239 38148 1277
rect 38148 1239 38200 1277
rect 38200 1239 38202 1277
rect 38146 1213 38202 1215
rect 38146 1161 38148 1213
rect 38148 1161 38200 1213
rect 38200 1161 38202 1213
rect 38146 1159 38202 1161
rect 38338 3133 38394 3135
rect 38338 3081 38340 3133
rect 38340 3081 38392 3133
rect 38392 3081 38394 3133
rect 38338 3079 38394 3081
rect 38338 3017 38340 3055
rect 38340 3017 38392 3055
rect 38392 3017 38394 3055
rect 38338 3005 38394 3017
rect 38338 2999 38340 3005
rect 38340 2999 38392 3005
rect 38392 2999 38394 3005
rect 38338 2953 38340 2975
rect 38340 2953 38392 2975
rect 38392 2953 38394 2975
rect 38338 2941 38394 2953
rect 38338 2919 38340 2941
rect 38340 2919 38392 2941
rect 38392 2919 38394 2941
rect 38338 2889 38340 2895
rect 38340 2889 38392 2895
rect 38392 2889 38394 2895
rect 38338 2877 38394 2889
rect 38338 2839 38340 2877
rect 38340 2839 38392 2877
rect 38392 2839 38394 2877
rect 38338 2813 38394 2815
rect 38338 2761 38340 2813
rect 38340 2761 38392 2813
rect 38392 2761 38394 2813
rect 38338 2759 38394 2761
rect 38338 2697 38340 2735
rect 38340 2697 38392 2735
rect 38392 2697 38394 2735
rect 38338 2685 38394 2697
rect 38338 2679 38340 2685
rect 38340 2679 38392 2685
rect 38392 2679 38394 2685
rect 38338 2633 38340 2655
rect 38340 2633 38392 2655
rect 38392 2633 38394 2655
rect 38338 2621 38394 2633
rect 38338 2599 38340 2621
rect 38340 2599 38392 2621
rect 38392 2599 38394 2621
rect 38338 2569 38340 2575
rect 38340 2569 38392 2575
rect 38392 2569 38394 2575
rect 38338 2557 38394 2569
rect 38338 2519 38340 2557
rect 38340 2519 38392 2557
rect 38392 2519 38394 2557
rect 38338 2493 38394 2495
rect 38338 2441 38340 2493
rect 38340 2441 38392 2493
rect 38392 2441 38394 2493
rect 38338 2439 38394 2441
rect 38338 2377 38340 2415
rect 38340 2377 38392 2415
rect 38392 2377 38394 2415
rect 38338 2365 38394 2377
rect 38338 2359 38340 2365
rect 38340 2359 38392 2365
rect 38392 2359 38394 2365
rect 38338 2313 38340 2335
rect 38340 2313 38392 2335
rect 38392 2313 38394 2335
rect 38338 2301 38394 2313
rect 38338 2279 38340 2301
rect 38340 2279 38392 2301
rect 38392 2279 38394 2301
rect 38338 2249 38340 2255
rect 38340 2249 38392 2255
rect 38392 2249 38394 2255
rect 38338 2237 38394 2249
rect 38338 2199 38340 2237
rect 38340 2199 38392 2237
rect 38392 2199 38394 2237
rect 38338 2173 38394 2175
rect 38338 2121 38340 2173
rect 38340 2121 38392 2173
rect 38392 2121 38394 2173
rect 38338 2119 38394 2121
rect 38338 2057 38340 2095
rect 38340 2057 38392 2095
rect 38392 2057 38394 2095
rect 38338 2045 38394 2057
rect 38338 2039 38340 2045
rect 38340 2039 38392 2045
rect 38392 2039 38394 2045
rect 38338 1993 38340 2015
rect 38340 1993 38392 2015
rect 38392 1993 38394 2015
rect 38338 1981 38394 1993
rect 38338 1959 38340 1981
rect 38340 1959 38392 1981
rect 38392 1959 38394 1981
rect 38338 1929 38340 1935
rect 38340 1929 38392 1935
rect 38392 1929 38394 1935
rect 38338 1917 38394 1929
rect 38338 1879 38340 1917
rect 38340 1879 38392 1917
rect 38392 1879 38394 1917
rect 38338 1853 38394 1855
rect 38338 1801 38340 1853
rect 38340 1801 38392 1853
rect 38392 1801 38394 1853
rect 38338 1799 38394 1801
rect 38338 1737 38340 1775
rect 38340 1737 38392 1775
rect 38392 1737 38394 1775
rect 38338 1725 38394 1737
rect 38338 1719 38340 1725
rect 38340 1719 38392 1725
rect 38392 1719 38394 1725
rect 38338 1673 38340 1695
rect 38340 1673 38392 1695
rect 38392 1673 38394 1695
rect 38338 1661 38394 1673
rect 38338 1639 38340 1661
rect 38340 1639 38392 1661
rect 38392 1639 38394 1661
rect 38338 1609 38340 1615
rect 38340 1609 38392 1615
rect 38392 1609 38394 1615
rect 38338 1597 38394 1609
rect 38338 1559 38340 1597
rect 38340 1559 38392 1597
rect 38392 1559 38394 1597
rect 38338 1533 38394 1535
rect 38338 1481 38340 1533
rect 38340 1481 38392 1533
rect 38392 1481 38394 1533
rect 38338 1479 38394 1481
rect 38338 1417 38340 1455
rect 38340 1417 38392 1455
rect 38392 1417 38394 1455
rect 38338 1405 38394 1417
rect 38338 1399 38340 1405
rect 38340 1399 38392 1405
rect 38392 1399 38394 1405
rect 38338 1353 38340 1375
rect 38340 1353 38392 1375
rect 38392 1353 38394 1375
rect 38338 1341 38394 1353
rect 38338 1319 38340 1341
rect 38340 1319 38392 1341
rect 38392 1319 38394 1341
rect 38338 1289 38340 1295
rect 38340 1289 38392 1295
rect 38392 1289 38394 1295
rect 38338 1277 38394 1289
rect 38338 1239 38340 1277
rect 38340 1239 38392 1277
rect 38392 1239 38394 1277
rect 38338 1213 38394 1215
rect 38338 1161 38340 1213
rect 38340 1161 38392 1213
rect 38392 1161 38394 1213
rect 38338 1159 38394 1161
rect 38530 3133 38586 3135
rect 38530 3081 38532 3133
rect 38532 3081 38584 3133
rect 38584 3081 38586 3133
rect 38530 3079 38586 3081
rect 38530 3017 38532 3055
rect 38532 3017 38584 3055
rect 38584 3017 38586 3055
rect 38530 3005 38586 3017
rect 38530 2999 38532 3005
rect 38532 2999 38584 3005
rect 38584 2999 38586 3005
rect 38530 2953 38532 2975
rect 38532 2953 38584 2975
rect 38584 2953 38586 2975
rect 38530 2941 38586 2953
rect 38530 2919 38532 2941
rect 38532 2919 38584 2941
rect 38584 2919 38586 2941
rect 38530 2889 38532 2895
rect 38532 2889 38584 2895
rect 38584 2889 38586 2895
rect 38530 2877 38586 2889
rect 38530 2839 38532 2877
rect 38532 2839 38584 2877
rect 38584 2839 38586 2877
rect 38530 2813 38586 2815
rect 38530 2761 38532 2813
rect 38532 2761 38584 2813
rect 38584 2761 38586 2813
rect 38530 2759 38586 2761
rect 38530 2697 38532 2735
rect 38532 2697 38584 2735
rect 38584 2697 38586 2735
rect 38530 2685 38586 2697
rect 38530 2679 38532 2685
rect 38532 2679 38584 2685
rect 38584 2679 38586 2685
rect 38530 2633 38532 2655
rect 38532 2633 38584 2655
rect 38584 2633 38586 2655
rect 38530 2621 38586 2633
rect 38530 2599 38532 2621
rect 38532 2599 38584 2621
rect 38584 2599 38586 2621
rect 38530 2569 38532 2575
rect 38532 2569 38584 2575
rect 38584 2569 38586 2575
rect 38530 2557 38586 2569
rect 38530 2519 38532 2557
rect 38532 2519 38584 2557
rect 38584 2519 38586 2557
rect 38530 2493 38586 2495
rect 38530 2441 38532 2493
rect 38532 2441 38584 2493
rect 38584 2441 38586 2493
rect 38530 2439 38586 2441
rect 38530 2377 38532 2415
rect 38532 2377 38584 2415
rect 38584 2377 38586 2415
rect 38530 2365 38586 2377
rect 38530 2359 38532 2365
rect 38532 2359 38584 2365
rect 38584 2359 38586 2365
rect 38530 2313 38532 2335
rect 38532 2313 38584 2335
rect 38584 2313 38586 2335
rect 38530 2301 38586 2313
rect 38530 2279 38532 2301
rect 38532 2279 38584 2301
rect 38584 2279 38586 2301
rect 38530 2249 38532 2255
rect 38532 2249 38584 2255
rect 38584 2249 38586 2255
rect 38530 2237 38586 2249
rect 38530 2199 38532 2237
rect 38532 2199 38584 2237
rect 38584 2199 38586 2237
rect 38530 2173 38586 2175
rect 38530 2121 38532 2173
rect 38532 2121 38584 2173
rect 38584 2121 38586 2173
rect 38530 2119 38586 2121
rect 38530 2057 38532 2095
rect 38532 2057 38584 2095
rect 38584 2057 38586 2095
rect 38530 2045 38586 2057
rect 38530 2039 38532 2045
rect 38532 2039 38584 2045
rect 38584 2039 38586 2045
rect 38530 1993 38532 2015
rect 38532 1993 38584 2015
rect 38584 1993 38586 2015
rect 38530 1981 38586 1993
rect 38530 1959 38532 1981
rect 38532 1959 38584 1981
rect 38584 1959 38586 1981
rect 38530 1929 38532 1935
rect 38532 1929 38584 1935
rect 38584 1929 38586 1935
rect 38530 1917 38586 1929
rect 38530 1879 38532 1917
rect 38532 1879 38584 1917
rect 38584 1879 38586 1917
rect 38530 1853 38586 1855
rect 38530 1801 38532 1853
rect 38532 1801 38584 1853
rect 38584 1801 38586 1853
rect 38530 1799 38586 1801
rect 38530 1737 38532 1775
rect 38532 1737 38584 1775
rect 38584 1737 38586 1775
rect 38530 1725 38586 1737
rect 38530 1719 38532 1725
rect 38532 1719 38584 1725
rect 38584 1719 38586 1725
rect 38530 1673 38532 1695
rect 38532 1673 38584 1695
rect 38584 1673 38586 1695
rect 38530 1661 38586 1673
rect 38530 1639 38532 1661
rect 38532 1639 38584 1661
rect 38584 1639 38586 1661
rect 38530 1609 38532 1615
rect 38532 1609 38584 1615
rect 38584 1609 38586 1615
rect 38530 1597 38586 1609
rect 38530 1559 38532 1597
rect 38532 1559 38584 1597
rect 38584 1559 38586 1597
rect 38530 1533 38586 1535
rect 38530 1481 38532 1533
rect 38532 1481 38584 1533
rect 38584 1481 38586 1533
rect 38530 1479 38586 1481
rect 38530 1417 38532 1455
rect 38532 1417 38584 1455
rect 38584 1417 38586 1455
rect 38530 1405 38586 1417
rect 38530 1399 38532 1405
rect 38532 1399 38584 1405
rect 38584 1399 38586 1405
rect 38530 1353 38532 1375
rect 38532 1353 38584 1375
rect 38584 1353 38586 1375
rect 38530 1341 38586 1353
rect 38530 1319 38532 1341
rect 38532 1319 38584 1341
rect 38584 1319 38586 1341
rect 38530 1289 38532 1295
rect 38532 1289 38584 1295
rect 38584 1289 38586 1295
rect 38530 1277 38586 1289
rect 38530 1239 38532 1277
rect 38532 1239 38584 1277
rect 38584 1239 38586 1277
rect 38530 1213 38586 1215
rect 38530 1161 38532 1213
rect 38532 1161 38584 1213
rect 38584 1161 38586 1213
rect 38530 1159 38586 1161
<< metal3 >>
rect 29116 3522 38592 3606
rect 29116 3135 29184 3522
rect 29116 3079 29122 3135
rect 29178 3079 29184 3135
rect 29116 3055 29184 3079
rect 29116 2999 29122 3055
rect 29178 2999 29184 3055
rect 29116 2975 29184 2999
rect 29116 2919 29122 2975
rect 29178 2919 29184 2975
rect 29116 2895 29184 2919
rect 29116 2839 29122 2895
rect 29178 2839 29184 2895
rect 29116 2815 29184 2839
rect 29116 2759 29122 2815
rect 29178 2759 29184 2815
rect 29116 2735 29184 2759
rect 29116 2679 29122 2735
rect 29178 2679 29184 2735
rect 29116 2655 29184 2679
rect 29116 2599 29122 2655
rect 29178 2599 29184 2655
rect 29116 2575 29184 2599
rect 29116 2519 29122 2575
rect 29178 2519 29184 2575
rect 29116 2495 29184 2519
rect 29116 2439 29122 2495
rect 29178 2439 29184 2495
rect 29116 2415 29184 2439
rect 29116 2359 29122 2415
rect 29178 2359 29184 2415
rect 29116 2335 29184 2359
rect 29116 2279 29122 2335
rect 29178 2279 29184 2335
rect 29116 2255 29184 2279
rect 29116 2199 29122 2255
rect 29178 2199 29184 2255
rect 29116 2175 29184 2199
rect 29116 2119 29122 2175
rect 29178 2119 29184 2175
rect 29116 2095 29184 2119
rect 29116 2039 29122 2095
rect 29178 2039 29184 2095
rect 29116 2015 29184 2039
rect 29116 1959 29122 2015
rect 29178 1959 29184 2015
rect 29116 1935 29184 1959
rect 29116 1879 29122 1935
rect 29178 1879 29184 1935
rect 29116 1855 29184 1879
rect 29116 1799 29122 1855
rect 29178 1799 29184 1855
rect 29116 1775 29184 1799
rect 29116 1719 29122 1775
rect 29178 1719 29184 1775
rect 29116 1695 29184 1719
rect 29116 1639 29122 1695
rect 29178 1639 29184 1695
rect 29116 1615 29184 1639
rect 29116 1559 29122 1615
rect 29178 1559 29184 1615
rect 29116 1535 29184 1559
rect 29116 1479 29122 1535
rect 29178 1479 29184 1535
rect 29116 1455 29184 1479
rect 29116 1399 29122 1455
rect 29178 1399 29184 1455
rect 29116 1375 29184 1399
rect 29116 1319 29122 1375
rect 29178 1319 29184 1375
rect 29116 1295 29184 1319
rect 29116 1239 29122 1295
rect 29178 1239 29184 1295
rect 29116 1215 29184 1239
rect 29116 1159 29122 1215
rect 29178 1159 29184 1215
rect 29116 1147 29184 1159
rect 29308 3135 29376 3522
rect 29308 3079 29314 3135
rect 29370 3079 29376 3135
rect 29308 3055 29376 3079
rect 29308 2999 29314 3055
rect 29370 2999 29376 3055
rect 29308 2975 29376 2999
rect 29308 2919 29314 2975
rect 29370 2919 29376 2975
rect 29308 2895 29376 2919
rect 29308 2839 29314 2895
rect 29370 2839 29376 2895
rect 29308 2815 29376 2839
rect 29308 2759 29314 2815
rect 29370 2759 29376 2815
rect 29308 2735 29376 2759
rect 29308 2679 29314 2735
rect 29370 2679 29376 2735
rect 29308 2655 29376 2679
rect 29308 2599 29314 2655
rect 29370 2599 29376 2655
rect 29308 2575 29376 2599
rect 29308 2519 29314 2575
rect 29370 2519 29376 2575
rect 29308 2495 29376 2519
rect 29308 2439 29314 2495
rect 29370 2439 29376 2495
rect 29308 2415 29376 2439
rect 29308 2359 29314 2415
rect 29370 2359 29376 2415
rect 29308 2335 29376 2359
rect 29308 2279 29314 2335
rect 29370 2279 29376 2335
rect 29308 2255 29376 2279
rect 29308 2199 29314 2255
rect 29370 2199 29376 2255
rect 29308 2175 29376 2199
rect 29308 2119 29314 2175
rect 29370 2119 29376 2175
rect 29308 2095 29376 2119
rect 29308 2039 29314 2095
rect 29370 2039 29376 2095
rect 29308 2015 29376 2039
rect 29308 1959 29314 2015
rect 29370 1959 29376 2015
rect 29308 1935 29376 1959
rect 29308 1879 29314 1935
rect 29370 1879 29376 1935
rect 29308 1855 29376 1879
rect 29308 1799 29314 1855
rect 29370 1799 29376 1855
rect 29308 1775 29376 1799
rect 29308 1719 29314 1775
rect 29370 1719 29376 1775
rect 29308 1695 29376 1719
rect 29308 1639 29314 1695
rect 29370 1639 29376 1695
rect 29308 1615 29376 1639
rect 29308 1559 29314 1615
rect 29370 1559 29376 1615
rect 29308 1535 29376 1559
rect 29308 1479 29314 1535
rect 29370 1479 29376 1535
rect 29308 1455 29376 1479
rect 29308 1399 29314 1455
rect 29370 1399 29376 1455
rect 29308 1375 29376 1399
rect 29308 1319 29314 1375
rect 29370 1319 29376 1375
rect 29308 1295 29376 1319
rect 29308 1239 29314 1295
rect 29370 1239 29376 1295
rect 29308 1215 29376 1239
rect 29308 1159 29314 1215
rect 29370 1159 29376 1215
rect 29308 1147 29376 1159
rect 29500 3135 29568 3522
rect 29500 3079 29506 3135
rect 29562 3079 29568 3135
rect 29500 3055 29568 3079
rect 29500 2999 29506 3055
rect 29562 2999 29568 3055
rect 29500 2975 29568 2999
rect 29500 2919 29506 2975
rect 29562 2919 29568 2975
rect 29500 2895 29568 2919
rect 29500 2839 29506 2895
rect 29562 2839 29568 2895
rect 29500 2815 29568 2839
rect 29500 2759 29506 2815
rect 29562 2759 29568 2815
rect 29500 2735 29568 2759
rect 29500 2679 29506 2735
rect 29562 2679 29568 2735
rect 29500 2655 29568 2679
rect 29500 2599 29506 2655
rect 29562 2599 29568 2655
rect 29500 2575 29568 2599
rect 29500 2519 29506 2575
rect 29562 2519 29568 2575
rect 29500 2495 29568 2519
rect 29500 2439 29506 2495
rect 29562 2439 29568 2495
rect 29500 2415 29568 2439
rect 29500 2359 29506 2415
rect 29562 2359 29568 2415
rect 29500 2335 29568 2359
rect 29500 2279 29506 2335
rect 29562 2279 29568 2335
rect 29500 2255 29568 2279
rect 29500 2199 29506 2255
rect 29562 2199 29568 2255
rect 29500 2175 29568 2199
rect 29500 2119 29506 2175
rect 29562 2119 29568 2175
rect 29500 2095 29568 2119
rect 29500 2039 29506 2095
rect 29562 2039 29568 2095
rect 29500 2015 29568 2039
rect 29500 1959 29506 2015
rect 29562 1959 29568 2015
rect 29500 1935 29568 1959
rect 29500 1879 29506 1935
rect 29562 1879 29568 1935
rect 29500 1855 29568 1879
rect 29500 1799 29506 1855
rect 29562 1799 29568 1855
rect 29500 1775 29568 1799
rect 29500 1719 29506 1775
rect 29562 1719 29568 1775
rect 29500 1695 29568 1719
rect 29500 1639 29506 1695
rect 29562 1639 29568 1695
rect 29500 1615 29568 1639
rect 29500 1559 29506 1615
rect 29562 1559 29568 1615
rect 29500 1535 29568 1559
rect 29500 1479 29506 1535
rect 29562 1479 29568 1535
rect 29500 1455 29568 1479
rect 29500 1399 29506 1455
rect 29562 1399 29568 1455
rect 29500 1375 29568 1399
rect 29500 1319 29506 1375
rect 29562 1319 29568 1375
rect 29500 1295 29568 1319
rect 29500 1239 29506 1295
rect 29562 1239 29568 1295
rect 29500 1215 29568 1239
rect 29500 1159 29506 1215
rect 29562 1159 29568 1215
rect 29500 1147 29568 1159
rect 29692 3135 29760 3522
rect 29692 3079 29698 3135
rect 29754 3079 29760 3135
rect 29692 3055 29760 3079
rect 29692 2999 29698 3055
rect 29754 2999 29760 3055
rect 29692 2975 29760 2999
rect 29692 2919 29698 2975
rect 29754 2919 29760 2975
rect 29692 2895 29760 2919
rect 29692 2839 29698 2895
rect 29754 2839 29760 2895
rect 29692 2815 29760 2839
rect 29692 2759 29698 2815
rect 29754 2759 29760 2815
rect 29692 2735 29760 2759
rect 29692 2679 29698 2735
rect 29754 2679 29760 2735
rect 29692 2655 29760 2679
rect 29692 2599 29698 2655
rect 29754 2599 29760 2655
rect 29692 2575 29760 2599
rect 29692 2519 29698 2575
rect 29754 2519 29760 2575
rect 29692 2495 29760 2519
rect 29692 2439 29698 2495
rect 29754 2439 29760 2495
rect 29692 2415 29760 2439
rect 29692 2359 29698 2415
rect 29754 2359 29760 2415
rect 29692 2335 29760 2359
rect 29692 2279 29698 2335
rect 29754 2279 29760 2335
rect 29692 2255 29760 2279
rect 29692 2199 29698 2255
rect 29754 2199 29760 2255
rect 29692 2175 29760 2199
rect 29692 2119 29698 2175
rect 29754 2119 29760 2175
rect 29692 2095 29760 2119
rect 29692 2039 29698 2095
rect 29754 2039 29760 2095
rect 29692 2015 29760 2039
rect 29692 1959 29698 2015
rect 29754 1959 29760 2015
rect 29692 1935 29760 1959
rect 29692 1879 29698 1935
rect 29754 1879 29760 1935
rect 29692 1855 29760 1879
rect 29692 1799 29698 1855
rect 29754 1799 29760 1855
rect 29692 1775 29760 1799
rect 29692 1719 29698 1775
rect 29754 1719 29760 1775
rect 29692 1695 29760 1719
rect 29692 1639 29698 1695
rect 29754 1639 29760 1695
rect 29692 1615 29760 1639
rect 29692 1559 29698 1615
rect 29754 1559 29760 1615
rect 29692 1535 29760 1559
rect 29692 1479 29698 1535
rect 29754 1479 29760 1535
rect 29692 1455 29760 1479
rect 29692 1399 29698 1455
rect 29754 1399 29760 1455
rect 29692 1375 29760 1399
rect 29692 1319 29698 1375
rect 29754 1319 29760 1375
rect 29692 1295 29760 1319
rect 29692 1239 29698 1295
rect 29754 1239 29760 1295
rect 29692 1215 29760 1239
rect 29692 1159 29698 1215
rect 29754 1159 29760 1215
rect 29692 1147 29760 1159
rect 29884 3135 29952 3522
rect 29884 3079 29890 3135
rect 29946 3079 29952 3135
rect 29884 3055 29952 3079
rect 29884 2999 29890 3055
rect 29946 2999 29952 3055
rect 29884 2975 29952 2999
rect 29884 2919 29890 2975
rect 29946 2919 29952 2975
rect 29884 2895 29952 2919
rect 29884 2839 29890 2895
rect 29946 2839 29952 2895
rect 29884 2815 29952 2839
rect 29884 2759 29890 2815
rect 29946 2759 29952 2815
rect 29884 2735 29952 2759
rect 29884 2679 29890 2735
rect 29946 2679 29952 2735
rect 29884 2655 29952 2679
rect 29884 2599 29890 2655
rect 29946 2599 29952 2655
rect 29884 2575 29952 2599
rect 29884 2519 29890 2575
rect 29946 2519 29952 2575
rect 29884 2495 29952 2519
rect 29884 2439 29890 2495
rect 29946 2439 29952 2495
rect 29884 2415 29952 2439
rect 29884 2359 29890 2415
rect 29946 2359 29952 2415
rect 29884 2335 29952 2359
rect 29884 2279 29890 2335
rect 29946 2279 29952 2335
rect 29884 2255 29952 2279
rect 29884 2199 29890 2255
rect 29946 2199 29952 2255
rect 29884 2175 29952 2199
rect 29884 2119 29890 2175
rect 29946 2119 29952 2175
rect 29884 2095 29952 2119
rect 29884 2039 29890 2095
rect 29946 2039 29952 2095
rect 29884 2015 29952 2039
rect 29884 1959 29890 2015
rect 29946 1959 29952 2015
rect 29884 1935 29952 1959
rect 29884 1879 29890 1935
rect 29946 1879 29952 1935
rect 29884 1855 29952 1879
rect 29884 1799 29890 1855
rect 29946 1799 29952 1855
rect 29884 1775 29952 1799
rect 29884 1719 29890 1775
rect 29946 1719 29952 1775
rect 29884 1695 29952 1719
rect 29884 1639 29890 1695
rect 29946 1639 29952 1695
rect 29884 1615 29952 1639
rect 29884 1559 29890 1615
rect 29946 1559 29952 1615
rect 29884 1535 29952 1559
rect 29884 1479 29890 1535
rect 29946 1479 29952 1535
rect 29884 1455 29952 1479
rect 29884 1399 29890 1455
rect 29946 1399 29952 1455
rect 29884 1375 29952 1399
rect 29884 1319 29890 1375
rect 29946 1319 29952 1375
rect 29884 1295 29952 1319
rect 29884 1239 29890 1295
rect 29946 1239 29952 1295
rect 29884 1215 29952 1239
rect 29884 1159 29890 1215
rect 29946 1159 29952 1215
rect 29884 1147 29952 1159
rect 30076 3135 30144 3522
rect 30076 3079 30082 3135
rect 30138 3079 30144 3135
rect 30076 3055 30144 3079
rect 30076 2999 30082 3055
rect 30138 2999 30144 3055
rect 30076 2975 30144 2999
rect 30076 2919 30082 2975
rect 30138 2919 30144 2975
rect 30076 2895 30144 2919
rect 30076 2839 30082 2895
rect 30138 2839 30144 2895
rect 30076 2815 30144 2839
rect 30076 2759 30082 2815
rect 30138 2759 30144 2815
rect 30076 2735 30144 2759
rect 30076 2679 30082 2735
rect 30138 2679 30144 2735
rect 30076 2655 30144 2679
rect 30076 2599 30082 2655
rect 30138 2599 30144 2655
rect 30076 2575 30144 2599
rect 30076 2519 30082 2575
rect 30138 2519 30144 2575
rect 30076 2495 30144 2519
rect 30076 2439 30082 2495
rect 30138 2439 30144 2495
rect 30076 2415 30144 2439
rect 30076 2359 30082 2415
rect 30138 2359 30144 2415
rect 30076 2335 30144 2359
rect 30076 2279 30082 2335
rect 30138 2279 30144 2335
rect 30076 2255 30144 2279
rect 30076 2199 30082 2255
rect 30138 2199 30144 2255
rect 30076 2175 30144 2199
rect 30076 2119 30082 2175
rect 30138 2119 30144 2175
rect 30076 2095 30144 2119
rect 30076 2039 30082 2095
rect 30138 2039 30144 2095
rect 30076 2015 30144 2039
rect 30076 1959 30082 2015
rect 30138 1959 30144 2015
rect 30076 1935 30144 1959
rect 30076 1879 30082 1935
rect 30138 1879 30144 1935
rect 30076 1855 30144 1879
rect 30076 1799 30082 1855
rect 30138 1799 30144 1855
rect 30076 1775 30144 1799
rect 30076 1719 30082 1775
rect 30138 1719 30144 1775
rect 30076 1695 30144 1719
rect 30076 1639 30082 1695
rect 30138 1639 30144 1695
rect 30076 1615 30144 1639
rect 30076 1559 30082 1615
rect 30138 1559 30144 1615
rect 30076 1535 30144 1559
rect 30076 1479 30082 1535
rect 30138 1479 30144 1535
rect 30076 1455 30144 1479
rect 30076 1399 30082 1455
rect 30138 1399 30144 1455
rect 30076 1375 30144 1399
rect 30076 1319 30082 1375
rect 30138 1319 30144 1375
rect 30076 1295 30144 1319
rect 30076 1239 30082 1295
rect 30138 1239 30144 1295
rect 30076 1215 30144 1239
rect 30076 1159 30082 1215
rect 30138 1159 30144 1215
rect 30076 1147 30144 1159
rect 30268 3135 30336 3522
rect 30268 3079 30274 3135
rect 30330 3079 30336 3135
rect 30268 3055 30336 3079
rect 30268 2999 30274 3055
rect 30330 2999 30336 3055
rect 30268 2975 30336 2999
rect 30268 2919 30274 2975
rect 30330 2919 30336 2975
rect 30268 2895 30336 2919
rect 30268 2839 30274 2895
rect 30330 2839 30336 2895
rect 30268 2815 30336 2839
rect 30268 2759 30274 2815
rect 30330 2759 30336 2815
rect 30268 2735 30336 2759
rect 30268 2679 30274 2735
rect 30330 2679 30336 2735
rect 30268 2655 30336 2679
rect 30268 2599 30274 2655
rect 30330 2599 30336 2655
rect 30268 2575 30336 2599
rect 30268 2519 30274 2575
rect 30330 2519 30336 2575
rect 30268 2495 30336 2519
rect 30268 2439 30274 2495
rect 30330 2439 30336 2495
rect 30268 2415 30336 2439
rect 30268 2359 30274 2415
rect 30330 2359 30336 2415
rect 30268 2335 30336 2359
rect 30268 2279 30274 2335
rect 30330 2279 30336 2335
rect 30268 2255 30336 2279
rect 30268 2199 30274 2255
rect 30330 2199 30336 2255
rect 30268 2175 30336 2199
rect 30268 2119 30274 2175
rect 30330 2119 30336 2175
rect 30268 2095 30336 2119
rect 30268 2039 30274 2095
rect 30330 2039 30336 2095
rect 30268 2015 30336 2039
rect 30268 1959 30274 2015
rect 30330 1959 30336 2015
rect 30268 1935 30336 1959
rect 30268 1879 30274 1935
rect 30330 1879 30336 1935
rect 30268 1855 30336 1879
rect 30268 1799 30274 1855
rect 30330 1799 30336 1855
rect 30268 1775 30336 1799
rect 30268 1719 30274 1775
rect 30330 1719 30336 1775
rect 30268 1695 30336 1719
rect 30268 1639 30274 1695
rect 30330 1639 30336 1695
rect 30268 1615 30336 1639
rect 30268 1559 30274 1615
rect 30330 1559 30336 1615
rect 30268 1535 30336 1559
rect 30268 1479 30274 1535
rect 30330 1479 30336 1535
rect 30268 1455 30336 1479
rect 30268 1399 30274 1455
rect 30330 1399 30336 1455
rect 30268 1375 30336 1399
rect 30268 1319 30274 1375
rect 30330 1319 30336 1375
rect 30268 1295 30336 1319
rect 30268 1239 30274 1295
rect 30330 1239 30336 1295
rect 30268 1215 30336 1239
rect 30268 1159 30274 1215
rect 30330 1159 30336 1215
rect 30268 1147 30336 1159
rect 30460 3135 30528 3522
rect 30460 3079 30466 3135
rect 30522 3079 30528 3135
rect 30460 3055 30528 3079
rect 30460 2999 30466 3055
rect 30522 2999 30528 3055
rect 30460 2975 30528 2999
rect 30460 2919 30466 2975
rect 30522 2919 30528 2975
rect 30460 2895 30528 2919
rect 30460 2839 30466 2895
rect 30522 2839 30528 2895
rect 30460 2815 30528 2839
rect 30460 2759 30466 2815
rect 30522 2759 30528 2815
rect 30460 2735 30528 2759
rect 30460 2679 30466 2735
rect 30522 2679 30528 2735
rect 30460 2655 30528 2679
rect 30460 2599 30466 2655
rect 30522 2599 30528 2655
rect 30460 2575 30528 2599
rect 30460 2519 30466 2575
rect 30522 2519 30528 2575
rect 30460 2495 30528 2519
rect 30460 2439 30466 2495
rect 30522 2439 30528 2495
rect 30460 2415 30528 2439
rect 30460 2359 30466 2415
rect 30522 2359 30528 2415
rect 30460 2335 30528 2359
rect 30460 2279 30466 2335
rect 30522 2279 30528 2335
rect 30460 2255 30528 2279
rect 30460 2199 30466 2255
rect 30522 2199 30528 2255
rect 30460 2175 30528 2199
rect 30460 2119 30466 2175
rect 30522 2119 30528 2175
rect 30460 2095 30528 2119
rect 30460 2039 30466 2095
rect 30522 2039 30528 2095
rect 30460 2015 30528 2039
rect 30460 1959 30466 2015
rect 30522 1959 30528 2015
rect 30460 1935 30528 1959
rect 30460 1879 30466 1935
rect 30522 1879 30528 1935
rect 30460 1855 30528 1879
rect 30460 1799 30466 1855
rect 30522 1799 30528 1855
rect 30460 1775 30528 1799
rect 30460 1719 30466 1775
rect 30522 1719 30528 1775
rect 30460 1695 30528 1719
rect 30460 1639 30466 1695
rect 30522 1639 30528 1695
rect 30460 1615 30528 1639
rect 30460 1559 30466 1615
rect 30522 1559 30528 1615
rect 30460 1535 30528 1559
rect 30460 1479 30466 1535
rect 30522 1479 30528 1535
rect 30460 1455 30528 1479
rect 30460 1399 30466 1455
rect 30522 1399 30528 1455
rect 30460 1375 30528 1399
rect 30460 1319 30466 1375
rect 30522 1319 30528 1375
rect 30460 1295 30528 1319
rect 30460 1239 30466 1295
rect 30522 1239 30528 1295
rect 30460 1215 30528 1239
rect 30460 1159 30466 1215
rect 30522 1159 30528 1215
rect 30460 1147 30528 1159
rect 30652 3135 30720 3522
rect 30652 3079 30658 3135
rect 30714 3079 30720 3135
rect 30652 3055 30720 3079
rect 30652 2999 30658 3055
rect 30714 2999 30720 3055
rect 30652 2975 30720 2999
rect 30652 2919 30658 2975
rect 30714 2919 30720 2975
rect 30652 2895 30720 2919
rect 30652 2839 30658 2895
rect 30714 2839 30720 2895
rect 30652 2815 30720 2839
rect 30652 2759 30658 2815
rect 30714 2759 30720 2815
rect 30652 2735 30720 2759
rect 30652 2679 30658 2735
rect 30714 2679 30720 2735
rect 30652 2655 30720 2679
rect 30652 2599 30658 2655
rect 30714 2599 30720 2655
rect 30652 2575 30720 2599
rect 30652 2519 30658 2575
rect 30714 2519 30720 2575
rect 30652 2495 30720 2519
rect 30652 2439 30658 2495
rect 30714 2439 30720 2495
rect 30652 2415 30720 2439
rect 30652 2359 30658 2415
rect 30714 2359 30720 2415
rect 30652 2335 30720 2359
rect 30652 2279 30658 2335
rect 30714 2279 30720 2335
rect 30652 2255 30720 2279
rect 30652 2199 30658 2255
rect 30714 2199 30720 2255
rect 30652 2175 30720 2199
rect 30652 2119 30658 2175
rect 30714 2119 30720 2175
rect 30652 2095 30720 2119
rect 30652 2039 30658 2095
rect 30714 2039 30720 2095
rect 30652 2015 30720 2039
rect 30652 1959 30658 2015
rect 30714 1959 30720 2015
rect 30652 1935 30720 1959
rect 30652 1879 30658 1935
rect 30714 1879 30720 1935
rect 30652 1855 30720 1879
rect 30652 1799 30658 1855
rect 30714 1799 30720 1855
rect 30652 1775 30720 1799
rect 30652 1719 30658 1775
rect 30714 1719 30720 1775
rect 30652 1695 30720 1719
rect 30652 1639 30658 1695
rect 30714 1639 30720 1695
rect 30652 1615 30720 1639
rect 30652 1559 30658 1615
rect 30714 1559 30720 1615
rect 30652 1535 30720 1559
rect 30652 1479 30658 1535
rect 30714 1479 30720 1535
rect 30652 1455 30720 1479
rect 30652 1399 30658 1455
rect 30714 1399 30720 1455
rect 30652 1375 30720 1399
rect 30652 1319 30658 1375
rect 30714 1319 30720 1375
rect 30652 1295 30720 1319
rect 30652 1239 30658 1295
rect 30714 1239 30720 1295
rect 30652 1215 30720 1239
rect 30652 1159 30658 1215
rect 30714 1159 30720 1215
rect 30652 1147 30720 1159
rect 30844 3135 30912 3522
rect 30844 3079 30850 3135
rect 30906 3079 30912 3135
rect 30844 3055 30912 3079
rect 30844 2999 30850 3055
rect 30906 2999 30912 3055
rect 30844 2975 30912 2999
rect 30844 2919 30850 2975
rect 30906 2919 30912 2975
rect 30844 2895 30912 2919
rect 30844 2839 30850 2895
rect 30906 2839 30912 2895
rect 30844 2815 30912 2839
rect 30844 2759 30850 2815
rect 30906 2759 30912 2815
rect 30844 2735 30912 2759
rect 30844 2679 30850 2735
rect 30906 2679 30912 2735
rect 30844 2655 30912 2679
rect 30844 2599 30850 2655
rect 30906 2599 30912 2655
rect 30844 2575 30912 2599
rect 30844 2519 30850 2575
rect 30906 2519 30912 2575
rect 30844 2495 30912 2519
rect 30844 2439 30850 2495
rect 30906 2439 30912 2495
rect 30844 2415 30912 2439
rect 30844 2359 30850 2415
rect 30906 2359 30912 2415
rect 30844 2335 30912 2359
rect 30844 2279 30850 2335
rect 30906 2279 30912 2335
rect 30844 2255 30912 2279
rect 30844 2199 30850 2255
rect 30906 2199 30912 2255
rect 30844 2175 30912 2199
rect 30844 2119 30850 2175
rect 30906 2119 30912 2175
rect 30844 2095 30912 2119
rect 30844 2039 30850 2095
rect 30906 2039 30912 2095
rect 30844 2015 30912 2039
rect 30844 1959 30850 2015
rect 30906 1959 30912 2015
rect 30844 1935 30912 1959
rect 30844 1879 30850 1935
rect 30906 1879 30912 1935
rect 30844 1855 30912 1879
rect 30844 1799 30850 1855
rect 30906 1799 30912 1855
rect 30844 1775 30912 1799
rect 30844 1719 30850 1775
rect 30906 1719 30912 1775
rect 30844 1695 30912 1719
rect 30844 1639 30850 1695
rect 30906 1639 30912 1695
rect 30844 1615 30912 1639
rect 30844 1559 30850 1615
rect 30906 1559 30912 1615
rect 30844 1535 30912 1559
rect 30844 1479 30850 1535
rect 30906 1479 30912 1535
rect 30844 1455 30912 1479
rect 30844 1399 30850 1455
rect 30906 1399 30912 1455
rect 30844 1375 30912 1399
rect 30844 1319 30850 1375
rect 30906 1319 30912 1375
rect 30844 1295 30912 1319
rect 30844 1239 30850 1295
rect 30906 1239 30912 1295
rect 30844 1215 30912 1239
rect 30844 1159 30850 1215
rect 30906 1159 30912 1215
rect 30844 1147 30912 1159
rect 31036 3135 31104 3522
rect 31036 3079 31042 3135
rect 31098 3079 31104 3135
rect 31036 3055 31104 3079
rect 31036 2999 31042 3055
rect 31098 2999 31104 3055
rect 31036 2975 31104 2999
rect 31036 2919 31042 2975
rect 31098 2919 31104 2975
rect 31036 2895 31104 2919
rect 31036 2839 31042 2895
rect 31098 2839 31104 2895
rect 31036 2815 31104 2839
rect 31036 2759 31042 2815
rect 31098 2759 31104 2815
rect 31036 2735 31104 2759
rect 31036 2679 31042 2735
rect 31098 2679 31104 2735
rect 31036 2655 31104 2679
rect 31036 2599 31042 2655
rect 31098 2599 31104 2655
rect 31036 2575 31104 2599
rect 31036 2519 31042 2575
rect 31098 2519 31104 2575
rect 31036 2495 31104 2519
rect 31036 2439 31042 2495
rect 31098 2439 31104 2495
rect 31036 2415 31104 2439
rect 31036 2359 31042 2415
rect 31098 2359 31104 2415
rect 31036 2335 31104 2359
rect 31036 2279 31042 2335
rect 31098 2279 31104 2335
rect 31036 2255 31104 2279
rect 31036 2199 31042 2255
rect 31098 2199 31104 2255
rect 31036 2175 31104 2199
rect 31036 2119 31042 2175
rect 31098 2119 31104 2175
rect 31036 2095 31104 2119
rect 31036 2039 31042 2095
rect 31098 2039 31104 2095
rect 31036 2015 31104 2039
rect 31036 1959 31042 2015
rect 31098 1959 31104 2015
rect 31036 1935 31104 1959
rect 31036 1879 31042 1935
rect 31098 1879 31104 1935
rect 31036 1855 31104 1879
rect 31036 1799 31042 1855
rect 31098 1799 31104 1855
rect 31036 1775 31104 1799
rect 31036 1719 31042 1775
rect 31098 1719 31104 1775
rect 31036 1695 31104 1719
rect 31036 1639 31042 1695
rect 31098 1639 31104 1695
rect 31036 1615 31104 1639
rect 31036 1559 31042 1615
rect 31098 1559 31104 1615
rect 31036 1535 31104 1559
rect 31036 1479 31042 1535
rect 31098 1479 31104 1535
rect 31036 1455 31104 1479
rect 31036 1399 31042 1455
rect 31098 1399 31104 1455
rect 31036 1375 31104 1399
rect 31036 1319 31042 1375
rect 31098 1319 31104 1375
rect 31036 1295 31104 1319
rect 31036 1239 31042 1295
rect 31098 1239 31104 1295
rect 31036 1215 31104 1239
rect 31036 1159 31042 1215
rect 31098 1159 31104 1215
rect 31036 1147 31104 1159
rect 31228 3135 31296 3522
rect 31228 3079 31234 3135
rect 31290 3079 31296 3135
rect 31228 3055 31296 3079
rect 31228 2999 31234 3055
rect 31290 2999 31296 3055
rect 31228 2975 31296 2999
rect 31228 2919 31234 2975
rect 31290 2919 31296 2975
rect 31228 2895 31296 2919
rect 31228 2839 31234 2895
rect 31290 2839 31296 2895
rect 31228 2815 31296 2839
rect 31228 2759 31234 2815
rect 31290 2759 31296 2815
rect 31228 2735 31296 2759
rect 31228 2679 31234 2735
rect 31290 2679 31296 2735
rect 31228 2655 31296 2679
rect 31228 2599 31234 2655
rect 31290 2599 31296 2655
rect 31228 2575 31296 2599
rect 31228 2519 31234 2575
rect 31290 2519 31296 2575
rect 31228 2495 31296 2519
rect 31228 2439 31234 2495
rect 31290 2439 31296 2495
rect 31228 2415 31296 2439
rect 31228 2359 31234 2415
rect 31290 2359 31296 2415
rect 31228 2335 31296 2359
rect 31228 2279 31234 2335
rect 31290 2279 31296 2335
rect 31228 2255 31296 2279
rect 31228 2199 31234 2255
rect 31290 2199 31296 2255
rect 31228 2175 31296 2199
rect 31228 2119 31234 2175
rect 31290 2119 31296 2175
rect 31228 2095 31296 2119
rect 31228 2039 31234 2095
rect 31290 2039 31296 2095
rect 31228 2015 31296 2039
rect 31228 1959 31234 2015
rect 31290 1959 31296 2015
rect 31228 1935 31296 1959
rect 31228 1879 31234 1935
rect 31290 1879 31296 1935
rect 31228 1855 31296 1879
rect 31228 1799 31234 1855
rect 31290 1799 31296 1855
rect 31228 1775 31296 1799
rect 31228 1719 31234 1775
rect 31290 1719 31296 1775
rect 31228 1695 31296 1719
rect 31228 1639 31234 1695
rect 31290 1639 31296 1695
rect 31228 1615 31296 1639
rect 31228 1559 31234 1615
rect 31290 1559 31296 1615
rect 31228 1535 31296 1559
rect 31228 1479 31234 1535
rect 31290 1479 31296 1535
rect 31228 1455 31296 1479
rect 31228 1399 31234 1455
rect 31290 1399 31296 1455
rect 31228 1375 31296 1399
rect 31228 1319 31234 1375
rect 31290 1319 31296 1375
rect 31228 1295 31296 1319
rect 31228 1239 31234 1295
rect 31290 1239 31296 1295
rect 31228 1215 31296 1239
rect 31228 1159 31234 1215
rect 31290 1159 31296 1215
rect 31228 1147 31296 1159
rect 31420 3135 31488 3522
rect 31420 3079 31426 3135
rect 31482 3079 31488 3135
rect 31420 3055 31488 3079
rect 31420 2999 31426 3055
rect 31482 2999 31488 3055
rect 31420 2975 31488 2999
rect 31420 2919 31426 2975
rect 31482 2919 31488 2975
rect 31420 2895 31488 2919
rect 31420 2839 31426 2895
rect 31482 2839 31488 2895
rect 31420 2815 31488 2839
rect 31420 2759 31426 2815
rect 31482 2759 31488 2815
rect 31420 2735 31488 2759
rect 31420 2679 31426 2735
rect 31482 2679 31488 2735
rect 31420 2655 31488 2679
rect 31420 2599 31426 2655
rect 31482 2599 31488 2655
rect 31420 2575 31488 2599
rect 31420 2519 31426 2575
rect 31482 2519 31488 2575
rect 31420 2495 31488 2519
rect 31420 2439 31426 2495
rect 31482 2439 31488 2495
rect 31420 2415 31488 2439
rect 31420 2359 31426 2415
rect 31482 2359 31488 2415
rect 31420 2335 31488 2359
rect 31420 2279 31426 2335
rect 31482 2279 31488 2335
rect 31420 2255 31488 2279
rect 31420 2199 31426 2255
rect 31482 2199 31488 2255
rect 31420 2175 31488 2199
rect 31420 2119 31426 2175
rect 31482 2119 31488 2175
rect 31420 2095 31488 2119
rect 31420 2039 31426 2095
rect 31482 2039 31488 2095
rect 31420 2015 31488 2039
rect 31420 1959 31426 2015
rect 31482 1959 31488 2015
rect 31420 1935 31488 1959
rect 31420 1879 31426 1935
rect 31482 1879 31488 1935
rect 31420 1855 31488 1879
rect 31420 1799 31426 1855
rect 31482 1799 31488 1855
rect 31420 1775 31488 1799
rect 31420 1719 31426 1775
rect 31482 1719 31488 1775
rect 31420 1695 31488 1719
rect 31420 1639 31426 1695
rect 31482 1639 31488 1695
rect 31420 1615 31488 1639
rect 31420 1559 31426 1615
rect 31482 1559 31488 1615
rect 31420 1535 31488 1559
rect 31420 1479 31426 1535
rect 31482 1479 31488 1535
rect 31420 1455 31488 1479
rect 31420 1399 31426 1455
rect 31482 1399 31488 1455
rect 31420 1375 31488 1399
rect 31420 1319 31426 1375
rect 31482 1319 31488 1375
rect 31420 1295 31488 1319
rect 31420 1239 31426 1295
rect 31482 1239 31488 1295
rect 31420 1215 31488 1239
rect 31420 1159 31426 1215
rect 31482 1159 31488 1215
rect 31420 1147 31488 1159
rect 31612 3135 31680 3522
rect 31612 3079 31618 3135
rect 31674 3079 31680 3135
rect 31612 3055 31680 3079
rect 31612 2999 31618 3055
rect 31674 2999 31680 3055
rect 31612 2975 31680 2999
rect 31612 2919 31618 2975
rect 31674 2919 31680 2975
rect 31612 2895 31680 2919
rect 31612 2839 31618 2895
rect 31674 2839 31680 2895
rect 31612 2815 31680 2839
rect 31612 2759 31618 2815
rect 31674 2759 31680 2815
rect 31612 2735 31680 2759
rect 31612 2679 31618 2735
rect 31674 2679 31680 2735
rect 31612 2655 31680 2679
rect 31612 2599 31618 2655
rect 31674 2599 31680 2655
rect 31612 2575 31680 2599
rect 31612 2519 31618 2575
rect 31674 2519 31680 2575
rect 31612 2495 31680 2519
rect 31612 2439 31618 2495
rect 31674 2439 31680 2495
rect 31612 2415 31680 2439
rect 31612 2359 31618 2415
rect 31674 2359 31680 2415
rect 31612 2335 31680 2359
rect 31612 2279 31618 2335
rect 31674 2279 31680 2335
rect 31612 2255 31680 2279
rect 31612 2199 31618 2255
rect 31674 2199 31680 2255
rect 31612 2175 31680 2199
rect 31612 2119 31618 2175
rect 31674 2119 31680 2175
rect 31612 2095 31680 2119
rect 31612 2039 31618 2095
rect 31674 2039 31680 2095
rect 31612 2015 31680 2039
rect 31612 1959 31618 2015
rect 31674 1959 31680 2015
rect 31612 1935 31680 1959
rect 31612 1879 31618 1935
rect 31674 1879 31680 1935
rect 31612 1855 31680 1879
rect 31612 1799 31618 1855
rect 31674 1799 31680 1855
rect 31612 1775 31680 1799
rect 31612 1719 31618 1775
rect 31674 1719 31680 1775
rect 31612 1695 31680 1719
rect 31612 1639 31618 1695
rect 31674 1639 31680 1695
rect 31612 1615 31680 1639
rect 31612 1559 31618 1615
rect 31674 1559 31680 1615
rect 31612 1535 31680 1559
rect 31612 1479 31618 1535
rect 31674 1479 31680 1535
rect 31612 1455 31680 1479
rect 31612 1399 31618 1455
rect 31674 1399 31680 1455
rect 31612 1375 31680 1399
rect 31612 1319 31618 1375
rect 31674 1319 31680 1375
rect 31612 1295 31680 1319
rect 31612 1239 31618 1295
rect 31674 1239 31680 1295
rect 31612 1215 31680 1239
rect 31612 1159 31618 1215
rect 31674 1159 31680 1215
rect 31612 1147 31680 1159
rect 31804 3135 31872 3522
rect 31804 3079 31810 3135
rect 31866 3079 31872 3135
rect 31804 3055 31872 3079
rect 31804 2999 31810 3055
rect 31866 2999 31872 3055
rect 31804 2975 31872 2999
rect 31804 2919 31810 2975
rect 31866 2919 31872 2975
rect 31804 2895 31872 2919
rect 31804 2839 31810 2895
rect 31866 2839 31872 2895
rect 31804 2815 31872 2839
rect 31804 2759 31810 2815
rect 31866 2759 31872 2815
rect 31804 2735 31872 2759
rect 31804 2679 31810 2735
rect 31866 2679 31872 2735
rect 31804 2655 31872 2679
rect 31804 2599 31810 2655
rect 31866 2599 31872 2655
rect 31804 2575 31872 2599
rect 31804 2519 31810 2575
rect 31866 2519 31872 2575
rect 31804 2495 31872 2519
rect 31804 2439 31810 2495
rect 31866 2439 31872 2495
rect 31804 2415 31872 2439
rect 31804 2359 31810 2415
rect 31866 2359 31872 2415
rect 31804 2335 31872 2359
rect 31804 2279 31810 2335
rect 31866 2279 31872 2335
rect 31804 2255 31872 2279
rect 31804 2199 31810 2255
rect 31866 2199 31872 2255
rect 31804 2175 31872 2199
rect 31804 2119 31810 2175
rect 31866 2119 31872 2175
rect 31804 2095 31872 2119
rect 31804 2039 31810 2095
rect 31866 2039 31872 2095
rect 31804 2015 31872 2039
rect 31804 1959 31810 2015
rect 31866 1959 31872 2015
rect 31804 1935 31872 1959
rect 31804 1879 31810 1935
rect 31866 1879 31872 1935
rect 31804 1855 31872 1879
rect 31804 1799 31810 1855
rect 31866 1799 31872 1855
rect 31804 1775 31872 1799
rect 31804 1719 31810 1775
rect 31866 1719 31872 1775
rect 31804 1695 31872 1719
rect 31804 1639 31810 1695
rect 31866 1639 31872 1695
rect 31804 1615 31872 1639
rect 31804 1559 31810 1615
rect 31866 1559 31872 1615
rect 31804 1535 31872 1559
rect 31804 1479 31810 1535
rect 31866 1479 31872 1535
rect 31804 1455 31872 1479
rect 31804 1399 31810 1455
rect 31866 1399 31872 1455
rect 31804 1375 31872 1399
rect 31804 1319 31810 1375
rect 31866 1319 31872 1375
rect 31804 1295 31872 1319
rect 31804 1239 31810 1295
rect 31866 1239 31872 1295
rect 31804 1215 31872 1239
rect 31804 1159 31810 1215
rect 31866 1159 31872 1215
rect 31804 1147 31872 1159
rect 31996 3135 32064 3522
rect 31996 3079 32002 3135
rect 32058 3079 32064 3135
rect 31996 3055 32064 3079
rect 31996 2999 32002 3055
rect 32058 2999 32064 3055
rect 31996 2975 32064 2999
rect 31996 2919 32002 2975
rect 32058 2919 32064 2975
rect 31996 2895 32064 2919
rect 31996 2839 32002 2895
rect 32058 2839 32064 2895
rect 31996 2815 32064 2839
rect 31996 2759 32002 2815
rect 32058 2759 32064 2815
rect 31996 2735 32064 2759
rect 31996 2679 32002 2735
rect 32058 2679 32064 2735
rect 31996 2655 32064 2679
rect 31996 2599 32002 2655
rect 32058 2599 32064 2655
rect 31996 2575 32064 2599
rect 31996 2519 32002 2575
rect 32058 2519 32064 2575
rect 31996 2495 32064 2519
rect 31996 2439 32002 2495
rect 32058 2439 32064 2495
rect 31996 2415 32064 2439
rect 31996 2359 32002 2415
rect 32058 2359 32064 2415
rect 31996 2335 32064 2359
rect 31996 2279 32002 2335
rect 32058 2279 32064 2335
rect 31996 2255 32064 2279
rect 31996 2199 32002 2255
rect 32058 2199 32064 2255
rect 31996 2175 32064 2199
rect 31996 2119 32002 2175
rect 32058 2119 32064 2175
rect 31996 2095 32064 2119
rect 31996 2039 32002 2095
rect 32058 2039 32064 2095
rect 31996 2015 32064 2039
rect 31996 1959 32002 2015
rect 32058 1959 32064 2015
rect 31996 1935 32064 1959
rect 31996 1879 32002 1935
rect 32058 1879 32064 1935
rect 31996 1855 32064 1879
rect 31996 1799 32002 1855
rect 32058 1799 32064 1855
rect 31996 1775 32064 1799
rect 31996 1719 32002 1775
rect 32058 1719 32064 1775
rect 31996 1695 32064 1719
rect 31996 1639 32002 1695
rect 32058 1639 32064 1695
rect 31996 1615 32064 1639
rect 31996 1559 32002 1615
rect 32058 1559 32064 1615
rect 31996 1535 32064 1559
rect 31996 1479 32002 1535
rect 32058 1479 32064 1535
rect 31996 1455 32064 1479
rect 31996 1399 32002 1455
rect 32058 1399 32064 1455
rect 31996 1375 32064 1399
rect 31996 1319 32002 1375
rect 32058 1319 32064 1375
rect 31996 1295 32064 1319
rect 31996 1239 32002 1295
rect 32058 1239 32064 1295
rect 31996 1215 32064 1239
rect 31996 1159 32002 1215
rect 32058 1159 32064 1215
rect 31996 1147 32064 1159
rect 32188 3135 32256 3522
rect 32188 3079 32194 3135
rect 32250 3079 32256 3135
rect 32188 3055 32256 3079
rect 32188 2999 32194 3055
rect 32250 2999 32256 3055
rect 32188 2975 32256 2999
rect 32188 2919 32194 2975
rect 32250 2919 32256 2975
rect 32188 2895 32256 2919
rect 32188 2839 32194 2895
rect 32250 2839 32256 2895
rect 32188 2815 32256 2839
rect 32188 2759 32194 2815
rect 32250 2759 32256 2815
rect 32188 2735 32256 2759
rect 32188 2679 32194 2735
rect 32250 2679 32256 2735
rect 32188 2655 32256 2679
rect 32188 2599 32194 2655
rect 32250 2599 32256 2655
rect 32188 2575 32256 2599
rect 32188 2519 32194 2575
rect 32250 2519 32256 2575
rect 32188 2495 32256 2519
rect 32188 2439 32194 2495
rect 32250 2439 32256 2495
rect 32188 2415 32256 2439
rect 32188 2359 32194 2415
rect 32250 2359 32256 2415
rect 32188 2335 32256 2359
rect 32188 2279 32194 2335
rect 32250 2279 32256 2335
rect 32188 2255 32256 2279
rect 32188 2199 32194 2255
rect 32250 2199 32256 2255
rect 32188 2175 32256 2199
rect 32188 2119 32194 2175
rect 32250 2119 32256 2175
rect 32188 2095 32256 2119
rect 32188 2039 32194 2095
rect 32250 2039 32256 2095
rect 32188 2015 32256 2039
rect 32188 1959 32194 2015
rect 32250 1959 32256 2015
rect 32188 1935 32256 1959
rect 32188 1879 32194 1935
rect 32250 1879 32256 1935
rect 32188 1855 32256 1879
rect 32188 1799 32194 1855
rect 32250 1799 32256 1855
rect 32188 1775 32256 1799
rect 32188 1719 32194 1775
rect 32250 1719 32256 1775
rect 32188 1695 32256 1719
rect 32188 1639 32194 1695
rect 32250 1639 32256 1695
rect 32188 1615 32256 1639
rect 32188 1559 32194 1615
rect 32250 1559 32256 1615
rect 32188 1535 32256 1559
rect 32188 1479 32194 1535
rect 32250 1479 32256 1535
rect 32188 1455 32256 1479
rect 32188 1399 32194 1455
rect 32250 1399 32256 1455
rect 32188 1375 32256 1399
rect 32188 1319 32194 1375
rect 32250 1319 32256 1375
rect 32188 1295 32256 1319
rect 32188 1239 32194 1295
rect 32250 1239 32256 1295
rect 32188 1215 32256 1239
rect 32188 1159 32194 1215
rect 32250 1159 32256 1215
rect 32188 1147 32256 1159
rect 32380 3135 32448 3522
rect 32380 3079 32386 3135
rect 32442 3079 32448 3135
rect 32380 3055 32448 3079
rect 32380 2999 32386 3055
rect 32442 2999 32448 3055
rect 32380 2975 32448 2999
rect 32380 2919 32386 2975
rect 32442 2919 32448 2975
rect 32380 2895 32448 2919
rect 32380 2839 32386 2895
rect 32442 2839 32448 2895
rect 32380 2815 32448 2839
rect 32380 2759 32386 2815
rect 32442 2759 32448 2815
rect 32380 2735 32448 2759
rect 32380 2679 32386 2735
rect 32442 2679 32448 2735
rect 32380 2655 32448 2679
rect 32380 2599 32386 2655
rect 32442 2599 32448 2655
rect 32380 2575 32448 2599
rect 32380 2519 32386 2575
rect 32442 2519 32448 2575
rect 32380 2495 32448 2519
rect 32380 2439 32386 2495
rect 32442 2439 32448 2495
rect 32380 2415 32448 2439
rect 32380 2359 32386 2415
rect 32442 2359 32448 2415
rect 32380 2335 32448 2359
rect 32380 2279 32386 2335
rect 32442 2279 32448 2335
rect 32380 2255 32448 2279
rect 32380 2199 32386 2255
rect 32442 2199 32448 2255
rect 32380 2175 32448 2199
rect 32380 2119 32386 2175
rect 32442 2119 32448 2175
rect 32380 2095 32448 2119
rect 32380 2039 32386 2095
rect 32442 2039 32448 2095
rect 32380 2015 32448 2039
rect 32380 1959 32386 2015
rect 32442 1959 32448 2015
rect 32380 1935 32448 1959
rect 32380 1879 32386 1935
rect 32442 1879 32448 1935
rect 32380 1855 32448 1879
rect 32380 1799 32386 1855
rect 32442 1799 32448 1855
rect 32380 1775 32448 1799
rect 32380 1719 32386 1775
rect 32442 1719 32448 1775
rect 32380 1695 32448 1719
rect 32380 1639 32386 1695
rect 32442 1639 32448 1695
rect 32380 1615 32448 1639
rect 32380 1559 32386 1615
rect 32442 1559 32448 1615
rect 32380 1535 32448 1559
rect 32380 1479 32386 1535
rect 32442 1479 32448 1535
rect 32380 1455 32448 1479
rect 32380 1399 32386 1455
rect 32442 1399 32448 1455
rect 32380 1375 32448 1399
rect 32380 1319 32386 1375
rect 32442 1319 32448 1375
rect 32380 1295 32448 1319
rect 32380 1239 32386 1295
rect 32442 1239 32448 1295
rect 32380 1215 32448 1239
rect 32380 1159 32386 1215
rect 32442 1159 32448 1215
rect 32380 1147 32448 1159
rect 32572 3135 32640 3522
rect 32572 3079 32578 3135
rect 32634 3079 32640 3135
rect 32572 3055 32640 3079
rect 32572 2999 32578 3055
rect 32634 2999 32640 3055
rect 32572 2975 32640 2999
rect 32572 2919 32578 2975
rect 32634 2919 32640 2975
rect 32572 2895 32640 2919
rect 32572 2839 32578 2895
rect 32634 2839 32640 2895
rect 32572 2815 32640 2839
rect 32572 2759 32578 2815
rect 32634 2759 32640 2815
rect 32572 2735 32640 2759
rect 32572 2679 32578 2735
rect 32634 2679 32640 2735
rect 32572 2655 32640 2679
rect 32572 2599 32578 2655
rect 32634 2599 32640 2655
rect 32572 2575 32640 2599
rect 32572 2519 32578 2575
rect 32634 2519 32640 2575
rect 32572 2495 32640 2519
rect 32572 2439 32578 2495
rect 32634 2439 32640 2495
rect 32572 2415 32640 2439
rect 32572 2359 32578 2415
rect 32634 2359 32640 2415
rect 32572 2335 32640 2359
rect 32572 2279 32578 2335
rect 32634 2279 32640 2335
rect 32572 2255 32640 2279
rect 32572 2199 32578 2255
rect 32634 2199 32640 2255
rect 32572 2175 32640 2199
rect 32572 2119 32578 2175
rect 32634 2119 32640 2175
rect 32572 2095 32640 2119
rect 32572 2039 32578 2095
rect 32634 2039 32640 2095
rect 32572 2015 32640 2039
rect 32572 1959 32578 2015
rect 32634 1959 32640 2015
rect 32572 1935 32640 1959
rect 32572 1879 32578 1935
rect 32634 1879 32640 1935
rect 32572 1855 32640 1879
rect 32572 1799 32578 1855
rect 32634 1799 32640 1855
rect 32572 1775 32640 1799
rect 32572 1719 32578 1775
rect 32634 1719 32640 1775
rect 32572 1695 32640 1719
rect 32572 1639 32578 1695
rect 32634 1639 32640 1695
rect 32572 1615 32640 1639
rect 32572 1559 32578 1615
rect 32634 1559 32640 1615
rect 32572 1535 32640 1559
rect 32572 1479 32578 1535
rect 32634 1479 32640 1535
rect 32572 1455 32640 1479
rect 32572 1399 32578 1455
rect 32634 1399 32640 1455
rect 32572 1375 32640 1399
rect 32572 1319 32578 1375
rect 32634 1319 32640 1375
rect 32572 1295 32640 1319
rect 32572 1239 32578 1295
rect 32634 1239 32640 1295
rect 32572 1215 32640 1239
rect 32572 1159 32578 1215
rect 32634 1159 32640 1215
rect 32572 1147 32640 1159
rect 32764 3135 32832 3522
rect 32764 3079 32770 3135
rect 32826 3079 32832 3135
rect 32764 3055 32832 3079
rect 32764 2999 32770 3055
rect 32826 2999 32832 3055
rect 32764 2975 32832 2999
rect 32764 2919 32770 2975
rect 32826 2919 32832 2975
rect 32764 2895 32832 2919
rect 32764 2839 32770 2895
rect 32826 2839 32832 2895
rect 32764 2815 32832 2839
rect 32764 2759 32770 2815
rect 32826 2759 32832 2815
rect 32764 2735 32832 2759
rect 32764 2679 32770 2735
rect 32826 2679 32832 2735
rect 32764 2655 32832 2679
rect 32764 2599 32770 2655
rect 32826 2599 32832 2655
rect 32764 2575 32832 2599
rect 32764 2519 32770 2575
rect 32826 2519 32832 2575
rect 32764 2495 32832 2519
rect 32764 2439 32770 2495
rect 32826 2439 32832 2495
rect 32764 2415 32832 2439
rect 32764 2359 32770 2415
rect 32826 2359 32832 2415
rect 32764 2335 32832 2359
rect 32764 2279 32770 2335
rect 32826 2279 32832 2335
rect 32764 2255 32832 2279
rect 32764 2199 32770 2255
rect 32826 2199 32832 2255
rect 32764 2175 32832 2199
rect 32764 2119 32770 2175
rect 32826 2119 32832 2175
rect 32764 2095 32832 2119
rect 32764 2039 32770 2095
rect 32826 2039 32832 2095
rect 32764 2015 32832 2039
rect 32764 1959 32770 2015
rect 32826 1959 32832 2015
rect 32764 1935 32832 1959
rect 32764 1879 32770 1935
rect 32826 1879 32832 1935
rect 32764 1855 32832 1879
rect 32764 1799 32770 1855
rect 32826 1799 32832 1855
rect 32764 1775 32832 1799
rect 32764 1719 32770 1775
rect 32826 1719 32832 1775
rect 32764 1695 32832 1719
rect 32764 1639 32770 1695
rect 32826 1639 32832 1695
rect 32764 1615 32832 1639
rect 32764 1559 32770 1615
rect 32826 1559 32832 1615
rect 32764 1535 32832 1559
rect 32764 1479 32770 1535
rect 32826 1479 32832 1535
rect 32764 1455 32832 1479
rect 32764 1399 32770 1455
rect 32826 1399 32832 1455
rect 32764 1375 32832 1399
rect 32764 1319 32770 1375
rect 32826 1319 32832 1375
rect 32764 1295 32832 1319
rect 32764 1239 32770 1295
rect 32826 1239 32832 1295
rect 32764 1215 32832 1239
rect 32764 1159 32770 1215
rect 32826 1159 32832 1215
rect 32764 1147 32832 1159
rect 32956 3135 33024 3522
rect 32956 3079 32962 3135
rect 33018 3079 33024 3135
rect 32956 3055 33024 3079
rect 32956 2999 32962 3055
rect 33018 2999 33024 3055
rect 32956 2975 33024 2999
rect 32956 2919 32962 2975
rect 33018 2919 33024 2975
rect 32956 2895 33024 2919
rect 32956 2839 32962 2895
rect 33018 2839 33024 2895
rect 32956 2815 33024 2839
rect 32956 2759 32962 2815
rect 33018 2759 33024 2815
rect 32956 2735 33024 2759
rect 32956 2679 32962 2735
rect 33018 2679 33024 2735
rect 32956 2655 33024 2679
rect 32956 2599 32962 2655
rect 33018 2599 33024 2655
rect 32956 2575 33024 2599
rect 32956 2519 32962 2575
rect 33018 2519 33024 2575
rect 32956 2495 33024 2519
rect 32956 2439 32962 2495
rect 33018 2439 33024 2495
rect 32956 2415 33024 2439
rect 32956 2359 32962 2415
rect 33018 2359 33024 2415
rect 32956 2335 33024 2359
rect 32956 2279 32962 2335
rect 33018 2279 33024 2335
rect 32956 2255 33024 2279
rect 32956 2199 32962 2255
rect 33018 2199 33024 2255
rect 32956 2175 33024 2199
rect 32956 2119 32962 2175
rect 33018 2119 33024 2175
rect 32956 2095 33024 2119
rect 32956 2039 32962 2095
rect 33018 2039 33024 2095
rect 32956 2015 33024 2039
rect 32956 1959 32962 2015
rect 33018 1959 33024 2015
rect 32956 1935 33024 1959
rect 32956 1879 32962 1935
rect 33018 1879 33024 1935
rect 32956 1855 33024 1879
rect 32956 1799 32962 1855
rect 33018 1799 33024 1855
rect 32956 1775 33024 1799
rect 32956 1719 32962 1775
rect 33018 1719 33024 1775
rect 32956 1695 33024 1719
rect 32956 1639 32962 1695
rect 33018 1639 33024 1695
rect 32956 1615 33024 1639
rect 32956 1559 32962 1615
rect 33018 1559 33024 1615
rect 32956 1535 33024 1559
rect 32956 1479 32962 1535
rect 33018 1479 33024 1535
rect 32956 1455 33024 1479
rect 32956 1399 32962 1455
rect 33018 1399 33024 1455
rect 32956 1375 33024 1399
rect 32956 1319 32962 1375
rect 33018 1319 33024 1375
rect 32956 1295 33024 1319
rect 32956 1239 32962 1295
rect 33018 1239 33024 1295
rect 32956 1215 33024 1239
rect 32956 1159 32962 1215
rect 33018 1159 33024 1215
rect 32956 1147 33024 1159
rect 33148 3135 33216 3522
rect 33148 3079 33154 3135
rect 33210 3079 33216 3135
rect 33148 3055 33216 3079
rect 33148 2999 33154 3055
rect 33210 2999 33216 3055
rect 33148 2975 33216 2999
rect 33148 2919 33154 2975
rect 33210 2919 33216 2975
rect 33148 2895 33216 2919
rect 33148 2839 33154 2895
rect 33210 2839 33216 2895
rect 33148 2815 33216 2839
rect 33148 2759 33154 2815
rect 33210 2759 33216 2815
rect 33148 2735 33216 2759
rect 33148 2679 33154 2735
rect 33210 2679 33216 2735
rect 33148 2655 33216 2679
rect 33148 2599 33154 2655
rect 33210 2599 33216 2655
rect 33148 2575 33216 2599
rect 33148 2519 33154 2575
rect 33210 2519 33216 2575
rect 33148 2495 33216 2519
rect 33148 2439 33154 2495
rect 33210 2439 33216 2495
rect 33148 2415 33216 2439
rect 33148 2359 33154 2415
rect 33210 2359 33216 2415
rect 33148 2335 33216 2359
rect 33148 2279 33154 2335
rect 33210 2279 33216 2335
rect 33148 2255 33216 2279
rect 33148 2199 33154 2255
rect 33210 2199 33216 2255
rect 33148 2175 33216 2199
rect 33148 2119 33154 2175
rect 33210 2119 33216 2175
rect 33148 2095 33216 2119
rect 33148 2039 33154 2095
rect 33210 2039 33216 2095
rect 33148 2015 33216 2039
rect 33148 1959 33154 2015
rect 33210 1959 33216 2015
rect 33148 1935 33216 1959
rect 33148 1879 33154 1935
rect 33210 1879 33216 1935
rect 33148 1855 33216 1879
rect 33148 1799 33154 1855
rect 33210 1799 33216 1855
rect 33148 1775 33216 1799
rect 33148 1719 33154 1775
rect 33210 1719 33216 1775
rect 33148 1695 33216 1719
rect 33148 1639 33154 1695
rect 33210 1639 33216 1695
rect 33148 1615 33216 1639
rect 33148 1559 33154 1615
rect 33210 1559 33216 1615
rect 33148 1535 33216 1559
rect 33148 1479 33154 1535
rect 33210 1479 33216 1535
rect 33148 1455 33216 1479
rect 33148 1399 33154 1455
rect 33210 1399 33216 1455
rect 33148 1375 33216 1399
rect 33148 1319 33154 1375
rect 33210 1319 33216 1375
rect 33148 1295 33216 1319
rect 33148 1239 33154 1295
rect 33210 1239 33216 1295
rect 33148 1215 33216 1239
rect 33148 1159 33154 1215
rect 33210 1159 33216 1215
rect 33148 1147 33216 1159
rect 33340 3135 33408 3522
rect 33340 3079 33346 3135
rect 33402 3079 33408 3135
rect 33340 3055 33408 3079
rect 33340 2999 33346 3055
rect 33402 2999 33408 3055
rect 33340 2975 33408 2999
rect 33340 2919 33346 2975
rect 33402 2919 33408 2975
rect 33340 2895 33408 2919
rect 33340 2839 33346 2895
rect 33402 2839 33408 2895
rect 33340 2815 33408 2839
rect 33340 2759 33346 2815
rect 33402 2759 33408 2815
rect 33340 2735 33408 2759
rect 33340 2679 33346 2735
rect 33402 2679 33408 2735
rect 33340 2655 33408 2679
rect 33340 2599 33346 2655
rect 33402 2599 33408 2655
rect 33340 2575 33408 2599
rect 33340 2519 33346 2575
rect 33402 2519 33408 2575
rect 33340 2495 33408 2519
rect 33340 2439 33346 2495
rect 33402 2439 33408 2495
rect 33340 2415 33408 2439
rect 33340 2359 33346 2415
rect 33402 2359 33408 2415
rect 33340 2335 33408 2359
rect 33340 2279 33346 2335
rect 33402 2279 33408 2335
rect 33340 2255 33408 2279
rect 33340 2199 33346 2255
rect 33402 2199 33408 2255
rect 33340 2175 33408 2199
rect 33340 2119 33346 2175
rect 33402 2119 33408 2175
rect 33340 2095 33408 2119
rect 33340 2039 33346 2095
rect 33402 2039 33408 2095
rect 33340 2015 33408 2039
rect 33340 1959 33346 2015
rect 33402 1959 33408 2015
rect 33340 1935 33408 1959
rect 33340 1879 33346 1935
rect 33402 1879 33408 1935
rect 33340 1855 33408 1879
rect 33340 1799 33346 1855
rect 33402 1799 33408 1855
rect 33340 1775 33408 1799
rect 33340 1719 33346 1775
rect 33402 1719 33408 1775
rect 33340 1695 33408 1719
rect 33340 1639 33346 1695
rect 33402 1639 33408 1695
rect 33340 1615 33408 1639
rect 33340 1559 33346 1615
rect 33402 1559 33408 1615
rect 33340 1535 33408 1559
rect 33340 1479 33346 1535
rect 33402 1479 33408 1535
rect 33340 1455 33408 1479
rect 33340 1399 33346 1455
rect 33402 1399 33408 1455
rect 33340 1375 33408 1399
rect 33340 1319 33346 1375
rect 33402 1319 33408 1375
rect 33340 1295 33408 1319
rect 33340 1239 33346 1295
rect 33402 1239 33408 1295
rect 33340 1215 33408 1239
rect 33340 1159 33346 1215
rect 33402 1159 33408 1215
rect 33340 1147 33408 1159
rect 33532 3135 33600 3522
rect 33532 3079 33538 3135
rect 33594 3079 33600 3135
rect 33532 3055 33600 3079
rect 33532 2999 33538 3055
rect 33594 2999 33600 3055
rect 33532 2975 33600 2999
rect 33532 2919 33538 2975
rect 33594 2919 33600 2975
rect 33532 2895 33600 2919
rect 33532 2839 33538 2895
rect 33594 2839 33600 2895
rect 33532 2815 33600 2839
rect 33532 2759 33538 2815
rect 33594 2759 33600 2815
rect 33532 2735 33600 2759
rect 33532 2679 33538 2735
rect 33594 2679 33600 2735
rect 33532 2655 33600 2679
rect 33532 2599 33538 2655
rect 33594 2599 33600 2655
rect 33532 2575 33600 2599
rect 33532 2519 33538 2575
rect 33594 2519 33600 2575
rect 33532 2495 33600 2519
rect 33532 2439 33538 2495
rect 33594 2439 33600 2495
rect 33532 2415 33600 2439
rect 33532 2359 33538 2415
rect 33594 2359 33600 2415
rect 33532 2335 33600 2359
rect 33532 2279 33538 2335
rect 33594 2279 33600 2335
rect 33532 2255 33600 2279
rect 33532 2199 33538 2255
rect 33594 2199 33600 2255
rect 33532 2175 33600 2199
rect 33532 2119 33538 2175
rect 33594 2119 33600 2175
rect 33532 2095 33600 2119
rect 33532 2039 33538 2095
rect 33594 2039 33600 2095
rect 33532 2015 33600 2039
rect 33532 1959 33538 2015
rect 33594 1959 33600 2015
rect 33532 1935 33600 1959
rect 33532 1879 33538 1935
rect 33594 1879 33600 1935
rect 33532 1855 33600 1879
rect 33532 1799 33538 1855
rect 33594 1799 33600 1855
rect 33532 1775 33600 1799
rect 33532 1719 33538 1775
rect 33594 1719 33600 1775
rect 33532 1695 33600 1719
rect 33532 1639 33538 1695
rect 33594 1639 33600 1695
rect 33532 1615 33600 1639
rect 33532 1559 33538 1615
rect 33594 1559 33600 1615
rect 33532 1535 33600 1559
rect 33532 1479 33538 1535
rect 33594 1479 33600 1535
rect 33532 1455 33600 1479
rect 33532 1399 33538 1455
rect 33594 1399 33600 1455
rect 33532 1375 33600 1399
rect 33532 1319 33538 1375
rect 33594 1319 33600 1375
rect 33532 1295 33600 1319
rect 33532 1239 33538 1295
rect 33594 1239 33600 1295
rect 33532 1215 33600 1239
rect 33532 1159 33538 1215
rect 33594 1159 33600 1215
rect 33532 1147 33600 1159
rect 33724 3135 33792 3522
rect 33724 3079 33730 3135
rect 33786 3079 33792 3135
rect 33724 3055 33792 3079
rect 33724 2999 33730 3055
rect 33786 2999 33792 3055
rect 33724 2975 33792 2999
rect 33724 2919 33730 2975
rect 33786 2919 33792 2975
rect 33724 2895 33792 2919
rect 33724 2839 33730 2895
rect 33786 2839 33792 2895
rect 33724 2815 33792 2839
rect 33724 2759 33730 2815
rect 33786 2759 33792 2815
rect 33724 2735 33792 2759
rect 33724 2679 33730 2735
rect 33786 2679 33792 2735
rect 33724 2655 33792 2679
rect 33724 2599 33730 2655
rect 33786 2599 33792 2655
rect 33724 2575 33792 2599
rect 33724 2519 33730 2575
rect 33786 2519 33792 2575
rect 33724 2495 33792 2519
rect 33724 2439 33730 2495
rect 33786 2439 33792 2495
rect 33724 2415 33792 2439
rect 33724 2359 33730 2415
rect 33786 2359 33792 2415
rect 33724 2335 33792 2359
rect 33724 2279 33730 2335
rect 33786 2279 33792 2335
rect 33724 2255 33792 2279
rect 33724 2199 33730 2255
rect 33786 2199 33792 2255
rect 33724 2175 33792 2199
rect 33724 2119 33730 2175
rect 33786 2119 33792 2175
rect 33724 2095 33792 2119
rect 33724 2039 33730 2095
rect 33786 2039 33792 2095
rect 33724 2015 33792 2039
rect 33724 1959 33730 2015
rect 33786 1959 33792 2015
rect 33724 1935 33792 1959
rect 33724 1879 33730 1935
rect 33786 1879 33792 1935
rect 33724 1855 33792 1879
rect 33724 1799 33730 1855
rect 33786 1799 33792 1855
rect 33724 1775 33792 1799
rect 33724 1719 33730 1775
rect 33786 1719 33792 1775
rect 33724 1695 33792 1719
rect 33724 1639 33730 1695
rect 33786 1639 33792 1695
rect 33724 1615 33792 1639
rect 33724 1559 33730 1615
rect 33786 1559 33792 1615
rect 33724 1535 33792 1559
rect 33724 1479 33730 1535
rect 33786 1479 33792 1535
rect 33724 1455 33792 1479
rect 33724 1399 33730 1455
rect 33786 1399 33792 1455
rect 33724 1375 33792 1399
rect 33724 1319 33730 1375
rect 33786 1319 33792 1375
rect 33724 1295 33792 1319
rect 33724 1239 33730 1295
rect 33786 1239 33792 1295
rect 33724 1215 33792 1239
rect 33724 1159 33730 1215
rect 33786 1159 33792 1215
rect 33724 1147 33792 1159
rect 33916 3135 33984 3522
rect 33916 3079 33922 3135
rect 33978 3079 33984 3135
rect 33916 3055 33984 3079
rect 33916 2999 33922 3055
rect 33978 2999 33984 3055
rect 33916 2975 33984 2999
rect 33916 2919 33922 2975
rect 33978 2919 33984 2975
rect 33916 2895 33984 2919
rect 33916 2839 33922 2895
rect 33978 2839 33984 2895
rect 33916 2815 33984 2839
rect 33916 2759 33922 2815
rect 33978 2759 33984 2815
rect 33916 2735 33984 2759
rect 33916 2679 33922 2735
rect 33978 2679 33984 2735
rect 33916 2655 33984 2679
rect 33916 2599 33922 2655
rect 33978 2599 33984 2655
rect 33916 2575 33984 2599
rect 33916 2519 33922 2575
rect 33978 2519 33984 2575
rect 33916 2495 33984 2519
rect 33916 2439 33922 2495
rect 33978 2439 33984 2495
rect 33916 2415 33984 2439
rect 33916 2359 33922 2415
rect 33978 2359 33984 2415
rect 33916 2335 33984 2359
rect 33916 2279 33922 2335
rect 33978 2279 33984 2335
rect 33916 2255 33984 2279
rect 33916 2199 33922 2255
rect 33978 2199 33984 2255
rect 33916 2175 33984 2199
rect 33916 2119 33922 2175
rect 33978 2119 33984 2175
rect 33916 2095 33984 2119
rect 33916 2039 33922 2095
rect 33978 2039 33984 2095
rect 33916 2015 33984 2039
rect 33916 1959 33922 2015
rect 33978 1959 33984 2015
rect 33916 1935 33984 1959
rect 33916 1879 33922 1935
rect 33978 1879 33984 1935
rect 33916 1855 33984 1879
rect 33916 1799 33922 1855
rect 33978 1799 33984 1855
rect 33916 1775 33984 1799
rect 33916 1719 33922 1775
rect 33978 1719 33984 1775
rect 33916 1695 33984 1719
rect 33916 1639 33922 1695
rect 33978 1639 33984 1695
rect 33916 1615 33984 1639
rect 33916 1559 33922 1615
rect 33978 1559 33984 1615
rect 33916 1535 33984 1559
rect 33916 1479 33922 1535
rect 33978 1479 33984 1535
rect 33916 1455 33984 1479
rect 33916 1399 33922 1455
rect 33978 1399 33984 1455
rect 33916 1375 33984 1399
rect 33916 1319 33922 1375
rect 33978 1319 33984 1375
rect 33916 1295 33984 1319
rect 33916 1239 33922 1295
rect 33978 1239 33984 1295
rect 33916 1215 33984 1239
rect 33916 1159 33922 1215
rect 33978 1159 33984 1215
rect 33916 1147 33984 1159
rect 34108 3135 34176 3522
rect 34108 3079 34114 3135
rect 34170 3079 34176 3135
rect 34108 3055 34176 3079
rect 34108 2999 34114 3055
rect 34170 2999 34176 3055
rect 34108 2975 34176 2999
rect 34108 2919 34114 2975
rect 34170 2919 34176 2975
rect 34108 2895 34176 2919
rect 34108 2839 34114 2895
rect 34170 2839 34176 2895
rect 34108 2815 34176 2839
rect 34108 2759 34114 2815
rect 34170 2759 34176 2815
rect 34108 2735 34176 2759
rect 34108 2679 34114 2735
rect 34170 2679 34176 2735
rect 34108 2655 34176 2679
rect 34108 2599 34114 2655
rect 34170 2599 34176 2655
rect 34108 2575 34176 2599
rect 34108 2519 34114 2575
rect 34170 2519 34176 2575
rect 34108 2495 34176 2519
rect 34108 2439 34114 2495
rect 34170 2439 34176 2495
rect 34108 2415 34176 2439
rect 34108 2359 34114 2415
rect 34170 2359 34176 2415
rect 34108 2335 34176 2359
rect 34108 2279 34114 2335
rect 34170 2279 34176 2335
rect 34108 2255 34176 2279
rect 34108 2199 34114 2255
rect 34170 2199 34176 2255
rect 34108 2175 34176 2199
rect 34108 2119 34114 2175
rect 34170 2119 34176 2175
rect 34108 2095 34176 2119
rect 34108 2039 34114 2095
rect 34170 2039 34176 2095
rect 34108 2015 34176 2039
rect 34108 1959 34114 2015
rect 34170 1959 34176 2015
rect 34108 1935 34176 1959
rect 34108 1879 34114 1935
rect 34170 1879 34176 1935
rect 34108 1855 34176 1879
rect 34108 1799 34114 1855
rect 34170 1799 34176 1855
rect 34108 1775 34176 1799
rect 34108 1719 34114 1775
rect 34170 1719 34176 1775
rect 34108 1695 34176 1719
rect 34108 1639 34114 1695
rect 34170 1639 34176 1695
rect 34108 1615 34176 1639
rect 34108 1559 34114 1615
rect 34170 1559 34176 1615
rect 34108 1535 34176 1559
rect 34108 1479 34114 1535
rect 34170 1479 34176 1535
rect 34108 1455 34176 1479
rect 34108 1399 34114 1455
rect 34170 1399 34176 1455
rect 34108 1375 34176 1399
rect 34108 1319 34114 1375
rect 34170 1319 34176 1375
rect 34108 1295 34176 1319
rect 34108 1239 34114 1295
rect 34170 1239 34176 1295
rect 34108 1215 34176 1239
rect 34108 1159 34114 1215
rect 34170 1159 34176 1215
rect 34108 1147 34176 1159
rect 34300 3135 34368 3522
rect 34300 3079 34306 3135
rect 34362 3079 34368 3135
rect 34300 3055 34368 3079
rect 34300 2999 34306 3055
rect 34362 2999 34368 3055
rect 34300 2975 34368 2999
rect 34300 2919 34306 2975
rect 34362 2919 34368 2975
rect 34300 2895 34368 2919
rect 34300 2839 34306 2895
rect 34362 2839 34368 2895
rect 34300 2815 34368 2839
rect 34300 2759 34306 2815
rect 34362 2759 34368 2815
rect 34300 2735 34368 2759
rect 34300 2679 34306 2735
rect 34362 2679 34368 2735
rect 34300 2655 34368 2679
rect 34300 2599 34306 2655
rect 34362 2599 34368 2655
rect 34300 2575 34368 2599
rect 34300 2519 34306 2575
rect 34362 2519 34368 2575
rect 34300 2495 34368 2519
rect 34300 2439 34306 2495
rect 34362 2439 34368 2495
rect 34300 2415 34368 2439
rect 34300 2359 34306 2415
rect 34362 2359 34368 2415
rect 34300 2335 34368 2359
rect 34300 2279 34306 2335
rect 34362 2279 34368 2335
rect 34300 2255 34368 2279
rect 34300 2199 34306 2255
rect 34362 2199 34368 2255
rect 34300 2175 34368 2199
rect 34300 2119 34306 2175
rect 34362 2119 34368 2175
rect 34300 2095 34368 2119
rect 34300 2039 34306 2095
rect 34362 2039 34368 2095
rect 34300 2015 34368 2039
rect 34300 1959 34306 2015
rect 34362 1959 34368 2015
rect 34300 1935 34368 1959
rect 34300 1879 34306 1935
rect 34362 1879 34368 1935
rect 34300 1855 34368 1879
rect 34300 1799 34306 1855
rect 34362 1799 34368 1855
rect 34300 1775 34368 1799
rect 34300 1719 34306 1775
rect 34362 1719 34368 1775
rect 34300 1695 34368 1719
rect 34300 1639 34306 1695
rect 34362 1639 34368 1695
rect 34300 1615 34368 1639
rect 34300 1559 34306 1615
rect 34362 1559 34368 1615
rect 34300 1535 34368 1559
rect 34300 1479 34306 1535
rect 34362 1479 34368 1535
rect 34300 1455 34368 1479
rect 34300 1399 34306 1455
rect 34362 1399 34368 1455
rect 34300 1375 34368 1399
rect 34300 1319 34306 1375
rect 34362 1319 34368 1375
rect 34300 1295 34368 1319
rect 34300 1239 34306 1295
rect 34362 1239 34368 1295
rect 34300 1215 34368 1239
rect 34300 1159 34306 1215
rect 34362 1159 34368 1215
rect 34300 1147 34368 1159
rect 34492 3135 34560 3522
rect 34492 3079 34498 3135
rect 34554 3079 34560 3135
rect 34492 3055 34560 3079
rect 34492 2999 34498 3055
rect 34554 2999 34560 3055
rect 34492 2975 34560 2999
rect 34492 2919 34498 2975
rect 34554 2919 34560 2975
rect 34492 2895 34560 2919
rect 34492 2839 34498 2895
rect 34554 2839 34560 2895
rect 34492 2815 34560 2839
rect 34492 2759 34498 2815
rect 34554 2759 34560 2815
rect 34492 2735 34560 2759
rect 34492 2679 34498 2735
rect 34554 2679 34560 2735
rect 34492 2655 34560 2679
rect 34492 2599 34498 2655
rect 34554 2599 34560 2655
rect 34492 2575 34560 2599
rect 34492 2519 34498 2575
rect 34554 2519 34560 2575
rect 34492 2495 34560 2519
rect 34492 2439 34498 2495
rect 34554 2439 34560 2495
rect 34492 2415 34560 2439
rect 34492 2359 34498 2415
rect 34554 2359 34560 2415
rect 34492 2335 34560 2359
rect 34492 2279 34498 2335
rect 34554 2279 34560 2335
rect 34492 2255 34560 2279
rect 34492 2199 34498 2255
rect 34554 2199 34560 2255
rect 34492 2175 34560 2199
rect 34492 2119 34498 2175
rect 34554 2119 34560 2175
rect 34492 2095 34560 2119
rect 34492 2039 34498 2095
rect 34554 2039 34560 2095
rect 34492 2015 34560 2039
rect 34492 1959 34498 2015
rect 34554 1959 34560 2015
rect 34492 1935 34560 1959
rect 34492 1879 34498 1935
rect 34554 1879 34560 1935
rect 34492 1855 34560 1879
rect 34492 1799 34498 1855
rect 34554 1799 34560 1855
rect 34492 1775 34560 1799
rect 34492 1719 34498 1775
rect 34554 1719 34560 1775
rect 34492 1695 34560 1719
rect 34492 1639 34498 1695
rect 34554 1639 34560 1695
rect 34492 1615 34560 1639
rect 34492 1559 34498 1615
rect 34554 1559 34560 1615
rect 34492 1535 34560 1559
rect 34492 1479 34498 1535
rect 34554 1479 34560 1535
rect 34492 1455 34560 1479
rect 34492 1399 34498 1455
rect 34554 1399 34560 1455
rect 34492 1375 34560 1399
rect 34492 1319 34498 1375
rect 34554 1319 34560 1375
rect 34492 1295 34560 1319
rect 34492 1239 34498 1295
rect 34554 1239 34560 1295
rect 34492 1215 34560 1239
rect 34492 1159 34498 1215
rect 34554 1159 34560 1215
rect 34492 1147 34560 1159
rect 34684 3135 34752 3522
rect 34684 3079 34690 3135
rect 34746 3079 34752 3135
rect 34684 3055 34752 3079
rect 34684 2999 34690 3055
rect 34746 2999 34752 3055
rect 34684 2975 34752 2999
rect 34684 2919 34690 2975
rect 34746 2919 34752 2975
rect 34684 2895 34752 2919
rect 34684 2839 34690 2895
rect 34746 2839 34752 2895
rect 34684 2815 34752 2839
rect 34684 2759 34690 2815
rect 34746 2759 34752 2815
rect 34684 2735 34752 2759
rect 34684 2679 34690 2735
rect 34746 2679 34752 2735
rect 34684 2655 34752 2679
rect 34684 2599 34690 2655
rect 34746 2599 34752 2655
rect 34684 2575 34752 2599
rect 34684 2519 34690 2575
rect 34746 2519 34752 2575
rect 34684 2495 34752 2519
rect 34684 2439 34690 2495
rect 34746 2439 34752 2495
rect 34684 2415 34752 2439
rect 34684 2359 34690 2415
rect 34746 2359 34752 2415
rect 34684 2335 34752 2359
rect 34684 2279 34690 2335
rect 34746 2279 34752 2335
rect 34684 2255 34752 2279
rect 34684 2199 34690 2255
rect 34746 2199 34752 2255
rect 34684 2175 34752 2199
rect 34684 2119 34690 2175
rect 34746 2119 34752 2175
rect 34684 2095 34752 2119
rect 34684 2039 34690 2095
rect 34746 2039 34752 2095
rect 34684 2015 34752 2039
rect 34684 1959 34690 2015
rect 34746 1959 34752 2015
rect 34684 1935 34752 1959
rect 34684 1879 34690 1935
rect 34746 1879 34752 1935
rect 34684 1855 34752 1879
rect 34684 1799 34690 1855
rect 34746 1799 34752 1855
rect 34684 1775 34752 1799
rect 34684 1719 34690 1775
rect 34746 1719 34752 1775
rect 34684 1695 34752 1719
rect 34684 1639 34690 1695
rect 34746 1639 34752 1695
rect 34684 1615 34752 1639
rect 34684 1559 34690 1615
rect 34746 1559 34752 1615
rect 34684 1535 34752 1559
rect 34684 1479 34690 1535
rect 34746 1479 34752 1535
rect 34684 1455 34752 1479
rect 34684 1399 34690 1455
rect 34746 1399 34752 1455
rect 34684 1375 34752 1399
rect 34684 1319 34690 1375
rect 34746 1319 34752 1375
rect 34684 1295 34752 1319
rect 34684 1239 34690 1295
rect 34746 1239 34752 1295
rect 34684 1215 34752 1239
rect 34684 1159 34690 1215
rect 34746 1159 34752 1215
rect 34684 1147 34752 1159
rect 34876 3135 34944 3522
rect 34876 3079 34882 3135
rect 34938 3079 34944 3135
rect 34876 3055 34944 3079
rect 34876 2999 34882 3055
rect 34938 2999 34944 3055
rect 34876 2975 34944 2999
rect 34876 2919 34882 2975
rect 34938 2919 34944 2975
rect 34876 2895 34944 2919
rect 34876 2839 34882 2895
rect 34938 2839 34944 2895
rect 34876 2815 34944 2839
rect 34876 2759 34882 2815
rect 34938 2759 34944 2815
rect 34876 2735 34944 2759
rect 34876 2679 34882 2735
rect 34938 2679 34944 2735
rect 34876 2655 34944 2679
rect 34876 2599 34882 2655
rect 34938 2599 34944 2655
rect 34876 2575 34944 2599
rect 34876 2519 34882 2575
rect 34938 2519 34944 2575
rect 34876 2495 34944 2519
rect 34876 2439 34882 2495
rect 34938 2439 34944 2495
rect 34876 2415 34944 2439
rect 34876 2359 34882 2415
rect 34938 2359 34944 2415
rect 34876 2335 34944 2359
rect 34876 2279 34882 2335
rect 34938 2279 34944 2335
rect 34876 2255 34944 2279
rect 34876 2199 34882 2255
rect 34938 2199 34944 2255
rect 34876 2175 34944 2199
rect 34876 2119 34882 2175
rect 34938 2119 34944 2175
rect 34876 2095 34944 2119
rect 34876 2039 34882 2095
rect 34938 2039 34944 2095
rect 34876 2015 34944 2039
rect 34876 1959 34882 2015
rect 34938 1959 34944 2015
rect 34876 1935 34944 1959
rect 34876 1879 34882 1935
rect 34938 1879 34944 1935
rect 34876 1855 34944 1879
rect 34876 1799 34882 1855
rect 34938 1799 34944 1855
rect 34876 1775 34944 1799
rect 34876 1719 34882 1775
rect 34938 1719 34944 1775
rect 34876 1695 34944 1719
rect 34876 1639 34882 1695
rect 34938 1639 34944 1695
rect 34876 1615 34944 1639
rect 34876 1559 34882 1615
rect 34938 1559 34944 1615
rect 34876 1535 34944 1559
rect 34876 1479 34882 1535
rect 34938 1479 34944 1535
rect 34876 1455 34944 1479
rect 34876 1399 34882 1455
rect 34938 1399 34944 1455
rect 34876 1375 34944 1399
rect 34876 1319 34882 1375
rect 34938 1319 34944 1375
rect 34876 1295 34944 1319
rect 34876 1239 34882 1295
rect 34938 1239 34944 1295
rect 34876 1215 34944 1239
rect 34876 1159 34882 1215
rect 34938 1159 34944 1215
rect 34876 1147 34944 1159
rect 35068 3135 35136 3522
rect 35068 3079 35074 3135
rect 35130 3079 35136 3135
rect 35068 3055 35136 3079
rect 35068 2999 35074 3055
rect 35130 2999 35136 3055
rect 35068 2975 35136 2999
rect 35068 2919 35074 2975
rect 35130 2919 35136 2975
rect 35068 2895 35136 2919
rect 35068 2839 35074 2895
rect 35130 2839 35136 2895
rect 35068 2815 35136 2839
rect 35068 2759 35074 2815
rect 35130 2759 35136 2815
rect 35068 2735 35136 2759
rect 35068 2679 35074 2735
rect 35130 2679 35136 2735
rect 35068 2655 35136 2679
rect 35068 2599 35074 2655
rect 35130 2599 35136 2655
rect 35068 2575 35136 2599
rect 35068 2519 35074 2575
rect 35130 2519 35136 2575
rect 35068 2495 35136 2519
rect 35068 2439 35074 2495
rect 35130 2439 35136 2495
rect 35068 2415 35136 2439
rect 35068 2359 35074 2415
rect 35130 2359 35136 2415
rect 35068 2335 35136 2359
rect 35068 2279 35074 2335
rect 35130 2279 35136 2335
rect 35068 2255 35136 2279
rect 35068 2199 35074 2255
rect 35130 2199 35136 2255
rect 35068 2175 35136 2199
rect 35068 2119 35074 2175
rect 35130 2119 35136 2175
rect 35068 2095 35136 2119
rect 35068 2039 35074 2095
rect 35130 2039 35136 2095
rect 35068 2015 35136 2039
rect 35068 1959 35074 2015
rect 35130 1959 35136 2015
rect 35068 1935 35136 1959
rect 35068 1879 35074 1935
rect 35130 1879 35136 1935
rect 35068 1855 35136 1879
rect 35068 1799 35074 1855
rect 35130 1799 35136 1855
rect 35068 1775 35136 1799
rect 35068 1719 35074 1775
rect 35130 1719 35136 1775
rect 35068 1695 35136 1719
rect 35068 1639 35074 1695
rect 35130 1639 35136 1695
rect 35068 1615 35136 1639
rect 35068 1559 35074 1615
rect 35130 1559 35136 1615
rect 35068 1535 35136 1559
rect 35068 1479 35074 1535
rect 35130 1479 35136 1535
rect 35068 1455 35136 1479
rect 35068 1399 35074 1455
rect 35130 1399 35136 1455
rect 35068 1375 35136 1399
rect 35068 1319 35074 1375
rect 35130 1319 35136 1375
rect 35068 1295 35136 1319
rect 35068 1239 35074 1295
rect 35130 1239 35136 1295
rect 35068 1215 35136 1239
rect 35068 1159 35074 1215
rect 35130 1159 35136 1215
rect 35068 1147 35136 1159
rect 35260 3135 35328 3522
rect 35260 3079 35266 3135
rect 35322 3079 35328 3135
rect 35260 3055 35328 3079
rect 35260 2999 35266 3055
rect 35322 2999 35328 3055
rect 35260 2975 35328 2999
rect 35260 2919 35266 2975
rect 35322 2919 35328 2975
rect 35260 2895 35328 2919
rect 35260 2839 35266 2895
rect 35322 2839 35328 2895
rect 35260 2815 35328 2839
rect 35260 2759 35266 2815
rect 35322 2759 35328 2815
rect 35260 2735 35328 2759
rect 35260 2679 35266 2735
rect 35322 2679 35328 2735
rect 35260 2655 35328 2679
rect 35260 2599 35266 2655
rect 35322 2599 35328 2655
rect 35260 2575 35328 2599
rect 35260 2519 35266 2575
rect 35322 2519 35328 2575
rect 35260 2495 35328 2519
rect 35260 2439 35266 2495
rect 35322 2439 35328 2495
rect 35260 2415 35328 2439
rect 35260 2359 35266 2415
rect 35322 2359 35328 2415
rect 35260 2335 35328 2359
rect 35260 2279 35266 2335
rect 35322 2279 35328 2335
rect 35260 2255 35328 2279
rect 35260 2199 35266 2255
rect 35322 2199 35328 2255
rect 35260 2175 35328 2199
rect 35260 2119 35266 2175
rect 35322 2119 35328 2175
rect 35260 2095 35328 2119
rect 35260 2039 35266 2095
rect 35322 2039 35328 2095
rect 35260 2015 35328 2039
rect 35260 1959 35266 2015
rect 35322 1959 35328 2015
rect 35260 1935 35328 1959
rect 35260 1879 35266 1935
rect 35322 1879 35328 1935
rect 35260 1855 35328 1879
rect 35260 1799 35266 1855
rect 35322 1799 35328 1855
rect 35260 1775 35328 1799
rect 35260 1719 35266 1775
rect 35322 1719 35328 1775
rect 35260 1695 35328 1719
rect 35260 1639 35266 1695
rect 35322 1639 35328 1695
rect 35260 1615 35328 1639
rect 35260 1559 35266 1615
rect 35322 1559 35328 1615
rect 35260 1535 35328 1559
rect 35260 1479 35266 1535
rect 35322 1479 35328 1535
rect 35260 1455 35328 1479
rect 35260 1399 35266 1455
rect 35322 1399 35328 1455
rect 35260 1375 35328 1399
rect 35260 1319 35266 1375
rect 35322 1319 35328 1375
rect 35260 1295 35328 1319
rect 35260 1239 35266 1295
rect 35322 1239 35328 1295
rect 35260 1215 35328 1239
rect 35260 1159 35266 1215
rect 35322 1159 35328 1215
rect 35260 1147 35328 1159
rect 35452 3135 35520 3522
rect 35452 3079 35458 3135
rect 35514 3079 35520 3135
rect 35452 3055 35520 3079
rect 35452 2999 35458 3055
rect 35514 2999 35520 3055
rect 35452 2975 35520 2999
rect 35452 2919 35458 2975
rect 35514 2919 35520 2975
rect 35452 2895 35520 2919
rect 35452 2839 35458 2895
rect 35514 2839 35520 2895
rect 35452 2815 35520 2839
rect 35452 2759 35458 2815
rect 35514 2759 35520 2815
rect 35452 2735 35520 2759
rect 35452 2679 35458 2735
rect 35514 2679 35520 2735
rect 35452 2655 35520 2679
rect 35452 2599 35458 2655
rect 35514 2599 35520 2655
rect 35452 2575 35520 2599
rect 35452 2519 35458 2575
rect 35514 2519 35520 2575
rect 35452 2495 35520 2519
rect 35452 2439 35458 2495
rect 35514 2439 35520 2495
rect 35452 2415 35520 2439
rect 35452 2359 35458 2415
rect 35514 2359 35520 2415
rect 35452 2335 35520 2359
rect 35452 2279 35458 2335
rect 35514 2279 35520 2335
rect 35452 2255 35520 2279
rect 35452 2199 35458 2255
rect 35514 2199 35520 2255
rect 35452 2175 35520 2199
rect 35452 2119 35458 2175
rect 35514 2119 35520 2175
rect 35452 2095 35520 2119
rect 35452 2039 35458 2095
rect 35514 2039 35520 2095
rect 35452 2015 35520 2039
rect 35452 1959 35458 2015
rect 35514 1959 35520 2015
rect 35452 1935 35520 1959
rect 35452 1879 35458 1935
rect 35514 1879 35520 1935
rect 35452 1855 35520 1879
rect 35452 1799 35458 1855
rect 35514 1799 35520 1855
rect 35452 1775 35520 1799
rect 35452 1719 35458 1775
rect 35514 1719 35520 1775
rect 35452 1695 35520 1719
rect 35452 1639 35458 1695
rect 35514 1639 35520 1695
rect 35452 1615 35520 1639
rect 35452 1559 35458 1615
rect 35514 1559 35520 1615
rect 35452 1535 35520 1559
rect 35452 1479 35458 1535
rect 35514 1479 35520 1535
rect 35452 1455 35520 1479
rect 35452 1399 35458 1455
rect 35514 1399 35520 1455
rect 35452 1375 35520 1399
rect 35452 1319 35458 1375
rect 35514 1319 35520 1375
rect 35452 1295 35520 1319
rect 35452 1239 35458 1295
rect 35514 1239 35520 1295
rect 35452 1215 35520 1239
rect 35452 1159 35458 1215
rect 35514 1159 35520 1215
rect 35452 1147 35520 1159
rect 35644 3135 35712 3522
rect 35644 3079 35650 3135
rect 35706 3079 35712 3135
rect 35644 3055 35712 3079
rect 35644 2999 35650 3055
rect 35706 2999 35712 3055
rect 35644 2975 35712 2999
rect 35644 2919 35650 2975
rect 35706 2919 35712 2975
rect 35644 2895 35712 2919
rect 35644 2839 35650 2895
rect 35706 2839 35712 2895
rect 35644 2815 35712 2839
rect 35644 2759 35650 2815
rect 35706 2759 35712 2815
rect 35644 2735 35712 2759
rect 35644 2679 35650 2735
rect 35706 2679 35712 2735
rect 35644 2655 35712 2679
rect 35644 2599 35650 2655
rect 35706 2599 35712 2655
rect 35644 2575 35712 2599
rect 35644 2519 35650 2575
rect 35706 2519 35712 2575
rect 35644 2495 35712 2519
rect 35644 2439 35650 2495
rect 35706 2439 35712 2495
rect 35644 2415 35712 2439
rect 35644 2359 35650 2415
rect 35706 2359 35712 2415
rect 35644 2335 35712 2359
rect 35644 2279 35650 2335
rect 35706 2279 35712 2335
rect 35644 2255 35712 2279
rect 35644 2199 35650 2255
rect 35706 2199 35712 2255
rect 35644 2175 35712 2199
rect 35644 2119 35650 2175
rect 35706 2119 35712 2175
rect 35644 2095 35712 2119
rect 35644 2039 35650 2095
rect 35706 2039 35712 2095
rect 35644 2015 35712 2039
rect 35644 1959 35650 2015
rect 35706 1959 35712 2015
rect 35644 1935 35712 1959
rect 35644 1879 35650 1935
rect 35706 1879 35712 1935
rect 35644 1855 35712 1879
rect 35644 1799 35650 1855
rect 35706 1799 35712 1855
rect 35644 1775 35712 1799
rect 35644 1719 35650 1775
rect 35706 1719 35712 1775
rect 35644 1695 35712 1719
rect 35644 1639 35650 1695
rect 35706 1639 35712 1695
rect 35644 1615 35712 1639
rect 35644 1559 35650 1615
rect 35706 1559 35712 1615
rect 35644 1535 35712 1559
rect 35644 1479 35650 1535
rect 35706 1479 35712 1535
rect 35644 1455 35712 1479
rect 35644 1399 35650 1455
rect 35706 1399 35712 1455
rect 35644 1375 35712 1399
rect 35644 1319 35650 1375
rect 35706 1319 35712 1375
rect 35644 1295 35712 1319
rect 35644 1239 35650 1295
rect 35706 1239 35712 1295
rect 35644 1215 35712 1239
rect 35644 1159 35650 1215
rect 35706 1159 35712 1215
rect 35644 1147 35712 1159
rect 35836 3135 35904 3522
rect 35836 3079 35842 3135
rect 35898 3079 35904 3135
rect 35836 3055 35904 3079
rect 35836 2999 35842 3055
rect 35898 2999 35904 3055
rect 35836 2975 35904 2999
rect 35836 2919 35842 2975
rect 35898 2919 35904 2975
rect 35836 2895 35904 2919
rect 35836 2839 35842 2895
rect 35898 2839 35904 2895
rect 35836 2815 35904 2839
rect 35836 2759 35842 2815
rect 35898 2759 35904 2815
rect 35836 2735 35904 2759
rect 35836 2679 35842 2735
rect 35898 2679 35904 2735
rect 35836 2655 35904 2679
rect 35836 2599 35842 2655
rect 35898 2599 35904 2655
rect 35836 2575 35904 2599
rect 35836 2519 35842 2575
rect 35898 2519 35904 2575
rect 35836 2495 35904 2519
rect 35836 2439 35842 2495
rect 35898 2439 35904 2495
rect 35836 2415 35904 2439
rect 35836 2359 35842 2415
rect 35898 2359 35904 2415
rect 35836 2335 35904 2359
rect 35836 2279 35842 2335
rect 35898 2279 35904 2335
rect 35836 2255 35904 2279
rect 35836 2199 35842 2255
rect 35898 2199 35904 2255
rect 35836 2175 35904 2199
rect 35836 2119 35842 2175
rect 35898 2119 35904 2175
rect 35836 2095 35904 2119
rect 35836 2039 35842 2095
rect 35898 2039 35904 2095
rect 35836 2015 35904 2039
rect 35836 1959 35842 2015
rect 35898 1959 35904 2015
rect 35836 1935 35904 1959
rect 35836 1879 35842 1935
rect 35898 1879 35904 1935
rect 35836 1855 35904 1879
rect 35836 1799 35842 1855
rect 35898 1799 35904 1855
rect 35836 1775 35904 1799
rect 35836 1719 35842 1775
rect 35898 1719 35904 1775
rect 35836 1695 35904 1719
rect 35836 1639 35842 1695
rect 35898 1639 35904 1695
rect 35836 1615 35904 1639
rect 35836 1559 35842 1615
rect 35898 1559 35904 1615
rect 35836 1535 35904 1559
rect 35836 1479 35842 1535
rect 35898 1479 35904 1535
rect 35836 1455 35904 1479
rect 35836 1399 35842 1455
rect 35898 1399 35904 1455
rect 35836 1375 35904 1399
rect 35836 1319 35842 1375
rect 35898 1319 35904 1375
rect 35836 1295 35904 1319
rect 35836 1239 35842 1295
rect 35898 1239 35904 1295
rect 35836 1215 35904 1239
rect 35836 1159 35842 1215
rect 35898 1159 35904 1215
rect 35836 1147 35904 1159
rect 36028 3135 36096 3522
rect 36028 3079 36034 3135
rect 36090 3079 36096 3135
rect 36028 3055 36096 3079
rect 36028 2999 36034 3055
rect 36090 2999 36096 3055
rect 36028 2975 36096 2999
rect 36028 2919 36034 2975
rect 36090 2919 36096 2975
rect 36028 2895 36096 2919
rect 36028 2839 36034 2895
rect 36090 2839 36096 2895
rect 36028 2815 36096 2839
rect 36028 2759 36034 2815
rect 36090 2759 36096 2815
rect 36028 2735 36096 2759
rect 36028 2679 36034 2735
rect 36090 2679 36096 2735
rect 36028 2655 36096 2679
rect 36028 2599 36034 2655
rect 36090 2599 36096 2655
rect 36028 2575 36096 2599
rect 36028 2519 36034 2575
rect 36090 2519 36096 2575
rect 36028 2495 36096 2519
rect 36028 2439 36034 2495
rect 36090 2439 36096 2495
rect 36028 2415 36096 2439
rect 36028 2359 36034 2415
rect 36090 2359 36096 2415
rect 36028 2335 36096 2359
rect 36028 2279 36034 2335
rect 36090 2279 36096 2335
rect 36028 2255 36096 2279
rect 36028 2199 36034 2255
rect 36090 2199 36096 2255
rect 36028 2175 36096 2199
rect 36028 2119 36034 2175
rect 36090 2119 36096 2175
rect 36028 2095 36096 2119
rect 36028 2039 36034 2095
rect 36090 2039 36096 2095
rect 36028 2015 36096 2039
rect 36028 1959 36034 2015
rect 36090 1959 36096 2015
rect 36028 1935 36096 1959
rect 36028 1879 36034 1935
rect 36090 1879 36096 1935
rect 36028 1855 36096 1879
rect 36028 1799 36034 1855
rect 36090 1799 36096 1855
rect 36028 1775 36096 1799
rect 36028 1719 36034 1775
rect 36090 1719 36096 1775
rect 36028 1695 36096 1719
rect 36028 1639 36034 1695
rect 36090 1639 36096 1695
rect 36028 1615 36096 1639
rect 36028 1559 36034 1615
rect 36090 1559 36096 1615
rect 36028 1535 36096 1559
rect 36028 1479 36034 1535
rect 36090 1479 36096 1535
rect 36028 1455 36096 1479
rect 36028 1399 36034 1455
rect 36090 1399 36096 1455
rect 36028 1375 36096 1399
rect 36028 1319 36034 1375
rect 36090 1319 36096 1375
rect 36028 1295 36096 1319
rect 36028 1239 36034 1295
rect 36090 1239 36096 1295
rect 36028 1215 36096 1239
rect 36028 1159 36034 1215
rect 36090 1159 36096 1215
rect 36028 1147 36096 1159
rect 36220 3135 36288 3522
rect 36220 3079 36226 3135
rect 36282 3079 36288 3135
rect 36220 3055 36288 3079
rect 36220 2999 36226 3055
rect 36282 2999 36288 3055
rect 36220 2975 36288 2999
rect 36220 2919 36226 2975
rect 36282 2919 36288 2975
rect 36220 2895 36288 2919
rect 36220 2839 36226 2895
rect 36282 2839 36288 2895
rect 36220 2815 36288 2839
rect 36220 2759 36226 2815
rect 36282 2759 36288 2815
rect 36220 2735 36288 2759
rect 36220 2679 36226 2735
rect 36282 2679 36288 2735
rect 36220 2655 36288 2679
rect 36220 2599 36226 2655
rect 36282 2599 36288 2655
rect 36220 2575 36288 2599
rect 36220 2519 36226 2575
rect 36282 2519 36288 2575
rect 36220 2495 36288 2519
rect 36220 2439 36226 2495
rect 36282 2439 36288 2495
rect 36220 2415 36288 2439
rect 36220 2359 36226 2415
rect 36282 2359 36288 2415
rect 36220 2335 36288 2359
rect 36220 2279 36226 2335
rect 36282 2279 36288 2335
rect 36220 2255 36288 2279
rect 36220 2199 36226 2255
rect 36282 2199 36288 2255
rect 36220 2175 36288 2199
rect 36220 2119 36226 2175
rect 36282 2119 36288 2175
rect 36220 2095 36288 2119
rect 36220 2039 36226 2095
rect 36282 2039 36288 2095
rect 36220 2015 36288 2039
rect 36220 1959 36226 2015
rect 36282 1959 36288 2015
rect 36220 1935 36288 1959
rect 36220 1879 36226 1935
rect 36282 1879 36288 1935
rect 36220 1855 36288 1879
rect 36220 1799 36226 1855
rect 36282 1799 36288 1855
rect 36220 1775 36288 1799
rect 36220 1719 36226 1775
rect 36282 1719 36288 1775
rect 36220 1695 36288 1719
rect 36220 1639 36226 1695
rect 36282 1639 36288 1695
rect 36220 1615 36288 1639
rect 36220 1559 36226 1615
rect 36282 1559 36288 1615
rect 36220 1535 36288 1559
rect 36220 1479 36226 1535
rect 36282 1479 36288 1535
rect 36220 1455 36288 1479
rect 36220 1399 36226 1455
rect 36282 1399 36288 1455
rect 36220 1375 36288 1399
rect 36220 1319 36226 1375
rect 36282 1319 36288 1375
rect 36220 1295 36288 1319
rect 36220 1239 36226 1295
rect 36282 1239 36288 1295
rect 36220 1215 36288 1239
rect 36220 1159 36226 1215
rect 36282 1159 36288 1215
rect 36220 1147 36288 1159
rect 36412 3135 36480 3522
rect 36412 3079 36418 3135
rect 36474 3079 36480 3135
rect 36412 3055 36480 3079
rect 36412 2999 36418 3055
rect 36474 2999 36480 3055
rect 36412 2975 36480 2999
rect 36412 2919 36418 2975
rect 36474 2919 36480 2975
rect 36412 2895 36480 2919
rect 36412 2839 36418 2895
rect 36474 2839 36480 2895
rect 36412 2815 36480 2839
rect 36412 2759 36418 2815
rect 36474 2759 36480 2815
rect 36412 2735 36480 2759
rect 36412 2679 36418 2735
rect 36474 2679 36480 2735
rect 36412 2655 36480 2679
rect 36412 2599 36418 2655
rect 36474 2599 36480 2655
rect 36412 2575 36480 2599
rect 36412 2519 36418 2575
rect 36474 2519 36480 2575
rect 36412 2495 36480 2519
rect 36412 2439 36418 2495
rect 36474 2439 36480 2495
rect 36412 2415 36480 2439
rect 36412 2359 36418 2415
rect 36474 2359 36480 2415
rect 36412 2335 36480 2359
rect 36412 2279 36418 2335
rect 36474 2279 36480 2335
rect 36412 2255 36480 2279
rect 36412 2199 36418 2255
rect 36474 2199 36480 2255
rect 36412 2175 36480 2199
rect 36412 2119 36418 2175
rect 36474 2119 36480 2175
rect 36412 2095 36480 2119
rect 36412 2039 36418 2095
rect 36474 2039 36480 2095
rect 36412 2015 36480 2039
rect 36412 1959 36418 2015
rect 36474 1959 36480 2015
rect 36412 1935 36480 1959
rect 36412 1879 36418 1935
rect 36474 1879 36480 1935
rect 36412 1855 36480 1879
rect 36412 1799 36418 1855
rect 36474 1799 36480 1855
rect 36412 1775 36480 1799
rect 36412 1719 36418 1775
rect 36474 1719 36480 1775
rect 36412 1695 36480 1719
rect 36412 1639 36418 1695
rect 36474 1639 36480 1695
rect 36412 1615 36480 1639
rect 36412 1559 36418 1615
rect 36474 1559 36480 1615
rect 36412 1535 36480 1559
rect 36412 1479 36418 1535
rect 36474 1479 36480 1535
rect 36412 1455 36480 1479
rect 36412 1399 36418 1455
rect 36474 1399 36480 1455
rect 36412 1375 36480 1399
rect 36412 1319 36418 1375
rect 36474 1319 36480 1375
rect 36412 1295 36480 1319
rect 36412 1239 36418 1295
rect 36474 1239 36480 1295
rect 36412 1215 36480 1239
rect 36412 1159 36418 1215
rect 36474 1159 36480 1215
rect 36412 1147 36480 1159
rect 36604 3135 36672 3522
rect 36604 3079 36610 3135
rect 36666 3079 36672 3135
rect 36604 3055 36672 3079
rect 36604 2999 36610 3055
rect 36666 2999 36672 3055
rect 36604 2975 36672 2999
rect 36604 2919 36610 2975
rect 36666 2919 36672 2975
rect 36604 2895 36672 2919
rect 36604 2839 36610 2895
rect 36666 2839 36672 2895
rect 36604 2815 36672 2839
rect 36604 2759 36610 2815
rect 36666 2759 36672 2815
rect 36604 2735 36672 2759
rect 36604 2679 36610 2735
rect 36666 2679 36672 2735
rect 36604 2655 36672 2679
rect 36604 2599 36610 2655
rect 36666 2599 36672 2655
rect 36604 2575 36672 2599
rect 36604 2519 36610 2575
rect 36666 2519 36672 2575
rect 36604 2495 36672 2519
rect 36604 2439 36610 2495
rect 36666 2439 36672 2495
rect 36604 2415 36672 2439
rect 36604 2359 36610 2415
rect 36666 2359 36672 2415
rect 36604 2335 36672 2359
rect 36604 2279 36610 2335
rect 36666 2279 36672 2335
rect 36604 2255 36672 2279
rect 36604 2199 36610 2255
rect 36666 2199 36672 2255
rect 36604 2175 36672 2199
rect 36604 2119 36610 2175
rect 36666 2119 36672 2175
rect 36604 2095 36672 2119
rect 36604 2039 36610 2095
rect 36666 2039 36672 2095
rect 36604 2015 36672 2039
rect 36604 1959 36610 2015
rect 36666 1959 36672 2015
rect 36604 1935 36672 1959
rect 36604 1879 36610 1935
rect 36666 1879 36672 1935
rect 36604 1855 36672 1879
rect 36604 1799 36610 1855
rect 36666 1799 36672 1855
rect 36604 1775 36672 1799
rect 36604 1719 36610 1775
rect 36666 1719 36672 1775
rect 36604 1695 36672 1719
rect 36604 1639 36610 1695
rect 36666 1639 36672 1695
rect 36604 1615 36672 1639
rect 36604 1559 36610 1615
rect 36666 1559 36672 1615
rect 36604 1535 36672 1559
rect 36604 1479 36610 1535
rect 36666 1479 36672 1535
rect 36604 1455 36672 1479
rect 36604 1399 36610 1455
rect 36666 1399 36672 1455
rect 36604 1375 36672 1399
rect 36604 1319 36610 1375
rect 36666 1319 36672 1375
rect 36604 1295 36672 1319
rect 36604 1239 36610 1295
rect 36666 1239 36672 1295
rect 36604 1215 36672 1239
rect 36604 1159 36610 1215
rect 36666 1159 36672 1215
rect 36604 1147 36672 1159
rect 36796 3135 36864 3522
rect 36796 3079 36802 3135
rect 36858 3079 36864 3135
rect 36796 3055 36864 3079
rect 36796 2999 36802 3055
rect 36858 2999 36864 3055
rect 36796 2975 36864 2999
rect 36796 2919 36802 2975
rect 36858 2919 36864 2975
rect 36796 2895 36864 2919
rect 36796 2839 36802 2895
rect 36858 2839 36864 2895
rect 36796 2815 36864 2839
rect 36796 2759 36802 2815
rect 36858 2759 36864 2815
rect 36796 2735 36864 2759
rect 36796 2679 36802 2735
rect 36858 2679 36864 2735
rect 36796 2655 36864 2679
rect 36796 2599 36802 2655
rect 36858 2599 36864 2655
rect 36796 2575 36864 2599
rect 36796 2519 36802 2575
rect 36858 2519 36864 2575
rect 36796 2495 36864 2519
rect 36796 2439 36802 2495
rect 36858 2439 36864 2495
rect 36796 2415 36864 2439
rect 36796 2359 36802 2415
rect 36858 2359 36864 2415
rect 36796 2335 36864 2359
rect 36796 2279 36802 2335
rect 36858 2279 36864 2335
rect 36796 2255 36864 2279
rect 36796 2199 36802 2255
rect 36858 2199 36864 2255
rect 36796 2175 36864 2199
rect 36796 2119 36802 2175
rect 36858 2119 36864 2175
rect 36796 2095 36864 2119
rect 36796 2039 36802 2095
rect 36858 2039 36864 2095
rect 36796 2015 36864 2039
rect 36796 1959 36802 2015
rect 36858 1959 36864 2015
rect 36796 1935 36864 1959
rect 36796 1879 36802 1935
rect 36858 1879 36864 1935
rect 36796 1855 36864 1879
rect 36796 1799 36802 1855
rect 36858 1799 36864 1855
rect 36796 1775 36864 1799
rect 36796 1719 36802 1775
rect 36858 1719 36864 1775
rect 36796 1695 36864 1719
rect 36796 1639 36802 1695
rect 36858 1639 36864 1695
rect 36796 1615 36864 1639
rect 36796 1559 36802 1615
rect 36858 1559 36864 1615
rect 36796 1535 36864 1559
rect 36796 1479 36802 1535
rect 36858 1479 36864 1535
rect 36796 1455 36864 1479
rect 36796 1399 36802 1455
rect 36858 1399 36864 1455
rect 36796 1375 36864 1399
rect 36796 1319 36802 1375
rect 36858 1319 36864 1375
rect 36796 1295 36864 1319
rect 36796 1239 36802 1295
rect 36858 1239 36864 1295
rect 36796 1215 36864 1239
rect 36796 1159 36802 1215
rect 36858 1159 36864 1215
rect 36796 1147 36864 1159
rect 36988 3135 37056 3522
rect 36988 3079 36994 3135
rect 37050 3079 37056 3135
rect 36988 3055 37056 3079
rect 36988 2999 36994 3055
rect 37050 2999 37056 3055
rect 36988 2975 37056 2999
rect 36988 2919 36994 2975
rect 37050 2919 37056 2975
rect 36988 2895 37056 2919
rect 36988 2839 36994 2895
rect 37050 2839 37056 2895
rect 36988 2815 37056 2839
rect 36988 2759 36994 2815
rect 37050 2759 37056 2815
rect 36988 2735 37056 2759
rect 36988 2679 36994 2735
rect 37050 2679 37056 2735
rect 36988 2655 37056 2679
rect 36988 2599 36994 2655
rect 37050 2599 37056 2655
rect 36988 2575 37056 2599
rect 36988 2519 36994 2575
rect 37050 2519 37056 2575
rect 36988 2495 37056 2519
rect 36988 2439 36994 2495
rect 37050 2439 37056 2495
rect 36988 2415 37056 2439
rect 36988 2359 36994 2415
rect 37050 2359 37056 2415
rect 36988 2335 37056 2359
rect 36988 2279 36994 2335
rect 37050 2279 37056 2335
rect 36988 2255 37056 2279
rect 36988 2199 36994 2255
rect 37050 2199 37056 2255
rect 36988 2175 37056 2199
rect 36988 2119 36994 2175
rect 37050 2119 37056 2175
rect 36988 2095 37056 2119
rect 36988 2039 36994 2095
rect 37050 2039 37056 2095
rect 36988 2015 37056 2039
rect 36988 1959 36994 2015
rect 37050 1959 37056 2015
rect 36988 1935 37056 1959
rect 36988 1879 36994 1935
rect 37050 1879 37056 1935
rect 36988 1855 37056 1879
rect 36988 1799 36994 1855
rect 37050 1799 37056 1855
rect 36988 1775 37056 1799
rect 36988 1719 36994 1775
rect 37050 1719 37056 1775
rect 36988 1695 37056 1719
rect 36988 1639 36994 1695
rect 37050 1639 37056 1695
rect 36988 1615 37056 1639
rect 36988 1559 36994 1615
rect 37050 1559 37056 1615
rect 36988 1535 37056 1559
rect 36988 1479 36994 1535
rect 37050 1479 37056 1535
rect 36988 1455 37056 1479
rect 36988 1399 36994 1455
rect 37050 1399 37056 1455
rect 36988 1375 37056 1399
rect 36988 1319 36994 1375
rect 37050 1319 37056 1375
rect 36988 1295 37056 1319
rect 36988 1239 36994 1295
rect 37050 1239 37056 1295
rect 36988 1215 37056 1239
rect 36988 1159 36994 1215
rect 37050 1159 37056 1215
rect 36988 1147 37056 1159
rect 37180 3135 37248 3522
rect 37180 3079 37186 3135
rect 37242 3079 37248 3135
rect 37180 3055 37248 3079
rect 37180 2999 37186 3055
rect 37242 2999 37248 3055
rect 37180 2975 37248 2999
rect 37180 2919 37186 2975
rect 37242 2919 37248 2975
rect 37180 2895 37248 2919
rect 37180 2839 37186 2895
rect 37242 2839 37248 2895
rect 37180 2815 37248 2839
rect 37180 2759 37186 2815
rect 37242 2759 37248 2815
rect 37180 2735 37248 2759
rect 37180 2679 37186 2735
rect 37242 2679 37248 2735
rect 37180 2655 37248 2679
rect 37180 2599 37186 2655
rect 37242 2599 37248 2655
rect 37180 2575 37248 2599
rect 37180 2519 37186 2575
rect 37242 2519 37248 2575
rect 37180 2495 37248 2519
rect 37180 2439 37186 2495
rect 37242 2439 37248 2495
rect 37180 2415 37248 2439
rect 37180 2359 37186 2415
rect 37242 2359 37248 2415
rect 37180 2335 37248 2359
rect 37180 2279 37186 2335
rect 37242 2279 37248 2335
rect 37180 2255 37248 2279
rect 37180 2199 37186 2255
rect 37242 2199 37248 2255
rect 37180 2175 37248 2199
rect 37180 2119 37186 2175
rect 37242 2119 37248 2175
rect 37180 2095 37248 2119
rect 37180 2039 37186 2095
rect 37242 2039 37248 2095
rect 37180 2015 37248 2039
rect 37180 1959 37186 2015
rect 37242 1959 37248 2015
rect 37180 1935 37248 1959
rect 37180 1879 37186 1935
rect 37242 1879 37248 1935
rect 37180 1855 37248 1879
rect 37180 1799 37186 1855
rect 37242 1799 37248 1855
rect 37180 1775 37248 1799
rect 37180 1719 37186 1775
rect 37242 1719 37248 1775
rect 37180 1695 37248 1719
rect 37180 1639 37186 1695
rect 37242 1639 37248 1695
rect 37180 1615 37248 1639
rect 37180 1559 37186 1615
rect 37242 1559 37248 1615
rect 37180 1535 37248 1559
rect 37180 1479 37186 1535
rect 37242 1479 37248 1535
rect 37180 1455 37248 1479
rect 37180 1399 37186 1455
rect 37242 1399 37248 1455
rect 37180 1375 37248 1399
rect 37180 1319 37186 1375
rect 37242 1319 37248 1375
rect 37180 1295 37248 1319
rect 37180 1239 37186 1295
rect 37242 1239 37248 1295
rect 37180 1215 37248 1239
rect 37180 1159 37186 1215
rect 37242 1159 37248 1215
rect 37180 1147 37248 1159
rect 37372 3135 37440 3522
rect 37372 3079 37378 3135
rect 37434 3079 37440 3135
rect 37372 3055 37440 3079
rect 37372 2999 37378 3055
rect 37434 2999 37440 3055
rect 37372 2975 37440 2999
rect 37372 2919 37378 2975
rect 37434 2919 37440 2975
rect 37372 2895 37440 2919
rect 37372 2839 37378 2895
rect 37434 2839 37440 2895
rect 37372 2815 37440 2839
rect 37372 2759 37378 2815
rect 37434 2759 37440 2815
rect 37372 2735 37440 2759
rect 37372 2679 37378 2735
rect 37434 2679 37440 2735
rect 37372 2655 37440 2679
rect 37372 2599 37378 2655
rect 37434 2599 37440 2655
rect 37372 2575 37440 2599
rect 37372 2519 37378 2575
rect 37434 2519 37440 2575
rect 37372 2495 37440 2519
rect 37372 2439 37378 2495
rect 37434 2439 37440 2495
rect 37372 2415 37440 2439
rect 37372 2359 37378 2415
rect 37434 2359 37440 2415
rect 37372 2335 37440 2359
rect 37372 2279 37378 2335
rect 37434 2279 37440 2335
rect 37372 2255 37440 2279
rect 37372 2199 37378 2255
rect 37434 2199 37440 2255
rect 37372 2175 37440 2199
rect 37372 2119 37378 2175
rect 37434 2119 37440 2175
rect 37372 2095 37440 2119
rect 37372 2039 37378 2095
rect 37434 2039 37440 2095
rect 37372 2015 37440 2039
rect 37372 1959 37378 2015
rect 37434 1959 37440 2015
rect 37372 1935 37440 1959
rect 37372 1879 37378 1935
rect 37434 1879 37440 1935
rect 37372 1855 37440 1879
rect 37372 1799 37378 1855
rect 37434 1799 37440 1855
rect 37372 1775 37440 1799
rect 37372 1719 37378 1775
rect 37434 1719 37440 1775
rect 37372 1695 37440 1719
rect 37372 1639 37378 1695
rect 37434 1639 37440 1695
rect 37372 1615 37440 1639
rect 37372 1559 37378 1615
rect 37434 1559 37440 1615
rect 37372 1535 37440 1559
rect 37372 1479 37378 1535
rect 37434 1479 37440 1535
rect 37372 1455 37440 1479
rect 37372 1399 37378 1455
rect 37434 1399 37440 1455
rect 37372 1375 37440 1399
rect 37372 1319 37378 1375
rect 37434 1319 37440 1375
rect 37372 1295 37440 1319
rect 37372 1239 37378 1295
rect 37434 1239 37440 1295
rect 37372 1215 37440 1239
rect 37372 1159 37378 1215
rect 37434 1159 37440 1215
rect 37372 1147 37440 1159
rect 37564 3135 37632 3522
rect 37564 3079 37570 3135
rect 37626 3079 37632 3135
rect 37564 3055 37632 3079
rect 37564 2999 37570 3055
rect 37626 2999 37632 3055
rect 37564 2975 37632 2999
rect 37564 2919 37570 2975
rect 37626 2919 37632 2975
rect 37564 2895 37632 2919
rect 37564 2839 37570 2895
rect 37626 2839 37632 2895
rect 37564 2815 37632 2839
rect 37564 2759 37570 2815
rect 37626 2759 37632 2815
rect 37564 2735 37632 2759
rect 37564 2679 37570 2735
rect 37626 2679 37632 2735
rect 37564 2655 37632 2679
rect 37564 2599 37570 2655
rect 37626 2599 37632 2655
rect 37564 2575 37632 2599
rect 37564 2519 37570 2575
rect 37626 2519 37632 2575
rect 37564 2495 37632 2519
rect 37564 2439 37570 2495
rect 37626 2439 37632 2495
rect 37564 2415 37632 2439
rect 37564 2359 37570 2415
rect 37626 2359 37632 2415
rect 37564 2335 37632 2359
rect 37564 2279 37570 2335
rect 37626 2279 37632 2335
rect 37564 2255 37632 2279
rect 37564 2199 37570 2255
rect 37626 2199 37632 2255
rect 37564 2175 37632 2199
rect 37564 2119 37570 2175
rect 37626 2119 37632 2175
rect 37564 2095 37632 2119
rect 37564 2039 37570 2095
rect 37626 2039 37632 2095
rect 37564 2015 37632 2039
rect 37564 1959 37570 2015
rect 37626 1959 37632 2015
rect 37564 1935 37632 1959
rect 37564 1879 37570 1935
rect 37626 1879 37632 1935
rect 37564 1855 37632 1879
rect 37564 1799 37570 1855
rect 37626 1799 37632 1855
rect 37564 1775 37632 1799
rect 37564 1719 37570 1775
rect 37626 1719 37632 1775
rect 37564 1695 37632 1719
rect 37564 1639 37570 1695
rect 37626 1639 37632 1695
rect 37564 1615 37632 1639
rect 37564 1559 37570 1615
rect 37626 1559 37632 1615
rect 37564 1535 37632 1559
rect 37564 1479 37570 1535
rect 37626 1479 37632 1535
rect 37564 1455 37632 1479
rect 37564 1399 37570 1455
rect 37626 1399 37632 1455
rect 37564 1375 37632 1399
rect 37564 1319 37570 1375
rect 37626 1319 37632 1375
rect 37564 1295 37632 1319
rect 37564 1239 37570 1295
rect 37626 1239 37632 1295
rect 37564 1215 37632 1239
rect 37564 1159 37570 1215
rect 37626 1159 37632 1215
rect 37564 1147 37632 1159
rect 37756 3135 37824 3522
rect 37756 3079 37762 3135
rect 37818 3079 37824 3135
rect 37756 3055 37824 3079
rect 37756 2999 37762 3055
rect 37818 2999 37824 3055
rect 37756 2975 37824 2999
rect 37756 2919 37762 2975
rect 37818 2919 37824 2975
rect 37756 2895 37824 2919
rect 37756 2839 37762 2895
rect 37818 2839 37824 2895
rect 37756 2815 37824 2839
rect 37756 2759 37762 2815
rect 37818 2759 37824 2815
rect 37756 2735 37824 2759
rect 37756 2679 37762 2735
rect 37818 2679 37824 2735
rect 37756 2655 37824 2679
rect 37756 2599 37762 2655
rect 37818 2599 37824 2655
rect 37756 2575 37824 2599
rect 37756 2519 37762 2575
rect 37818 2519 37824 2575
rect 37756 2495 37824 2519
rect 37756 2439 37762 2495
rect 37818 2439 37824 2495
rect 37756 2415 37824 2439
rect 37756 2359 37762 2415
rect 37818 2359 37824 2415
rect 37756 2335 37824 2359
rect 37756 2279 37762 2335
rect 37818 2279 37824 2335
rect 37756 2255 37824 2279
rect 37756 2199 37762 2255
rect 37818 2199 37824 2255
rect 37756 2175 37824 2199
rect 37756 2119 37762 2175
rect 37818 2119 37824 2175
rect 37756 2095 37824 2119
rect 37756 2039 37762 2095
rect 37818 2039 37824 2095
rect 37756 2015 37824 2039
rect 37756 1959 37762 2015
rect 37818 1959 37824 2015
rect 37756 1935 37824 1959
rect 37756 1879 37762 1935
rect 37818 1879 37824 1935
rect 37756 1855 37824 1879
rect 37756 1799 37762 1855
rect 37818 1799 37824 1855
rect 37756 1775 37824 1799
rect 37756 1719 37762 1775
rect 37818 1719 37824 1775
rect 37756 1695 37824 1719
rect 37756 1639 37762 1695
rect 37818 1639 37824 1695
rect 37756 1615 37824 1639
rect 37756 1559 37762 1615
rect 37818 1559 37824 1615
rect 37756 1535 37824 1559
rect 37756 1479 37762 1535
rect 37818 1479 37824 1535
rect 37756 1455 37824 1479
rect 37756 1399 37762 1455
rect 37818 1399 37824 1455
rect 37756 1375 37824 1399
rect 37756 1319 37762 1375
rect 37818 1319 37824 1375
rect 37756 1295 37824 1319
rect 37756 1239 37762 1295
rect 37818 1239 37824 1295
rect 37756 1215 37824 1239
rect 37756 1159 37762 1215
rect 37818 1159 37824 1215
rect 37756 1147 37824 1159
rect 37948 3135 38016 3522
rect 37948 3079 37954 3135
rect 38010 3079 38016 3135
rect 37948 3055 38016 3079
rect 37948 2999 37954 3055
rect 38010 2999 38016 3055
rect 37948 2975 38016 2999
rect 37948 2919 37954 2975
rect 38010 2919 38016 2975
rect 37948 2895 38016 2919
rect 37948 2839 37954 2895
rect 38010 2839 38016 2895
rect 37948 2815 38016 2839
rect 37948 2759 37954 2815
rect 38010 2759 38016 2815
rect 37948 2735 38016 2759
rect 37948 2679 37954 2735
rect 38010 2679 38016 2735
rect 37948 2655 38016 2679
rect 37948 2599 37954 2655
rect 38010 2599 38016 2655
rect 37948 2575 38016 2599
rect 37948 2519 37954 2575
rect 38010 2519 38016 2575
rect 37948 2495 38016 2519
rect 37948 2439 37954 2495
rect 38010 2439 38016 2495
rect 37948 2415 38016 2439
rect 37948 2359 37954 2415
rect 38010 2359 38016 2415
rect 37948 2335 38016 2359
rect 37948 2279 37954 2335
rect 38010 2279 38016 2335
rect 37948 2255 38016 2279
rect 37948 2199 37954 2255
rect 38010 2199 38016 2255
rect 37948 2175 38016 2199
rect 37948 2119 37954 2175
rect 38010 2119 38016 2175
rect 37948 2095 38016 2119
rect 37948 2039 37954 2095
rect 38010 2039 38016 2095
rect 37948 2015 38016 2039
rect 37948 1959 37954 2015
rect 38010 1959 38016 2015
rect 37948 1935 38016 1959
rect 37948 1879 37954 1935
rect 38010 1879 38016 1935
rect 37948 1855 38016 1879
rect 37948 1799 37954 1855
rect 38010 1799 38016 1855
rect 37948 1775 38016 1799
rect 37948 1719 37954 1775
rect 38010 1719 38016 1775
rect 37948 1695 38016 1719
rect 37948 1639 37954 1695
rect 38010 1639 38016 1695
rect 37948 1615 38016 1639
rect 37948 1559 37954 1615
rect 38010 1559 38016 1615
rect 37948 1535 38016 1559
rect 37948 1479 37954 1535
rect 38010 1479 38016 1535
rect 37948 1455 38016 1479
rect 37948 1399 37954 1455
rect 38010 1399 38016 1455
rect 37948 1375 38016 1399
rect 37948 1319 37954 1375
rect 38010 1319 38016 1375
rect 37948 1295 38016 1319
rect 37948 1239 37954 1295
rect 38010 1239 38016 1295
rect 37948 1215 38016 1239
rect 37948 1159 37954 1215
rect 38010 1159 38016 1215
rect 37948 1147 38016 1159
rect 38140 3135 38208 3522
rect 38140 3079 38146 3135
rect 38202 3079 38208 3135
rect 38140 3055 38208 3079
rect 38140 2999 38146 3055
rect 38202 2999 38208 3055
rect 38140 2975 38208 2999
rect 38140 2919 38146 2975
rect 38202 2919 38208 2975
rect 38140 2895 38208 2919
rect 38140 2839 38146 2895
rect 38202 2839 38208 2895
rect 38140 2815 38208 2839
rect 38140 2759 38146 2815
rect 38202 2759 38208 2815
rect 38140 2735 38208 2759
rect 38140 2679 38146 2735
rect 38202 2679 38208 2735
rect 38140 2655 38208 2679
rect 38140 2599 38146 2655
rect 38202 2599 38208 2655
rect 38140 2575 38208 2599
rect 38140 2519 38146 2575
rect 38202 2519 38208 2575
rect 38140 2495 38208 2519
rect 38140 2439 38146 2495
rect 38202 2439 38208 2495
rect 38140 2415 38208 2439
rect 38140 2359 38146 2415
rect 38202 2359 38208 2415
rect 38140 2335 38208 2359
rect 38140 2279 38146 2335
rect 38202 2279 38208 2335
rect 38140 2255 38208 2279
rect 38140 2199 38146 2255
rect 38202 2199 38208 2255
rect 38140 2175 38208 2199
rect 38140 2119 38146 2175
rect 38202 2119 38208 2175
rect 38140 2095 38208 2119
rect 38140 2039 38146 2095
rect 38202 2039 38208 2095
rect 38140 2015 38208 2039
rect 38140 1959 38146 2015
rect 38202 1959 38208 2015
rect 38140 1935 38208 1959
rect 38140 1879 38146 1935
rect 38202 1879 38208 1935
rect 38140 1855 38208 1879
rect 38140 1799 38146 1855
rect 38202 1799 38208 1855
rect 38140 1775 38208 1799
rect 38140 1719 38146 1775
rect 38202 1719 38208 1775
rect 38140 1695 38208 1719
rect 38140 1639 38146 1695
rect 38202 1639 38208 1695
rect 38140 1615 38208 1639
rect 38140 1559 38146 1615
rect 38202 1559 38208 1615
rect 38140 1535 38208 1559
rect 38140 1479 38146 1535
rect 38202 1479 38208 1535
rect 38140 1455 38208 1479
rect 38140 1399 38146 1455
rect 38202 1399 38208 1455
rect 38140 1375 38208 1399
rect 38140 1319 38146 1375
rect 38202 1319 38208 1375
rect 38140 1295 38208 1319
rect 38140 1239 38146 1295
rect 38202 1239 38208 1295
rect 38140 1215 38208 1239
rect 38140 1159 38146 1215
rect 38202 1159 38208 1215
rect 38140 1147 38208 1159
rect 38332 3135 38400 3522
rect 38332 3079 38338 3135
rect 38394 3079 38400 3135
rect 38332 3055 38400 3079
rect 38332 2999 38338 3055
rect 38394 2999 38400 3055
rect 38332 2975 38400 2999
rect 38332 2919 38338 2975
rect 38394 2919 38400 2975
rect 38332 2895 38400 2919
rect 38332 2839 38338 2895
rect 38394 2839 38400 2895
rect 38332 2815 38400 2839
rect 38332 2759 38338 2815
rect 38394 2759 38400 2815
rect 38332 2735 38400 2759
rect 38332 2679 38338 2735
rect 38394 2679 38400 2735
rect 38332 2655 38400 2679
rect 38332 2599 38338 2655
rect 38394 2599 38400 2655
rect 38332 2575 38400 2599
rect 38332 2519 38338 2575
rect 38394 2519 38400 2575
rect 38332 2495 38400 2519
rect 38332 2439 38338 2495
rect 38394 2439 38400 2495
rect 38332 2415 38400 2439
rect 38332 2359 38338 2415
rect 38394 2359 38400 2415
rect 38332 2335 38400 2359
rect 38332 2279 38338 2335
rect 38394 2279 38400 2335
rect 38332 2255 38400 2279
rect 38332 2199 38338 2255
rect 38394 2199 38400 2255
rect 38332 2175 38400 2199
rect 38332 2119 38338 2175
rect 38394 2119 38400 2175
rect 38332 2095 38400 2119
rect 38332 2039 38338 2095
rect 38394 2039 38400 2095
rect 38332 2015 38400 2039
rect 38332 1959 38338 2015
rect 38394 1959 38400 2015
rect 38332 1935 38400 1959
rect 38332 1879 38338 1935
rect 38394 1879 38400 1935
rect 38332 1855 38400 1879
rect 38332 1799 38338 1855
rect 38394 1799 38400 1855
rect 38332 1775 38400 1799
rect 38332 1719 38338 1775
rect 38394 1719 38400 1775
rect 38332 1695 38400 1719
rect 38332 1639 38338 1695
rect 38394 1639 38400 1695
rect 38332 1615 38400 1639
rect 38332 1559 38338 1615
rect 38394 1559 38400 1615
rect 38332 1535 38400 1559
rect 38332 1479 38338 1535
rect 38394 1479 38400 1535
rect 38332 1455 38400 1479
rect 38332 1399 38338 1455
rect 38394 1399 38400 1455
rect 38332 1375 38400 1399
rect 38332 1319 38338 1375
rect 38394 1319 38400 1375
rect 38332 1295 38400 1319
rect 38332 1239 38338 1295
rect 38394 1239 38400 1295
rect 38332 1215 38400 1239
rect 38332 1159 38338 1215
rect 38394 1159 38400 1215
rect 38332 1147 38400 1159
rect 38524 3135 38592 3522
rect 38524 3079 38530 3135
rect 38586 3079 38592 3135
rect 38524 3055 38592 3079
rect 38524 2999 38530 3055
rect 38586 2999 38592 3055
rect 38524 2975 38592 2999
rect 38524 2919 38530 2975
rect 38586 2919 38592 2975
rect 38524 2895 38592 2919
rect 38524 2839 38530 2895
rect 38586 2839 38592 2895
rect 38524 2815 38592 2839
rect 38524 2759 38530 2815
rect 38586 2759 38592 2815
rect 38524 2735 38592 2759
rect 38524 2679 38530 2735
rect 38586 2679 38592 2735
rect 38524 2655 38592 2679
rect 38524 2599 38530 2655
rect 38586 2599 38592 2655
rect 38524 2575 38592 2599
rect 38524 2519 38530 2575
rect 38586 2519 38592 2575
rect 38524 2495 38592 2519
rect 38524 2439 38530 2495
rect 38586 2439 38592 2495
rect 38524 2415 38592 2439
rect 38524 2359 38530 2415
rect 38586 2359 38592 2415
rect 38524 2335 38592 2359
rect 38524 2279 38530 2335
rect 38586 2279 38592 2335
rect 38524 2255 38592 2279
rect 38524 2199 38530 2255
rect 38586 2199 38592 2255
rect 38524 2175 38592 2199
rect 38524 2119 38530 2175
rect 38586 2119 38592 2175
rect 38524 2095 38592 2119
rect 38524 2039 38530 2095
rect 38586 2039 38592 2095
rect 38524 2015 38592 2039
rect 38524 1959 38530 2015
rect 38586 1959 38592 2015
rect 38524 1935 38592 1959
rect 38524 1879 38530 1935
rect 38586 1879 38592 1935
rect 38524 1855 38592 1879
rect 38524 1799 38530 1855
rect 38586 1799 38592 1855
rect 38524 1775 38592 1799
rect 38524 1719 38530 1775
rect 38586 1719 38592 1775
rect 38524 1695 38592 1719
rect 38524 1639 38530 1695
rect 38586 1639 38592 1695
rect 38524 1615 38592 1639
rect 38524 1559 38530 1615
rect 38586 1559 38592 1615
rect 38524 1535 38592 1559
rect 38524 1479 38530 1535
rect 38586 1479 38592 1535
rect 38524 1455 38592 1479
rect 38524 1399 38530 1455
rect 38586 1399 38592 1455
rect 38524 1375 38592 1399
rect 38524 1319 38530 1375
rect 38586 1319 38592 1375
rect 38524 1295 38592 1319
rect 38524 1239 38530 1295
rect 38586 1239 38592 1295
rect 38524 1215 38592 1239
rect 38524 1159 38530 1215
rect 38586 1159 38592 1215
rect 38524 1147 38592 1159
use sky130_fd_pr__nfet_01v8_spf0jm  sky130_fd_pr__nfet_01v8_spf0jm_0
timestamp 1611881054
transform 1 0 33854 0 1 2147
box -4931 -1174 4931 1174
<< end >>
