magic
tech sky130A
magscale 1 2
timestamp 1607995095
<< pwell >>
rect -2457 -1530 2457 1530
<< nmos >>
rect -2261 -1320 -1861 1320
rect -1803 -1320 -1403 1320
rect -1345 -1320 -945 1320
rect -887 -1320 -487 1320
rect -429 -1320 -29 1320
rect 29 -1320 429 1320
rect 487 -1320 887 1320
rect 945 -1320 1345 1320
rect 1403 -1320 1803 1320
rect 1861 -1320 2261 1320
<< ndiff >>
rect -2319 1308 -2261 1320
rect -2319 -1308 -2307 1308
rect -2273 -1308 -2261 1308
rect -2319 -1320 -2261 -1308
rect -1861 1308 -1803 1320
rect -1861 -1308 -1849 1308
rect -1815 -1308 -1803 1308
rect -1861 -1320 -1803 -1308
rect -1403 1308 -1345 1320
rect -1403 -1308 -1391 1308
rect -1357 -1308 -1345 1308
rect -1403 -1320 -1345 -1308
rect -945 1308 -887 1320
rect -945 -1308 -933 1308
rect -899 -1308 -887 1308
rect -945 -1320 -887 -1308
rect -487 1308 -429 1320
rect -487 -1308 -475 1308
rect -441 -1308 -429 1308
rect -487 -1320 -429 -1308
rect -29 1308 29 1320
rect -29 -1308 -17 1308
rect 17 -1308 29 1308
rect -29 -1320 29 -1308
rect 429 1308 487 1320
rect 429 -1308 441 1308
rect 475 -1308 487 1308
rect 429 -1320 487 -1308
rect 887 1308 945 1320
rect 887 -1308 899 1308
rect 933 -1308 945 1308
rect 887 -1320 945 -1308
rect 1345 1308 1403 1320
rect 1345 -1308 1357 1308
rect 1391 -1308 1403 1308
rect 1345 -1320 1403 -1308
rect 1803 1308 1861 1320
rect 1803 -1308 1815 1308
rect 1849 -1308 1861 1308
rect 1803 -1320 1861 -1308
rect 2261 1308 2319 1320
rect 2261 -1308 2273 1308
rect 2307 -1308 2319 1308
rect 2261 -1320 2319 -1308
<< ndiffc >>
rect -2307 -1308 -2273 1308
rect -1849 -1308 -1815 1308
rect -1391 -1308 -1357 1308
rect -933 -1308 -899 1308
rect -475 -1308 -441 1308
rect -17 -1308 17 1308
rect 441 -1308 475 1308
rect 899 -1308 933 1308
rect 1357 -1308 1391 1308
rect 1815 -1308 1849 1308
rect 2273 -1308 2307 1308
<< psubdiff >>
rect -2421 1460 -2325 1494
rect 2325 1460 2421 1494
rect -2421 1398 -2387 1460
rect 2387 1398 2421 1460
rect -2421 -1460 -2387 -1398
rect 2387 -1460 2421 -1398
rect -2421 -1494 -2325 -1460
rect 2325 -1494 2421 -1460
<< psubdiffcont >>
rect -2325 1460 2325 1494
rect -2421 -1398 -2387 1398
rect 2387 -1398 2421 1398
rect -2325 -1494 2325 -1460
<< poly >>
rect -2114 1392 -2008 1408
rect -2114 1375 -2098 1392
rect -2261 1358 -2098 1375
rect -2024 1375 -2008 1392
rect -1656 1392 -1550 1408
rect -1656 1375 -1640 1392
rect -2024 1358 -1861 1375
rect -2261 1320 -1861 1358
rect -1803 1358 -1640 1375
rect -1566 1375 -1550 1392
rect -1198 1392 -1092 1408
rect -1198 1375 -1182 1392
rect -1566 1358 -1403 1375
rect -1803 1320 -1403 1358
rect -1345 1358 -1182 1375
rect -1108 1375 -1092 1392
rect -740 1392 -634 1408
rect -740 1375 -724 1392
rect -1108 1358 -945 1375
rect -1345 1320 -945 1358
rect -887 1358 -724 1375
rect -650 1375 -634 1392
rect -282 1392 -176 1408
rect -282 1375 -266 1392
rect -650 1358 -487 1375
rect -887 1320 -487 1358
rect -429 1358 -266 1375
rect -192 1375 -176 1392
rect 176 1392 282 1408
rect 176 1375 192 1392
rect -192 1358 -29 1375
rect -429 1320 -29 1358
rect 29 1358 192 1375
rect 266 1375 282 1392
rect 634 1392 740 1408
rect 634 1375 650 1392
rect 266 1358 429 1375
rect 29 1320 429 1358
rect 487 1358 650 1375
rect 724 1375 740 1392
rect 1092 1392 1198 1408
rect 1092 1375 1108 1392
rect 724 1358 887 1375
rect 487 1320 887 1358
rect 945 1358 1108 1375
rect 1182 1375 1198 1392
rect 1550 1392 1656 1408
rect 1550 1375 1566 1392
rect 1182 1358 1345 1375
rect 945 1320 1345 1358
rect 1403 1358 1566 1375
rect 1640 1375 1656 1392
rect 2008 1392 2114 1408
rect 2008 1375 2024 1392
rect 1640 1358 1803 1375
rect 1403 1320 1803 1358
rect 1861 1358 2024 1375
rect 2098 1375 2114 1392
rect 2098 1358 2261 1375
rect 1861 1320 2261 1358
rect -2261 -1358 -1861 -1320
rect -2261 -1375 -2098 -1358
rect -2114 -1392 -2098 -1375
rect -2024 -1375 -1861 -1358
rect -1803 -1358 -1403 -1320
rect -1803 -1375 -1640 -1358
rect -2024 -1392 -2008 -1375
rect -2114 -1408 -2008 -1392
rect -1656 -1392 -1640 -1375
rect -1566 -1375 -1403 -1358
rect -1345 -1358 -945 -1320
rect -1345 -1375 -1182 -1358
rect -1566 -1392 -1550 -1375
rect -1656 -1408 -1550 -1392
rect -1198 -1392 -1182 -1375
rect -1108 -1375 -945 -1358
rect -887 -1358 -487 -1320
rect -887 -1375 -724 -1358
rect -1108 -1392 -1092 -1375
rect -1198 -1408 -1092 -1392
rect -740 -1392 -724 -1375
rect -650 -1375 -487 -1358
rect -429 -1358 -29 -1320
rect -429 -1375 -266 -1358
rect -650 -1392 -634 -1375
rect -740 -1408 -634 -1392
rect -282 -1392 -266 -1375
rect -192 -1375 -29 -1358
rect 29 -1358 429 -1320
rect 29 -1375 192 -1358
rect -192 -1392 -176 -1375
rect -282 -1408 -176 -1392
rect 176 -1392 192 -1375
rect 266 -1375 429 -1358
rect 487 -1358 887 -1320
rect 487 -1375 650 -1358
rect 266 -1392 282 -1375
rect 176 -1408 282 -1392
rect 634 -1392 650 -1375
rect 724 -1375 887 -1358
rect 945 -1358 1345 -1320
rect 945 -1375 1108 -1358
rect 724 -1392 740 -1375
rect 634 -1408 740 -1392
rect 1092 -1392 1108 -1375
rect 1182 -1375 1345 -1358
rect 1403 -1358 1803 -1320
rect 1403 -1375 1566 -1358
rect 1182 -1392 1198 -1375
rect 1092 -1408 1198 -1392
rect 1550 -1392 1566 -1375
rect 1640 -1375 1803 -1358
rect 1861 -1358 2261 -1320
rect 1861 -1375 2024 -1358
rect 1640 -1392 1656 -1375
rect 1550 -1408 1656 -1392
rect 2008 -1392 2024 -1375
rect 2098 -1375 2261 -1358
rect 2098 -1392 2114 -1375
rect 2008 -1408 2114 -1392
<< polycont >>
rect -2098 1358 -2024 1392
rect -1640 1358 -1566 1392
rect -1182 1358 -1108 1392
rect -724 1358 -650 1392
rect -266 1358 -192 1392
rect 192 1358 266 1392
rect 650 1358 724 1392
rect 1108 1358 1182 1392
rect 1566 1358 1640 1392
rect 2024 1358 2098 1392
rect -2098 -1392 -2024 -1358
rect -1640 -1392 -1566 -1358
rect -1182 -1392 -1108 -1358
rect -724 -1392 -650 -1358
rect -266 -1392 -192 -1358
rect 192 -1392 266 -1358
rect 650 -1392 724 -1358
rect 1108 -1392 1182 -1358
rect 1566 -1392 1640 -1358
rect 2024 -1392 2098 -1358
<< locali >>
rect -2421 1460 -2325 1494
rect 2325 1460 2421 1494
rect -2421 1398 -2387 1460
rect 2387 1398 2421 1460
rect -2114 1358 -2098 1392
rect -2024 1358 -2008 1392
rect -1656 1358 -1640 1392
rect -1566 1358 -1550 1392
rect -1198 1358 -1182 1392
rect -1108 1358 -1092 1392
rect -740 1358 -724 1392
rect -650 1358 -634 1392
rect -282 1358 -266 1392
rect -192 1358 -176 1392
rect 176 1358 192 1392
rect 266 1358 282 1392
rect 634 1358 650 1392
rect 724 1358 740 1392
rect 1092 1358 1108 1392
rect 1182 1358 1198 1392
rect 1550 1358 1566 1392
rect 1640 1358 1656 1392
rect 2008 1358 2024 1392
rect 2098 1358 2114 1392
rect -2307 1308 -2273 1324
rect -2307 -1324 -2273 -1308
rect -1849 1308 -1815 1324
rect -1849 -1324 -1815 -1308
rect -1391 1308 -1357 1324
rect -1391 -1324 -1357 -1308
rect -933 1308 -899 1324
rect -933 -1324 -899 -1308
rect -475 1308 -441 1324
rect -475 -1324 -441 -1308
rect -17 1308 17 1324
rect -17 -1324 17 -1308
rect 441 1308 475 1324
rect 441 -1324 475 -1308
rect 899 1308 933 1324
rect 899 -1324 933 -1308
rect 1357 1308 1391 1324
rect 1357 -1324 1391 -1308
rect 1815 1308 1849 1324
rect 1815 -1324 1849 -1308
rect 2273 1308 2307 1324
rect 2273 -1324 2307 -1308
rect -2114 -1392 -2098 -1358
rect -2024 -1392 -2008 -1358
rect -1656 -1392 -1640 -1358
rect -1566 -1392 -1550 -1358
rect -1198 -1392 -1182 -1358
rect -1108 -1392 -1092 -1358
rect -740 -1392 -724 -1358
rect -650 -1392 -634 -1358
rect -282 -1392 -266 -1358
rect -192 -1392 -176 -1358
rect 176 -1392 192 -1358
rect 266 -1392 282 -1358
rect 634 -1392 650 -1358
rect 724 -1392 740 -1358
rect 1092 -1392 1108 -1358
rect 1182 -1392 1198 -1358
rect 1550 -1392 1566 -1358
rect 1640 -1392 1656 -1358
rect 2008 -1392 2024 -1358
rect 2098 -1392 2114 -1358
rect -2421 -1494 -2387 -1398
rect 2387 -1494 2421 -1398
<< viali >>
rect -2307 -1308 -2273 1308
rect -1849 -1308 -1815 1308
rect -1391 -1308 -1357 1308
rect -933 -1308 -899 1308
rect -475 -1308 -441 1308
rect -17 -1308 17 1308
rect 441 -1308 475 1308
rect 899 -1308 933 1308
rect 1357 -1308 1391 1308
rect 1815 -1308 1849 1308
rect 2273 -1308 2307 1308
rect -2387 -1494 -2325 -1460
rect -2325 -1494 2325 -1460
rect 2325 -1494 2387 -1460
<< metal1 >>
rect -2313 1308 -2267 1320
rect -2313 -1308 -2307 1308
rect -2273 -1308 -2267 1308
rect -2313 -1320 -2267 -1308
rect -1855 1308 -1809 1320
rect -1855 -1308 -1849 1308
rect -1815 -1308 -1809 1308
rect -1855 -1320 -1809 -1308
rect -1397 1308 -1351 1320
rect -1397 -1308 -1391 1308
rect -1357 -1308 -1351 1308
rect -1397 -1320 -1351 -1308
rect -939 1308 -893 1320
rect -939 -1308 -933 1308
rect -899 -1308 -893 1308
rect -939 -1320 -893 -1308
rect -481 1308 -435 1320
rect -481 -1308 -475 1308
rect -441 -1308 -435 1308
rect -481 -1320 -435 -1308
rect -23 1308 23 1320
rect -23 -1308 -17 1308
rect 17 -1308 23 1308
rect -23 -1320 23 -1308
rect 435 1308 481 1320
rect 435 -1308 441 1308
rect 475 -1308 481 1308
rect 435 -1320 481 -1308
rect 893 1308 939 1320
rect 893 -1308 899 1308
rect 933 -1308 939 1308
rect 893 -1320 939 -1308
rect 1351 1308 1397 1320
rect 1351 -1308 1357 1308
rect 1391 -1308 1397 1308
rect 1351 -1320 1397 -1308
rect 1809 1308 1855 1320
rect 1809 -1308 1815 1308
rect 1849 -1308 1855 1308
rect 1809 -1320 1855 -1308
rect 2267 1308 2313 1320
rect 2267 -1308 2273 1308
rect 2307 -1308 2313 1308
rect 2267 -1320 2313 -1308
rect -2399 -1460 2399 -1454
rect -2399 -1494 -2387 -1460
rect 2387 -1494 2399 -1460
rect -2399 -1500 2399 -1494
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -2404 -1477 2404 1477
string parameters w 13.2 l 2 m 1 nf 10 diffcov 100 polycov 20 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 100 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
