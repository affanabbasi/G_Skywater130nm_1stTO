magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -360 340 360 374
rect -360 -340 -326 340
rect 326 -340 360 340
rect -360 -374 360 -340
<< nmoslvt >>
rect -200 -200 200 200
<< ndiff >>
rect -258 187 -200 200
rect -258 153 -246 187
rect -212 153 -200 187
rect -258 119 -200 153
rect -258 85 -246 119
rect -212 85 -200 119
rect -258 51 -200 85
rect -258 17 -246 51
rect -212 17 -200 51
rect -258 -17 -200 17
rect -258 -51 -246 -17
rect -212 -51 -200 -17
rect -258 -85 -200 -51
rect -258 -119 -246 -85
rect -212 -119 -200 -85
rect -258 -153 -200 -119
rect -258 -187 -246 -153
rect -212 -187 -200 -153
rect -258 -200 -200 -187
rect 200 187 258 200
rect 200 153 212 187
rect 246 153 258 187
rect 200 119 258 153
rect 200 85 212 119
rect 246 85 258 119
rect 200 51 258 85
rect 200 17 212 51
rect 246 17 258 51
rect 200 -17 258 17
rect 200 -51 212 -17
rect 246 -51 258 -17
rect 200 -85 258 -51
rect 200 -119 212 -85
rect 246 -119 258 -85
rect 200 -153 258 -119
rect 200 -187 212 -153
rect 246 -187 258 -153
rect 200 -200 258 -187
<< ndiffc >>
rect -246 153 -212 187
rect -246 85 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -85
rect -246 -187 -212 -153
rect 212 153 246 187
rect 212 85 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -85
rect 212 -187 246 -153
<< psubdiff >>
rect -360 340 -255 374
rect -221 340 -187 374
rect -153 340 -119 374
rect -85 340 -51 374
rect -17 340 17 374
rect 51 340 85 374
rect 119 340 153 374
rect 187 340 221 374
rect 255 340 360 374
rect -360 255 -326 340
rect -360 187 -326 221
rect 326 255 360 340
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
rect 326 187 360 221
rect 326 119 360 153
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect 326 -153 360 -119
rect -360 -340 -326 -255
rect 326 -221 360 -187
rect 326 -340 360 -255
rect -360 -374 -255 -340
rect -221 -374 -187 -340
rect -153 -374 -119 -340
rect -85 -374 -51 -340
rect -17 -374 17 -340
rect 51 -374 85 -340
rect 119 -374 153 -340
rect 187 -374 221 -340
rect 255 -374 360 -340
<< psubdiffcont >>
rect -255 340 -221 374
rect -187 340 -153 374
rect -119 340 -85 374
rect -51 340 -17 374
rect 17 340 51 374
rect 85 340 119 374
rect 153 340 187 374
rect 221 340 255 374
rect -360 221 -326 255
rect 326 221 360 255
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect 326 153 360 187
rect 326 85 360 119
rect 326 17 360 51
rect 326 -51 360 -17
rect 326 -119 360 -85
rect 326 -187 360 -153
rect -360 -255 -326 -221
rect 326 -255 360 -221
rect -255 -374 -221 -340
rect -187 -374 -153 -340
rect -119 -374 -85 -340
rect -51 -374 -17 -340
rect 17 -374 51 -340
rect 85 -374 119 -340
rect 153 -374 187 -340
rect 221 -374 255 -340
<< poly >>
rect -200 272 200 288
rect -200 238 -153 272
rect -119 238 -85 272
rect -51 238 -17 272
rect 17 238 51 272
rect 85 238 119 272
rect 153 238 200 272
rect -200 200 200 238
rect -200 -238 200 -200
rect -200 -272 -153 -238
rect -119 -272 -85 -238
rect -51 -272 -17 -238
rect 17 -272 51 -238
rect 85 -272 119 -238
rect 153 -272 200 -238
rect -200 -288 200 -272
<< polycont >>
rect -153 238 -119 272
rect -85 238 -51 272
rect -17 238 17 272
rect 51 238 85 272
rect 119 238 153 272
rect -153 -272 -119 -238
rect -85 -272 -51 -238
rect -17 -272 17 -238
rect 51 -272 85 -238
rect 119 -272 153 -238
<< locali >>
rect -360 340 -255 374
rect -221 340 -187 374
rect -153 340 -119 374
rect -85 340 -51 374
rect -17 340 17 374
rect 51 340 85 374
rect 119 340 153 374
rect 187 340 221 374
rect 255 340 360 374
rect -360 255 -326 340
rect -200 238 -153 272
rect -119 238 -85 272
rect -51 238 -17 272
rect 17 238 51 272
rect 85 238 119 272
rect 153 238 200 272
rect 326 255 360 340
rect -360 187 -326 221
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
rect -246 187 -212 204
rect -246 119 -212 153
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect -246 -153 -212 -119
rect -246 -204 -212 -187
rect 212 187 246 204
rect 212 119 246 153
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
rect 212 -153 246 -119
rect 212 -204 246 -187
rect 326 187 360 221
rect 326 119 360 153
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect 326 -153 360 -119
rect 326 -221 360 -187
rect -360 -340 -326 -255
rect -200 -272 -153 -238
rect -119 -272 -85 -238
rect -51 -272 -17 -238
rect 17 -272 51 -238
rect 85 -272 119 -238
rect 153 -272 200 -238
rect 326 -340 360 -255
rect -360 -374 -255 -340
rect -221 -374 -187 -340
rect -153 -374 -119 -340
rect -85 -374 -51 -340
rect -17 -374 17 -340
rect 51 -374 85 -340
rect 119 -374 153 -340
rect 187 -374 221 -340
rect 255 -374 360 -340
<< properties >>
string FIXED_BBOX -342 -356 342 356
<< end >>
