magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -642 838 642 872
rect -642 -838 -608 838
rect 608 -838 642 838
rect -642 -872 642 -838
<< psubdiff >>
rect -642 838 -527 872
rect -493 838 -459 872
rect -425 838 -391 872
rect -357 838 -323 872
rect -289 838 -255 872
rect -221 838 -187 872
rect -153 838 -119 872
rect -85 838 -51 872
rect -17 838 17 872
rect 51 838 85 872
rect 119 838 153 872
rect 187 838 221 872
rect 255 838 289 872
rect 323 838 357 872
rect 391 838 425 872
rect 459 838 493 872
rect 527 838 642 872
rect -642 765 -608 838
rect 608 765 642 838
rect -642 697 -608 731
rect -642 629 -608 663
rect -642 561 -608 595
rect -642 493 -608 527
rect -642 425 -608 459
rect -642 357 -608 391
rect -642 289 -608 323
rect -642 221 -608 255
rect -642 153 -608 187
rect -642 85 -608 119
rect -642 17 -608 51
rect -642 -51 -608 -17
rect -642 -119 -608 -85
rect -642 -187 -608 -153
rect -642 -255 -608 -221
rect -642 -323 -608 -289
rect -642 -391 -608 -357
rect -642 -459 -608 -425
rect -642 -527 -608 -493
rect -642 -595 -608 -561
rect -642 -663 -608 -629
rect -642 -731 -608 -697
rect 608 697 642 731
rect 608 629 642 663
rect 608 561 642 595
rect 608 493 642 527
rect 608 425 642 459
rect 608 357 642 391
rect 608 289 642 323
rect 608 221 642 255
rect 608 153 642 187
rect 608 85 642 119
rect 608 17 642 51
rect 608 -51 642 -17
rect 608 -119 642 -85
rect 608 -187 642 -153
rect 608 -255 642 -221
rect 608 -323 642 -289
rect 608 -391 642 -357
rect 608 -459 642 -425
rect 608 -527 642 -493
rect 608 -595 642 -561
rect 608 -663 642 -629
rect 608 -731 642 -697
rect -642 -838 -608 -765
rect 608 -838 642 -765
rect -642 -872 -527 -838
rect -493 -872 -459 -838
rect -425 -872 -391 -838
rect -357 -872 -323 -838
rect -289 -872 -255 -838
rect -221 -872 -187 -838
rect -153 -872 -119 -838
rect -85 -872 -51 -838
rect -17 -872 17 -838
rect 51 -872 85 -838
rect 119 -872 153 -838
rect 187 -872 221 -838
rect 255 -872 289 -838
rect 323 -872 357 -838
rect 391 -872 425 -838
rect 459 -872 493 -838
rect 527 -872 642 -838
<< psubdiffcont >>
rect -527 838 -493 872
rect -459 838 -425 872
rect -391 838 -357 872
rect -323 838 -289 872
rect -255 838 -221 872
rect -187 838 -153 872
rect -119 838 -85 872
rect -51 838 -17 872
rect 17 838 51 872
rect 85 838 119 872
rect 153 838 187 872
rect 221 838 255 872
rect 289 838 323 872
rect 357 838 391 872
rect 425 838 459 872
rect 493 838 527 872
rect -642 731 -608 765
rect -642 663 -608 697
rect -642 595 -608 629
rect -642 527 -608 561
rect -642 459 -608 493
rect -642 391 -608 425
rect -642 323 -608 357
rect -642 255 -608 289
rect -642 187 -608 221
rect -642 119 -608 153
rect -642 51 -608 85
rect -642 -17 -608 17
rect -642 -85 -608 -51
rect -642 -153 -608 -119
rect -642 -221 -608 -187
rect -642 -289 -608 -255
rect -642 -357 -608 -323
rect -642 -425 -608 -391
rect -642 -493 -608 -459
rect -642 -561 -608 -527
rect -642 -629 -608 -595
rect -642 -697 -608 -663
rect -642 -765 -608 -731
rect 608 731 642 765
rect 608 663 642 697
rect 608 595 642 629
rect 608 527 642 561
rect 608 459 642 493
rect 608 391 642 425
rect 608 323 642 357
rect 608 255 642 289
rect 608 187 642 221
rect 608 119 642 153
rect 608 51 642 85
rect 608 -17 642 17
rect 608 -85 642 -51
rect 608 -153 642 -119
rect 608 -221 642 -187
rect 608 -289 642 -255
rect 608 -357 642 -323
rect 608 -425 642 -391
rect 608 -493 642 -459
rect 608 -561 642 -527
rect 608 -629 642 -595
rect 608 -697 642 -663
rect 608 -765 642 -731
rect -527 -872 -493 -838
rect -459 -872 -425 -838
rect -391 -872 -357 -838
rect -323 -872 -289 -838
rect -255 -872 -221 -838
rect -187 -872 -153 -838
rect -119 -872 -85 -838
rect -51 -872 -17 -838
rect 17 -872 51 -838
rect 85 -872 119 -838
rect 153 -872 187 -838
rect 221 -872 255 -838
rect 289 -872 323 -838
rect 357 -872 391 -838
rect 425 -872 459 -838
rect 493 -872 527 -838
<< xpolycontact >>
rect -512 310 -442 742
rect -512 -742 -442 -310
rect -194 310 -124 742
rect -194 -742 -124 -310
rect 124 310 194 742
rect 124 -742 194 -310
rect 442 310 512 742
rect 442 -742 512 -310
<< xpolyres >>
rect -512 -310 -442 310
rect -194 -310 -124 310
rect 124 -310 194 310
rect 442 -310 512 310
<< locali >>
rect -642 838 -527 872
rect -493 838 -459 872
rect -425 838 -391 872
rect -357 838 -323 872
rect -289 838 -255 872
rect -221 838 -187 872
rect -153 838 -119 872
rect -85 838 -51 872
rect -17 838 17 872
rect 51 838 85 872
rect 119 838 153 872
rect 187 838 221 872
rect 255 838 289 872
rect 323 838 357 872
rect 391 838 425 872
rect 459 838 493 872
rect 527 838 642 872
rect -642 765 -608 838
rect 608 765 642 838
rect -642 697 -608 731
rect -642 629 -608 663
rect -642 561 -608 595
rect -642 493 -608 527
rect -642 425 -608 459
rect -642 357 -608 391
rect -642 289 -608 323
rect 608 697 642 731
rect 608 629 642 663
rect 608 561 642 595
rect 608 493 642 527
rect 608 425 642 459
rect 608 357 642 391
rect -642 221 -608 255
rect -642 153 -608 187
rect -642 85 -608 119
rect -642 17 -608 51
rect -642 -51 -608 -17
rect -642 -119 -608 -85
rect -642 -187 -608 -153
rect -642 -255 -608 -221
rect -642 -323 -608 -289
rect 608 289 642 323
rect 608 221 642 255
rect 608 153 642 187
rect 608 85 642 119
rect 608 17 642 51
rect 608 -51 642 -17
rect 608 -119 642 -85
rect 608 -187 642 -153
rect 608 -255 642 -221
rect -642 -391 -608 -357
rect -642 -459 -608 -425
rect -642 -527 -608 -493
rect -642 -595 -608 -561
rect -642 -663 -608 -629
rect -642 -731 -608 -697
rect 608 -323 642 -289
rect 608 -391 642 -357
rect 608 -459 642 -425
rect 608 -527 642 -493
rect 608 -595 642 -561
rect 608 -663 642 -629
rect 608 -731 642 -697
rect -642 -838 -608 -765
rect 608 -838 642 -765
rect -642 -872 -527 -838
rect -493 -872 -459 -838
rect -425 -872 -391 -838
rect -357 -872 -323 -838
rect -289 -872 -255 -838
rect -221 -872 -187 -838
rect -153 -872 -119 -838
rect -85 -872 -51 -838
rect -17 -872 17 -838
rect 51 -872 85 -838
rect 119 -872 153 -838
rect 187 -872 221 -838
rect 255 -872 289 -838
rect 323 -872 357 -838
rect 391 -872 425 -838
rect 459 -872 493 -838
rect 527 -872 642 -838
<< properties >>
string FIXED_BBOX -624 -854 624 854
<< end >>
