magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< error_p >>
rect -738 600 566 652
rect -738 552 -686 600
rect -666 552 494 580
rect -638 500 494 552
rect -638 -500 -586 500
rect 414 -500 494 500
rect -638 -552 494 -500
rect 466 -580 494 -552
rect 514 -600 566 600
rect 466 -652 566 -600
<< metal3 >>
rect -786 672 786 700
rect -786 608 702 672
rect 766 608 786 672
rect -786 600 786 608
rect -786 -600 -686 600
rect 514 592 786 600
rect 514 528 702 592
rect 766 528 786 592
rect 514 512 786 528
rect 514 448 702 512
rect 766 448 786 512
rect 514 432 786 448
rect 514 368 702 432
rect 766 368 786 432
rect 514 352 786 368
rect 514 288 702 352
rect 766 288 786 352
rect 514 272 786 288
rect 514 208 702 272
rect 766 208 786 272
rect 514 192 786 208
rect 514 128 702 192
rect 766 128 786 192
rect 514 112 786 128
rect 514 48 702 112
rect 766 48 786 112
rect 514 32 786 48
rect 514 -32 702 32
rect 766 -32 786 32
rect 514 -48 786 -32
rect 514 -112 702 -48
rect 766 -112 786 -48
rect 514 -128 786 -112
rect 514 -192 702 -128
rect 766 -192 786 -128
rect 514 -208 786 -192
rect 514 -272 702 -208
rect 766 -272 786 -208
rect 514 -288 786 -272
rect 514 -352 702 -288
rect 766 -352 786 -288
rect 514 -368 786 -352
rect 514 -432 702 -368
rect 766 -432 786 -368
rect 514 -448 786 -432
rect 514 -512 702 -448
rect 766 -512 786 -448
rect 514 -528 786 -512
rect 514 -592 702 -528
rect 766 -592 786 -528
rect 514 -600 786 -592
rect -786 -608 786 -600
rect -786 -672 702 -608
rect 766 -672 786 -608
rect -786 -700 786 -672
<< via3 >>
rect 702 608 766 672
rect 702 528 766 592
rect 702 448 766 512
rect 702 368 766 432
rect 702 288 766 352
rect 702 208 766 272
rect 702 128 766 192
rect 702 48 766 112
rect 702 -32 766 32
rect 702 -112 766 -48
rect 702 -192 766 -128
rect 702 -272 766 -208
rect 702 -352 766 -288
rect 702 -432 766 -368
rect 702 -512 766 -448
rect 702 -592 766 -528
rect 702 -672 766 -608
<< mimcapcontact >>
rect -638 -552 466 552
<< metal4 >>
rect 686 672 782 688
rect 686 608 702 672
rect 766 608 782 672
rect 686 592 782 608
rect -647 552 475 561
rect -647 -552 -638 552
rect 466 -552 475 552
rect -647 -561 475 -552
rect 686 528 702 592
rect 766 528 782 592
rect 686 512 782 528
rect 686 448 702 512
rect 766 448 782 512
rect 686 432 782 448
rect 686 368 702 432
rect 766 368 782 432
rect 686 352 782 368
rect 686 288 702 352
rect 766 288 782 352
rect 686 272 782 288
rect 686 208 702 272
rect 766 208 782 272
rect 686 192 782 208
rect 686 128 702 192
rect 766 128 782 192
rect 686 112 782 128
rect 686 48 702 112
rect 766 48 782 112
rect 686 32 782 48
rect 686 -32 702 32
rect 766 -32 782 32
rect 686 -48 782 -32
rect 686 -112 702 -48
rect 766 -112 782 -48
rect 686 -128 782 -112
rect 686 -192 702 -128
rect 766 -192 782 -128
rect 686 -208 782 -192
rect 686 -272 702 -208
rect 766 -272 782 -208
rect 686 -288 782 -272
rect 686 -352 702 -288
rect 766 -352 782 -288
rect 686 -368 782 -352
rect 686 -432 702 -368
rect 766 -432 782 -368
rect 686 -448 782 -432
rect 686 -512 702 -448
rect 766 -512 782 -448
rect 686 -528 782 -512
rect 686 -592 702 -528
rect 766 -592 782 -528
rect 686 -608 782 -592
rect 686 -672 702 -608
rect 766 -672 782 -608
rect 686 -688 782 -672
<< properties >>
string FIXED_BBOX -786 -700 614 700
<< end >>
