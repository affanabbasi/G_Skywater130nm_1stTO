magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect -396 -1219 396 1219
<< pmoslvt >>
rect -200 -1000 200 1000
<< pdiff >>
rect -258 969 -200 1000
rect -258 935 -246 969
rect -212 935 -200 969
rect -258 901 -200 935
rect -258 867 -246 901
rect -212 867 -200 901
rect -258 833 -200 867
rect -258 799 -246 833
rect -212 799 -200 833
rect -258 765 -200 799
rect -258 731 -246 765
rect -212 731 -200 765
rect -258 697 -200 731
rect -258 663 -246 697
rect -212 663 -200 697
rect -258 629 -200 663
rect -258 595 -246 629
rect -212 595 -200 629
rect -258 561 -200 595
rect -258 527 -246 561
rect -212 527 -200 561
rect -258 493 -200 527
rect -258 459 -246 493
rect -212 459 -200 493
rect -258 425 -200 459
rect -258 391 -246 425
rect -212 391 -200 425
rect -258 357 -200 391
rect -258 323 -246 357
rect -212 323 -200 357
rect -258 289 -200 323
rect -258 255 -246 289
rect -212 255 -200 289
rect -258 221 -200 255
rect -258 187 -246 221
rect -212 187 -200 221
rect -258 153 -200 187
rect -258 119 -246 153
rect -212 119 -200 153
rect -258 85 -200 119
rect -258 51 -246 85
rect -212 51 -200 85
rect -258 17 -200 51
rect -258 -17 -246 17
rect -212 -17 -200 17
rect -258 -51 -200 -17
rect -258 -85 -246 -51
rect -212 -85 -200 -51
rect -258 -119 -200 -85
rect -258 -153 -246 -119
rect -212 -153 -200 -119
rect -258 -187 -200 -153
rect -258 -221 -246 -187
rect -212 -221 -200 -187
rect -258 -255 -200 -221
rect -258 -289 -246 -255
rect -212 -289 -200 -255
rect -258 -323 -200 -289
rect -258 -357 -246 -323
rect -212 -357 -200 -323
rect -258 -391 -200 -357
rect -258 -425 -246 -391
rect -212 -425 -200 -391
rect -258 -459 -200 -425
rect -258 -493 -246 -459
rect -212 -493 -200 -459
rect -258 -527 -200 -493
rect -258 -561 -246 -527
rect -212 -561 -200 -527
rect -258 -595 -200 -561
rect -258 -629 -246 -595
rect -212 -629 -200 -595
rect -258 -663 -200 -629
rect -258 -697 -246 -663
rect -212 -697 -200 -663
rect -258 -731 -200 -697
rect -258 -765 -246 -731
rect -212 -765 -200 -731
rect -258 -799 -200 -765
rect -258 -833 -246 -799
rect -212 -833 -200 -799
rect -258 -867 -200 -833
rect -258 -901 -246 -867
rect -212 -901 -200 -867
rect -258 -935 -200 -901
rect -258 -969 -246 -935
rect -212 -969 -200 -935
rect -258 -1000 -200 -969
rect 200 969 258 1000
rect 200 935 212 969
rect 246 935 258 969
rect 200 901 258 935
rect 200 867 212 901
rect 246 867 258 901
rect 200 833 258 867
rect 200 799 212 833
rect 246 799 258 833
rect 200 765 258 799
rect 200 731 212 765
rect 246 731 258 765
rect 200 697 258 731
rect 200 663 212 697
rect 246 663 258 697
rect 200 629 258 663
rect 200 595 212 629
rect 246 595 258 629
rect 200 561 258 595
rect 200 527 212 561
rect 246 527 258 561
rect 200 493 258 527
rect 200 459 212 493
rect 246 459 258 493
rect 200 425 258 459
rect 200 391 212 425
rect 246 391 258 425
rect 200 357 258 391
rect 200 323 212 357
rect 246 323 258 357
rect 200 289 258 323
rect 200 255 212 289
rect 246 255 258 289
rect 200 221 258 255
rect 200 187 212 221
rect 246 187 258 221
rect 200 153 258 187
rect 200 119 212 153
rect 246 119 258 153
rect 200 85 258 119
rect 200 51 212 85
rect 246 51 258 85
rect 200 17 258 51
rect 200 -17 212 17
rect 246 -17 258 17
rect 200 -51 258 -17
rect 200 -85 212 -51
rect 246 -85 258 -51
rect 200 -119 258 -85
rect 200 -153 212 -119
rect 246 -153 258 -119
rect 200 -187 258 -153
rect 200 -221 212 -187
rect 246 -221 258 -187
rect 200 -255 258 -221
rect 200 -289 212 -255
rect 246 -289 258 -255
rect 200 -323 258 -289
rect 200 -357 212 -323
rect 246 -357 258 -323
rect 200 -391 258 -357
rect 200 -425 212 -391
rect 246 -425 258 -391
rect 200 -459 258 -425
rect 200 -493 212 -459
rect 246 -493 258 -459
rect 200 -527 258 -493
rect 200 -561 212 -527
rect 246 -561 258 -527
rect 200 -595 258 -561
rect 200 -629 212 -595
rect 246 -629 258 -595
rect 200 -663 258 -629
rect 200 -697 212 -663
rect 246 -697 258 -663
rect 200 -731 258 -697
rect 200 -765 212 -731
rect 246 -765 258 -731
rect 200 -799 258 -765
rect 200 -833 212 -799
rect 246 -833 258 -799
rect 200 -867 258 -833
rect 200 -901 212 -867
rect 246 -901 258 -867
rect 200 -935 258 -901
rect 200 -969 212 -935
rect 246 -969 258 -935
rect 200 -1000 258 -969
<< pdiffc >>
rect -246 935 -212 969
rect -246 867 -212 901
rect -246 799 -212 833
rect -246 731 -212 765
rect -246 663 -212 697
rect -246 595 -212 629
rect -246 527 -212 561
rect -246 459 -212 493
rect -246 391 -212 425
rect -246 323 -212 357
rect -246 255 -212 289
rect -246 187 -212 221
rect -246 119 -212 153
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect -246 -153 -212 -119
rect -246 -221 -212 -187
rect -246 -289 -212 -255
rect -246 -357 -212 -323
rect -246 -425 -212 -391
rect -246 -493 -212 -459
rect -246 -561 -212 -527
rect -246 -629 -212 -595
rect -246 -697 -212 -663
rect -246 -765 -212 -731
rect -246 -833 -212 -799
rect -246 -901 -212 -867
rect -246 -969 -212 -935
rect 212 935 246 969
rect 212 867 246 901
rect 212 799 246 833
rect 212 731 246 765
rect 212 663 246 697
rect 212 595 246 629
rect 212 527 246 561
rect 212 459 246 493
rect 212 391 246 425
rect 212 323 246 357
rect 212 255 246 289
rect 212 187 246 221
rect 212 119 246 153
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
rect 212 -153 246 -119
rect 212 -221 246 -187
rect 212 -289 246 -255
rect 212 -357 246 -323
rect 212 -425 246 -391
rect 212 -493 246 -459
rect 212 -561 246 -527
rect 212 -629 246 -595
rect 212 -697 246 -663
rect 212 -765 246 -731
rect 212 -833 246 -799
rect 212 -901 246 -867
rect 212 -969 246 -935
<< nsubdiff >>
rect -360 1149 -255 1183
rect -221 1149 -187 1183
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect 187 1149 221 1183
rect 255 1149 360 1183
rect -360 1071 -326 1149
rect -360 1003 -326 1037
rect 326 1071 360 1149
rect 326 1003 360 1037
rect -360 935 -326 969
rect -360 867 -326 901
rect -360 799 -326 833
rect -360 731 -326 765
rect -360 663 -326 697
rect -360 595 -326 629
rect -360 527 -326 561
rect -360 459 -326 493
rect -360 391 -326 425
rect -360 323 -326 357
rect -360 255 -326 289
rect -360 187 -326 221
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
rect -360 -289 -326 -255
rect -360 -357 -326 -323
rect -360 -425 -326 -391
rect -360 -493 -326 -459
rect -360 -561 -326 -527
rect -360 -629 -326 -595
rect -360 -697 -326 -663
rect -360 -765 -326 -731
rect -360 -833 -326 -799
rect -360 -901 -326 -867
rect -360 -969 -326 -935
rect 326 935 360 969
rect 326 867 360 901
rect 326 799 360 833
rect 326 731 360 765
rect 326 663 360 697
rect 326 595 360 629
rect 326 527 360 561
rect 326 459 360 493
rect 326 391 360 425
rect 326 323 360 357
rect 326 255 360 289
rect 326 187 360 221
rect 326 119 360 153
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect 326 -153 360 -119
rect 326 -221 360 -187
rect 326 -289 360 -255
rect 326 -357 360 -323
rect 326 -425 360 -391
rect 326 -493 360 -459
rect 326 -561 360 -527
rect 326 -629 360 -595
rect 326 -697 360 -663
rect 326 -765 360 -731
rect 326 -833 360 -799
rect 326 -901 360 -867
rect 326 -969 360 -935
rect -360 -1037 -326 -1003
rect -360 -1149 -326 -1071
rect 326 -1037 360 -1003
rect 326 -1149 360 -1071
rect -360 -1183 -255 -1149
rect -221 -1183 -187 -1149
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
rect 187 -1183 221 -1149
rect 255 -1183 360 -1149
<< nsubdiffcont >>
rect -255 1149 -221 1183
rect -187 1149 -153 1183
rect -119 1149 -85 1183
rect -51 1149 -17 1183
rect 17 1149 51 1183
rect 85 1149 119 1183
rect 153 1149 187 1183
rect 221 1149 255 1183
rect -360 1037 -326 1071
rect -360 969 -326 1003
rect 326 1037 360 1071
rect -360 901 -326 935
rect -360 833 -326 867
rect -360 765 -326 799
rect -360 697 -326 731
rect -360 629 -326 663
rect -360 561 -326 595
rect -360 493 -326 527
rect -360 425 -326 459
rect -360 357 -326 391
rect -360 289 -326 323
rect -360 221 -326 255
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect -360 -255 -326 -221
rect -360 -323 -326 -289
rect -360 -391 -326 -357
rect -360 -459 -326 -425
rect -360 -527 -326 -493
rect -360 -595 -326 -561
rect -360 -663 -326 -629
rect -360 -731 -326 -697
rect -360 -799 -326 -765
rect -360 -867 -326 -833
rect -360 -935 -326 -901
rect -360 -1003 -326 -969
rect 326 969 360 1003
rect 326 901 360 935
rect 326 833 360 867
rect 326 765 360 799
rect 326 697 360 731
rect 326 629 360 663
rect 326 561 360 595
rect 326 493 360 527
rect 326 425 360 459
rect 326 357 360 391
rect 326 289 360 323
rect 326 221 360 255
rect 326 153 360 187
rect 326 85 360 119
rect 326 17 360 51
rect 326 -51 360 -17
rect 326 -119 360 -85
rect 326 -187 360 -153
rect 326 -255 360 -221
rect 326 -323 360 -289
rect 326 -391 360 -357
rect 326 -459 360 -425
rect 326 -527 360 -493
rect 326 -595 360 -561
rect 326 -663 360 -629
rect 326 -731 360 -697
rect 326 -799 360 -765
rect 326 -867 360 -833
rect 326 -935 360 -901
rect -360 -1071 -326 -1037
rect 326 -1003 360 -969
rect 326 -1071 360 -1037
rect -255 -1183 -221 -1149
rect -187 -1183 -153 -1149
rect -119 -1183 -85 -1149
rect -51 -1183 -17 -1149
rect 17 -1183 51 -1149
rect 85 -1183 119 -1149
rect 153 -1183 187 -1149
rect 221 -1183 255 -1149
<< poly >>
rect -200 1081 200 1097
rect -200 1047 -153 1081
rect -119 1047 -85 1081
rect -51 1047 -17 1081
rect 17 1047 51 1081
rect 85 1047 119 1081
rect 153 1047 200 1081
rect -200 1000 200 1047
rect -200 -1047 200 -1000
rect -200 -1081 -153 -1047
rect -119 -1081 -85 -1047
rect -51 -1081 -17 -1047
rect 17 -1081 51 -1047
rect 85 -1081 119 -1047
rect 153 -1081 200 -1047
rect -200 -1097 200 -1081
<< polycont >>
rect -153 1047 -119 1081
rect -85 1047 -51 1081
rect -17 1047 17 1081
rect 51 1047 85 1081
rect 119 1047 153 1081
rect -153 -1081 -119 -1047
rect -85 -1081 -51 -1047
rect -17 -1081 17 -1047
rect 51 -1081 85 -1047
rect 119 -1081 153 -1047
<< locali >>
rect -360 1149 -255 1183
rect -221 1149 -187 1183
rect -153 1149 -119 1183
rect -85 1149 -51 1183
rect -17 1149 17 1183
rect 51 1149 85 1183
rect 119 1149 153 1183
rect 187 1149 221 1183
rect 255 1149 360 1183
rect -360 1071 -326 1149
rect -200 1047 -161 1081
rect -119 1047 -89 1081
rect -51 1047 -17 1081
rect 17 1047 51 1081
rect 89 1047 119 1081
rect 161 1047 200 1081
rect 326 1071 360 1149
rect -360 1003 -326 1037
rect -360 935 -326 969
rect -360 867 -326 901
rect -360 799 -326 833
rect -360 731 -326 765
rect -360 663 -326 697
rect -360 595 -326 629
rect -360 527 -326 561
rect -360 459 -326 493
rect -360 391 -326 425
rect -360 323 -326 357
rect -360 255 -326 289
rect -360 187 -326 221
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
rect -360 -289 -326 -255
rect -360 -357 -326 -323
rect -360 -425 -326 -391
rect -360 -493 -326 -459
rect -360 -561 -326 -527
rect -360 -629 -326 -595
rect -360 -697 -326 -663
rect -360 -765 -326 -731
rect -360 -833 -326 -799
rect -360 -901 -326 -867
rect -360 -969 -326 -935
rect -360 -1037 -326 -1003
rect -246 969 -212 1004
rect -246 901 -212 919
rect -246 833 -212 847
rect -246 765 -212 775
rect -246 697 -212 703
rect -246 629 -212 631
rect -246 593 -212 595
rect -246 521 -212 527
rect -246 449 -212 459
rect -246 377 -212 391
rect -246 305 -212 323
rect -246 233 -212 255
rect -246 161 -212 187
rect -246 89 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -89
rect -246 -187 -212 -161
rect -246 -255 -212 -233
rect -246 -323 -212 -305
rect -246 -391 -212 -377
rect -246 -459 -212 -449
rect -246 -527 -212 -521
rect -246 -595 -212 -593
rect -246 -631 -212 -629
rect -246 -703 -212 -697
rect -246 -775 -212 -765
rect -246 -847 -212 -833
rect -246 -919 -212 -901
rect -246 -1004 -212 -969
rect 212 969 246 1004
rect 212 901 246 919
rect 212 833 246 847
rect 212 765 246 775
rect 212 697 246 703
rect 212 629 246 631
rect 212 593 246 595
rect 212 521 246 527
rect 212 449 246 459
rect 212 377 246 391
rect 212 305 246 323
rect 212 233 246 255
rect 212 161 246 187
rect 212 89 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -89
rect 212 -187 246 -161
rect 212 -255 246 -233
rect 212 -323 246 -305
rect 212 -391 246 -377
rect 212 -459 246 -449
rect 212 -527 246 -521
rect 212 -595 246 -593
rect 212 -631 246 -629
rect 212 -703 246 -697
rect 212 -775 246 -765
rect 212 -847 246 -833
rect 212 -919 246 -901
rect 212 -1004 246 -969
rect 326 1003 360 1037
rect 326 935 360 969
rect 326 867 360 901
rect 326 799 360 833
rect 326 731 360 765
rect 326 663 360 697
rect 326 595 360 629
rect 326 527 360 561
rect 326 459 360 493
rect 326 391 360 425
rect 326 323 360 357
rect 326 255 360 289
rect 326 187 360 221
rect 326 119 360 153
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect 326 -153 360 -119
rect 326 -221 360 -187
rect 326 -289 360 -255
rect 326 -357 360 -323
rect 326 -425 360 -391
rect 326 -493 360 -459
rect 326 -561 360 -527
rect 326 -629 360 -595
rect 326 -697 360 -663
rect 326 -765 360 -731
rect 326 -833 360 -799
rect 326 -901 360 -867
rect 326 -969 360 -935
rect 326 -1037 360 -1003
rect -360 -1149 -326 -1071
rect -200 -1081 -161 -1047
rect -119 -1081 -89 -1047
rect -51 -1081 -17 -1047
rect 17 -1081 51 -1047
rect 89 -1081 119 -1047
rect 161 -1081 200 -1047
rect 326 -1149 360 -1071
rect -360 -1183 -255 -1149
rect -221 -1183 -187 -1149
rect -153 -1183 -119 -1149
rect -85 -1183 -51 -1149
rect -17 -1183 17 -1149
rect 51 -1183 85 -1149
rect 119 -1183 153 -1149
rect 187 -1183 221 -1149
rect 255 -1183 360 -1149
<< viali >>
rect -161 1047 -153 1081
rect -153 1047 -127 1081
rect -89 1047 -85 1081
rect -85 1047 -55 1081
rect -17 1047 17 1081
rect 55 1047 85 1081
rect 85 1047 89 1081
rect 127 1047 153 1081
rect 153 1047 161 1081
rect -246 935 -212 953
rect -246 919 -212 935
rect -246 867 -212 881
rect -246 847 -212 867
rect -246 799 -212 809
rect -246 775 -212 799
rect -246 731 -212 737
rect -246 703 -212 731
rect -246 663 -212 665
rect -246 631 -212 663
rect -246 561 -212 593
rect -246 559 -212 561
rect -246 493 -212 521
rect -246 487 -212 493
rect -246 425 -212 449
rect -246 415 -212 425
rect -246 357 -212 377
rect -246 343 -212 357
rect -246 289 -212 305
rect -246 271 -212 289
rect -246 221 -212 233
rect -246 199 -212 221
rect -246 153 -212 161
rect -246 127 -212 153
rect -246 85 -212 89
rect -246 55 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -55
rect -246 -89 -212 -85
rect -246 -153 -212 -127
rect -246 -161 -212 -153
rect -246 -221 -212 -199
rect -246 -233 -212 -221
rect -246 -289 -212 -271
rect -246 -305 -212 -289
rect -246 -357 -212 -343
rect -246 -377 -212 -357
rect -246 -425 -212 -415
rect -246 -449 -212 -425
rect -246 -493 -212 -487
rect -246 -521 -212 -493
rect -246 -561 -212 -559
rect -246 -593 -212 -561
rect -246 -663 -212 -631
rect -246 -665 -212 -663
rect -246 -731 -212 -703
rect -246 -737 -212 -731
rect -246 -799 -212 -775
rect -246 -809 -212 -799
rect -246 -867 -212 -847
rect -246 -881 -212 -867
rect -246 -935 -212 -919
rect -246 -953 -212 -935
rect 212 935 246 953
rect 212 919 246 935
rect 212 867 246 881
rect 212 847 246 867
rect 212 799 246 809
rect 212 775 246 799
rect 212 731 246 737
rect 212 703 246 731
rect 212 663 246 665
rect 212 631 246 663
rect 212 561 246 593
rect 212 559 246 561
rect 212 493 246 521
rect 212 487 246 493
rect 212 425 246 449
rect 212 415 246 425
rect 212 357 246 377
rect 212 343 246 357
rect 212 289 246 305
rect 212 271 246 289
rect 212 221 246 233
rect 212 199 246 221
rect 212 153 246 161
rect 212 127 246 153
rect 212 85 246 89
rect 212 55 246 85
rect 212 -17 246 17
rect 212 -85 246 -55
rect 212 -89 246 -85
rect 212 -153 246 -127
rect 212 -161 246 -153
rect 212 -221 246 -199
rect 212 -233 246 -221
rect 212 -289 246 -271
rect 212 -305 246 -289
rect 212 -357 246 -343
rect 212 -377 246 -357
rect 212 -425 246 -415
rect 212 -449 246 -425
rect 212 -493 246 -487
rect 212 -521 246 -493
rect 212 -561 246 -559
rect 212 -593 246 -561
rect 212 -663 246 -631
rect 212 -665 246 -663
rect 212 -731 246 -703
rect 212 -737 246 -731
rect 212 -799 246 -775
rect 212 -809 246 -799
rect 212 -867 246 -847
rect 212 -881 246 -867
rect 212 -935 246 -919
rect 212 -953 246 -935
rect -161 -1081 -153 -1047
rect -153 -1081 -127 -1047
rect -89 -1081 -85 -1047
rect -85 -1081 -55 -1047
rect -17 -1081 17 -1047
rect 55 -1081 85 -1047
rect 85 -1081 89 -1047
rect 127 -1081 153 -1047
rect 153 -1081 161 -1047
<< metal1 >>
rect -196 1081 196 1087
rect -196 1047 -161 1081
rect -127 1047 -89 1081
rect -55 1047 -17 1081
rect 17 1047 55 1081
rect 89 1047 127 1081
rect 161 1047 196 1081
rect -196 1041 196 1047
rect -252 953 -206 1000
rect -252 919 -246 953
rect -212 919 -206 953
rect -252 881 -206 919
rect -252 847 -246 881
rect -212 847 -206 881
rect -252 809 -206 847
rect -252 775 -246 809
rect -212 775 -206 809
rect -252 737 -206 775
rect -252 703 -246 737
rect -212 703 -206 737
rect -252 665 -206 703
rect -252 631 -246 665
rect -212 631 -206 665
rect -252 593 -206 631
rect -252 559 -246 593
rect -212 559 -206 593
rect -252 521 -206 559
rect -252 487 -246 521
rect -212 487 -206 521
rect -252 449 -206 487
rect -252 415 -246 449
rect -212 415 -206 449
rect -252 377 -206 415
rect -252 343 -246 377
rect -212 343 -206 377
rect -252 305 -206 343
rect -252 271 -246 305
rect -212 271 -206 305
rect -252 233 -206 271
rect -252 199 -246 233
rect -212 199 -206 233
rect -252 161 -206 199
rect -252 127 -246 161
rect -212 127 -206 161
rect -252 89 -206 127
rect -252 55 -246 89
rect -212 55 -206 89
rect -252 17 -206 55
rect -252 -17 -246 17
rect -212 -17 -206 17
rect -252 -55 -206 -17
rect -252 -89 -246 -55
rect -212 -89 -206 -55
rect -252 -127 -206 -89
rect -252 -161 -246 -127
rect -212 -161 -206 -127
rect -252 -199 -206 -161
rect -252 -233 -246 -199
rect -212 -233 -206 -199
rect -252 -271 -206 -233
rect -252 -305 -246 -271
rect -212 -305 -206 -271
rect -252 -343 -206 -305
rect -252 -377 -246 -343
rect -212 -377 -206 -343
rect -252 -415 -206 -377
rect -252 -449 -246 -415
rect -212 -449 -206 -415
rect -252 -487 -206 -449
rect -252 -521 -246 -487
rect -212 -521 -206 -487
rect -252 -559 -206 -521
rect -252 -593 -246 -559
rect -212 -593 -206 -559
rect -252 -631 -206 -593
rect -252 -665 -246 -631
rect -212 -665 -206 -631
rect -252 -703 -206 -665
rect -252 -737 -246 -703
rect -212 -737 -206 -703
rect -252 -775 -206 -737
rect -252 -809 -246 -775
rect -212 -809 -206 -775
rect -252 -847 -206 -809
rect -252 -881 -246 -847
rect -212 -881 -206 -847
rect -252 -919 -206 -881
rect -252 -953 -246 -919
rect -212 -953 -206 -919
rect -252 -1000 -206 -953
rect 206 953 252 1000
rect 206 919 212 953
rect 246 919 252 953
rect 206 881 252 919
rect 206 847 212 881
rect 246 847 252 881
rect 206 809 252 847
rect 206 775 212 809
rect 246 775 252 809
rect 206 737 252 775
rect 206 703 212 737
rect 246 703 252 737
rect 206 665 252 703
rect 206 631 212 665
rect 246 631 252 665
rect 206 593 252 631
rect 206 559 212 593
rect 246 559 252 593
rect 206 521 252 559
rect 206 487 212 521
rect 246 487 252 521
rect 206 449 252 487
rect 206 415 212 449
rect 246 415 252 449
rect 206 377 252 415
rect 206 343 212 377
rect 246 343 252 377
rect 206 305 252 343
rect 206 271 212 305
rect 246 271 252 305
rect 206 233 252 271
rect 206 199 212 233
rect 246 199 252 233
rect 206 161 252 199
rect 206 127 212 161
rect 246 127 252 161
rect 206 89 252 127
rect 206 55 212 89
rect 246 55 252 89
rect 206 17 252 55
rect 206 -17 212 17
rect 246 -17 252 17
rect 206 -55 252 -17
rect 206 -89 212 -55
rect 246 -89 252 -55
rect 206 -127 252 -89
rect 206 -161 212 -127
rect 246 -161 252 -127
rect 206 -199 252 -161
rect 206 -233 212 -199
rect 246 -233 252 -199
rect 206 -271 252 -233
rect 206 -305 212 -271
rect 246 -305 252 -271
rect 206 -343 252 -305
rect 206 -377 212 -343
rect 246 -377 252 -343
rect 206 -415 252 -377
rect 206 -449 212 -415
rect 246 -449 252 -415
rect 206 -487 252 -449
rect 206 -521 212 -487
rect 246 -521 252 -487
rect 206 -559 252 -521
rect 206 -593 212 -559
rect 246 -593 252 -559
rect 206 -631 252 -593
rect 206 -665 212 -631
rect 246 -665 252 -631
rect 206 -703 252 -665
rect 206 -737 212 -703
rect 246 -737 252 -703
rect 206 -775 252 -737
rect 206 -809 212 -775
rect 246 -809 252 -775
rect 206 -847 252 -809
rect 206 -881 212 -847
rect 246 -881 252 -847
rect 206 -919 252 -881
rect 206 -953 212 -919
rect 246 -953 252 -919
rect 206 -1000 252 -953
rect -196 -1047 196 -1041
rect -196 -1081 -161 -1047
rect -127 -1081 -89 -1047
rect -55 -1081 -17 -1047
rect 17 -1081 55 -1047
rect 89 -1081 127 -1047
rect 161 -1081 196 -1047
rect -196 -1087 196 -1081
<< properties >>
string FIXED_BBOX -343 -1166 343 1166
<< end >>
