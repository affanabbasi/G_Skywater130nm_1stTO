magic
tech sky130A
magscale 1 2
timestamp 1608050792
<< nwell >>
rect -1083 -1219 1083 1219
<< pmoslvt >>
rect -887 -1000 -487 1000
rect -429 -1000 -29 1000
rect 29 -1000 429 1000
rect 487 -1000 887 1000
<< pdiff >>
rect -945 988 -887 1000
rect -945 -988 -933 988
rect -899 -988 -887 988
rect -945 -1000 -887 -988
rect -487 988 -429 1000
rect -487 -988 -475 988
rect -441 -988 -429 988
rect -487 -1000 -429 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 429 988 487 1000
rect 429 -988 441 988
rect 475 -988 487 988
rect 429 -1000 487 -988
rect 887 988 945 1000
rect 887 -988 899 988
rect 933 -988 945 988
rect 887 -1000 945 -988
<< pdiffc >>
rect -933 -988 -899 988
rect -475 -988 -441 988
rect -17 -988 17 988
rect 441 -988 475 988
rect 899 -988 933 988
<< nsubdiff >>
rect -1047 1149 -951 1183
rect 951 1149 1047 1183
rect -1047 1087 -1013 1149
rect 1013 1087 1047 1149
rect -1047 -1149 -1013 -1087
rect 1013 -1149 1047 -1087
rect -1047 -1183 -951 -1149
rect 951 -1183 1047 -1149
<< nsubdiffcont >>
rect -951 1149 951 1183
rect -1047 -1087 -1013 1087
rect 1013 -1087 1047 1087
rect -951 -1183 951 -1149
<< poly >>
rect -740 1081 -634 1097
rect -740 1064 -724 1081
rect -887 1047 -724 1064
rect -650 1064 -634 1081
rect -282 1081 -176 1097
rect -282 1064 -266 1081
rect -650 1047 -487 1064
rect -887 1000 -487 1047
rect -429 1047 -266 1064
rect -192 1064 -176 1081
rect 176 1081 282 1097
rect 176 1064 192 1081
rect -192 1047 -29 1064
rect -429 1000 -29 1047
rect 29 1047 192 1064
rect 266 1064 282 1081
rect 634 1081 740 1097
rect 634 1064 650 1081
rect 266 1047 429 1064
rect 29 1000 429 1047
rect 487 1047 650 1064
rect 724 1064 740 1081
rect 724 1047 887 1064
rect 487 1000 887 1047
rect -887 -1047 -487 -1000
rect -887 -1064 -724 -1047
rect -740 -1081 -724 -1064
rect -650 -1064 -487 -1047
rect -429 -1047 -29 -1000
rect -429 -1064 -266 -1047
rect -650 -1081 -634 -1064
rect -740 -1097 -634 -1081
rect -282 -1081 -266 -1064
rect -192 -1064 -29 -1047
rect 29 -1047 429 -1000
rect 29 -1064 192 -1047
rect -192 -1081 -176 -1064
rect -282 -1097 -176 -1081
rect 176 -1081 192 -1064
rect 266 -1064 429 -1047
rect 487 -1047 887 -1000
rect 487 -1064 650 -1047
rect 266 -1081 282 -1064
rect 176 -1097 282 -1081
rect 634 -1081 650 -1064
rect 724 -1064 887 -1047
rect 724 -1081 740 -1064
rect 634 -1097 740 -1081
<< polycont >>
rect -724 1047 -650 1081
rect -266 1047 -192 1081
rect 192 1047 266 1081
rect 650 1047 724 1081
rect -724 -1081 -650 -1047
rect -266 -1081 -192 -1047
rect 192 -1081 266 -1047
rect 650 -1081 724 -1047
<< locali >>
rect -1047 1087 -1013 1183
rect 1013 1087 1047 1183
rect -740 1047 -724 1081
rect -650 1047 -634 1081
rect -282 1047 -266 1081
rect -192 1047 -176 1081
rect 176 1047 192 1081
rect 266 1047 282 1081
rect 634 1047 650 1081
rect 724 1047 740 1081
rect -933 988 -899 1004
rect -933 -1004 -899 -988
rect -475 988 -441 1004
rect -475 -1004 -441 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 441 988 475 1004
rect 441 -1004 475 -988
rect 899 988 933 1004
rect 899 -1004 933 -988
rect -740 -1081 -724 -1047
rect -650 -1081 -634 -1047
rect -282 -1081 -266 -1047
rect -192 -1081 -176 -1047
rect 176 -1081 192 -1047
rect 266 -1081 282 -1047
rect 634 -1081 650 -1047
rect 724 -1081 740 -1047
rect -1047 -1149 -1013 -1087
rect 1013 -1149 1047 -1087
rect -1047 -1183 -951 -1149
rect 951 -1183 1047 -1149
<< viali >>
rect -1013 1149 -951 1183
rect -951 1149 951 1183
rect 951 1149 1013 1183
rect -933 -988 -899 988
rect -475 -988 -441 988
rect -17 -988 17 988
rect 441 -988 475 988
rect 899 -988 933 988
<< metal1 >>
rect -1025 1183 1025 1189
rect -1025 1149 -1013 1183
rect 1013 1149 1025 1183
rect -1025 1143 1025 1149
rect -939 988 -893 1000
rect -939 -988 -933 988
rect -899 -988 -893 988
rect -939 -1000 -893 -988
rect -481 988 -435 1000
rect -481 -988 -475 988
rect -441 -988 -435 988
rect -481 -1000 -435 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 435 988 481 1000
rect 435 -988 441 988
rect 475 -988 481 988
rect 435 -1000 481 -988
rect 893 988 939 1000
rect 893 -988 899 988
rect 933 -988 939 988
rect 893 -1000 939 -988
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -1030 -1166 1030 1166
string parameters w 10 l 2 m 1 nf 4 diffcov 100 polycov 20 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 100 viagb 0 viagate 0 viadrn 100 viasrc 100
string library sky130
<< end >>
