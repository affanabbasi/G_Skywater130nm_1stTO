magic
tech sky130A
magscale 1 2
timestamp 1607669338
<< error_p >>
rect 20 126 78 132
rect 20 92 32 126
rect 20 86 78 92
rect -76 -92 -18 -86
rect -76 -126 -64 -92
rect -76 -132 -18 -126
use sky130_fd_pr__nfet_01v8_M2KAWZ  sky130_fd_pr__nfet_01v8_M2KAWZ_0
timestamp 1607669338
transform 1 0 1 0 1 0
box -263 -264 263 264
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -210 -212 210 212
string parameters w 0.55 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1
string library sky130
<< end >>
