magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -1596 1528 1596 1562
rect -1596 -1528 -1562 1528
rect 1562 -1528 1596 1528
rect -1596 -1562 1596 -1528
<< psubdiff >>
rect -1596 1528 -1479 1562
rect -1445 1528 -1411 1562
rect -1377 1528 -1343 1562
rect -1309 1528 -1275 1562
rect -1241 1528 -1207 1562
rect -1173 1528 -1139 1562
rect -1105 1528 -1071 1562
rect -1037 1528 -1003 1562
rect -969 1528 -935 1562
rect -901 1528 -867 1562
rect -833 1528 -799 1562
rect -765 1528 -731 1562
rect -697 1528 -663 1562
rect -629 1528 -595 1562
rect -561 1528 -527 1562
rect -493 1528 -459 1562
rect -425 1528 -391 1562
rect -357 1528 -323 1562
rect -289 1528 -255 1562
rect -221 1528 -187 1562
rect -153 1528 -119 1562
rect -85 1528 -51 1562
rect -17 1528 17 1562
rect 51 1528 85 1562
rect 119 1528 153 1562
rect 187 1528 221 1562
rect 255 1528 289 1562
rect 323 1528 357 1562
rect 391 1528 425 1562
rect 459 1528 493 1562
rect 527 1528 561 1562
rect 595 1528 629 1562
rect 663 1528 697 1562
rect 731 1528 765 1562
rect 799 1528 833 1562
rect 867 1528 901 1562
rect 935 1528 969 1562
rect 1003 1528 1037 1562
rect 1071 1528 1105 1562
rect 1139 1528 1173 1562
rect 1207 1528 1241 1562
rect 1275 1528 1309 1562
rect 1343 1528 1377 1562
rect 1411 1528 1445 1562
rect 1479 1528 1596 1562
rect -1596 1445 -1562 1528
rect 1562 1445 1596 1528
rect -1596 1377 -1562 1411
rect -1596 1309 -1562 1343
rect -1596 1241 -1562 1275
rect -1596 1173 -1562 1207
rect -1596 1105 -1562 1139
rect -1596 1037 -1562 1071
rect -1596 969 -1562 1003
rect -1596 901 -1562 935
rect -1596 833 -1562 867
rect -1596 765 -1562 799
rect -1596 697 -1562 731
rect -1596 629 -1562 663
rect -1596 561 -1562 595
rect -1596 493 -1562 527
rect -1596 425 -1562 459
rect -1596 357 -1562 391
rect -1596 289 -1562 323
rect -1596 221 -1562 255
rect -1596 153 -1562 187
rect -1596 85 -1562 119
rect -1596 17 -1562 51
rect -1596 -51 -1562 -17
rect -1596 -119 -1562 -85
rect -1596 -187 -1562 -153
rect -1596 -255 -1562 -221
rect -1596 -323 -1562 -289
rect -1596 -391 -1562 -357
rect -1596 -459 -1562 -425
rect -1596 -527 -1562 -493
rect -1596 -595 -1562 -561
rect -1596 -663 -1562 -629
rect -1596 -731 -1562 -697
rect -1596 -799 -1562 -765
rect -1596 -867 -1562 -833
rect -1596 -935 -1562 -901
rect -1596 -1003 -1562 -969
rect -1596 -1071 -1562 -1037
rect -1596 -1139 -1562 -1105
rect -1596 -1207 -1562 -1173
rect -1596 -1275 -1562 -1241
rect -1596 -1343 -1562 -1309
rect -1596 -1411 -1562 -1377
rect 1562 1377 1596 1411
rect 1562 1309 1596 1343
rect 1562 1241 1596 1275
rect 1562 1173 1596 1207
rect 1562 1105 1596 1139
rect 1562 1037 1596 1071
rect 1562 969 1596 1003
rect 1562 901 1596 935
rect 1562 833 1596 867
rect 1562 765 1596 799
rect 1562 697 1596 731
rect 1562 629 1596 663
rect 1562 561 1596 595
rect 1562 493 1596 527
rect 1562 425 1596 459
rect 1562 357 1596 391
rect 1562 289 1596 323
rect 1562 221 1596 255
rect 1562 153 1596 187
rect 1562 85 1596 119
rect 1562 17 1596 51
rect 1562 -51 1596 -17
rect 1562 -119 1596 -85
rect 1562 -187 1596 -153
rect 1562 -255 1596 -221
rect 1562 -323 1596 -289
rect 1562 -391 1596 -357
rect 1562 -459 1596 -425
rect 1562 -527 1596 -493
rect 1562 -595 1596 -561
rect 1562 -663 1596 -629
rect 1562 -731 1596 -697
rect 1562 -799 1596 -765
rect 1562 -867 1596 -833
rect 1562 -935 1596 -901
rect 1562 -1003 1596 -969
rect 1562 -1071 1596 -1037
rect 1562 -1139 1596 -1105
rect 1562 -1207 1596 -1173
rect 1562 -1275 1596 -1241
rect 1562 -1343 1596 -1309
rect 1562 -1411 1596 -1377
rect -1596 -1528 -1562 -1445
rect 1562 -1528 1596 -1445
rect -1596 -1562 -1479 -1528
rect -1445 -1562 -1411 -1528
rect -1377 -1562 -1343 -1528
rect -1309 -1562 -1275 -1528
rect -1241 -1562 -1207 -1528
rect -1173 -1562 -1139 -1528
rect -1105 -1562 -1071 -1528
rect -1037 -1562 -1003 -1528
rect -969 -1562 -935 -1528
rect -901 -1562 -867 -1528
rect -833 -1562 -799 -1528
rect -765 -1562 -731 -1528
rect -697 -1562 -663 -1528
rect -629 -1562 -595 -1528
rect -561 -1562 -527 -1528
rect -493 -1562 -459 -1528
rect -425 -1562 -391 -1528
rect -357 -1562 -323 -1528
rect -289 -1562 -255 -1528
rect -221 -1562 -187 -1528
rect -153 -1562 -119 -1528
rect -85 -1562 -51 -1528
rect -17 -1562 17 -1528
rect 51 -1562 85 -1528
rect 119 -1562 153 -1528
rect 187 -1562 221 -1528
rect 255 -1562 289 -1528
rect 323 -1562 357 -1528
rect 391 -1562 425 -1528
rect 459 -1562 493 -1528
rect 527 -1562 561 -1528
rect 595 -1562 629 -1528
rect 663 -1562 697 -1528
rect 731 -1562 765 -1528
rect 799 -1562 833 -1528
rect 867 -1562 901 -1528
rect 935 -1562 969 -1528
rect 1003 -1562 1037 -1528
rect 1071 -1562 1105 -1528
rect 1139 -1562 1173 -1528
rect 1207 -1562 1241 -1528
rect 1275 -1562 1309 -1528
rect 1343 -1562 1377 -1528
rect 1411 -1562 1445 -1528
rect 1479 -1562 1596 -1528
<< psubdiffcont >>
rect -1479 1528 -1445 1562
rect -1411 1528 -1377 1562
rect -1343 1528 -1309 1562
rect -1275 1528 -1241 1562
rect -1207 1528 -1173 1562
rect -1139 1528 -1105 1562
rect -1071 1528 -1037 1562
rect -1003 1528 -969 1562
rect -935 1528 -901 1562
rect -867 1528 -833 1562
rect -799 1528 -765 1562
rect -731 1528 -697 1562
rect -663 1528 -629 1562
rect -595 1528 -561 1562
rect -527 1528 -493 1562
rect -459 1528 -425 1562
rect -391 1528 -357 1562
rect -323 1528 -289 1562
rect -255 1528 -221 1562
rect -187 1528 -153 1562
rect -119 1528 -85 1562
rect -51 1528 -17 1562
rect 17 1528 51 1562
rect 85 1528 119 1562
rect 153 1528 187 1562
rect 221 1528 255 1562
rect 289 1528 323 1562
rect 357 1528 391 1562
rect 425 1528 459 1562
rect 493 1528 527 1562
rect 561 1528 595 1562
rect 629 1528 663 1562
rect 697 1528 731 1562
rect 765 1528 799 1562
rect 833 1528 867 1562
rect 901 1528 935 1562
rect 969 1528 1003 1562
rect 1037 1528 1071 1562
rect 1105 1528 1139 1562
rect 1173 1528 1207 1562
rect 1241 1528 1275 1562
rect 1309 1528 1343 1562
rect 1377 1528 1411 1562
rect 1445 1528 1479 1562
rect -1596 1411 -1562 1445
rect -1596 1343 -1562 1377
rect -1596 1275 -1562 1309
rect -1596 1207 -1562 1241
rect -1596 1139 -1562 1173
rect -1596 1071 -1562 1105
rect -1596 1003 -1562 1037
rect -1596 935 -1562 969
rect -1596 867 -1562 901
rect -1596 799 -1562 833
rect -1596 731 -1562 765
rect -1596 663 -1562 697
rect -1596 595 -1562 629
rect -1596 527 -1562 561
rect -1596 459 -1562 493
rect -1596 391 -1562 425
rect -1596 323 -1562 357
rect -1596 255 -1562 289
rect -1596 187 -1562 221
rect -1596 119 -1562 153
rect -1596 51 -1562 85
rect -1596 -17 -1562 17
rect -1596 -85 -1562 -51
rect -1596 -153 -1562 -119
rect -1596 -221 -1562 -187
rect -1596 -289 -1562 -255
rect -1596 -357 -1562 -323
rect -1596 -425 -1562 -391
rect -1596 -493 -1562 -459
rect -1596 -561 -1562 -527
rect -1596 -629 -1562 -595
rect -1596 -697 -1562 -663
rect -1596 -765 -1562 -731
rect -1596 -833 -1562 -799
rect -1596 -901 -1562 -867
rect -1596 -969 -1562 -935
rect -1596 -1037 -1562 -1003
rect -1596 -1105 -1562 -1071
rect -1596 -1173 -1562 -1139
rect -1596 -1241 -1562 -1207
rect -1596 -1309 -1562 -1275
rect -1596 -1377 -1562 -1343
rect -1596 -1445 -1562 -1411
rect 1562 1411 1596 1445
rect 1562 1343 1596 1377
rect 1562 1275 1596 1309
rect 1562 1207 1596 1241
rect 1562 1139 1596 1173
rect 1562 1071 1596 1105
rect 1562 1003 1596 1037
rect 1562 935 1596 969
rect 1562 867 1596 901
rect 1562 799 1596 833
rect 1562 731 1596 765
rect 1562 663 1596 697
rect 1562 595 1596 629
rect 1562 527 1596 561
rect 1562 459 1596 493
rect 1562 391 1596 425
rect 1562 323 1596 357
rect 1562 255 1596 289
rect 1562 187 1596 221
rect 1562 119 1596 153
rect 1562 51 1596 85
rect 1562 -17 1596 17
rect 1562 -85 1596 -51
rect 1562 -153 1596 -119
rect 1562 -221 1596 -187
rect 1562 -289 1596 -255
rect 1562 -357 1596 -323
rect 1562 -425 1596 -391
rect 1562 -493 1596 -459
rect 1562 -561 1596 -527
rect 1562 -629 1596 -595
rect 1562 -697 1596 -663
rect 1562 -765 1596 -731
rect 1562 -833 1596 -799
rect 1562 -901 1596 -867
rect 1562 -969 1596 -935
rect 1562 -1037 1596 -1003
rect 1562 -1105 1596 -1071
rect 1562 -1173 1596 -1139
rect 1562 -1241 1596 -1207
rect 1562 -1309 1596 -1275
rect 1562 -1377 1596 -1343
rect 1562 -1445 1596 -1411
rect -1479 -1562 -1445 -1528
rect -1411 -1562 -1377 -1528
rect -1343 -1562 -1309 -1528
rect -1275 -1562 -1241 -1528
rect -1207 -1562 -1173 -1528
rect -1139 -1562 -1105 -1528
rect -1071 -1562 -1037 -1528
rect -1003 -1562 -969 -1528
rect -935 -1562 -901 -1528
rect -867 -1562 -833 -1528
rect -799 -1562 -765 -1528
rect -731 -1562 -697 -1528
rect -663 -1562 -629 -1528
rect -595 -1562 -561 -1528
rect -527 -1562 -493 -1528
rect -459 -1562 -425 -1528
rect -391 -1562 -357 -1528
rect -323 -1562 -289 -1528
rect -255 -1562 -221 -1528
rect -187 -1562 -153 -1528
rect -119 -1562 -85 -1528
rect -51 -1562 -17 -1528
rect 17 -1562 51 -1528
rect 85 -1562 119 -1528
rect 153 -1562 187 -1528
rect 221 -1562 255 -1528
rect 289 -1562 323 -1528
rect 357 -1562 391 -1528
rect 425 -1562 459 -1528
rect 493 -1562 527 -1528
rect 561 -1562 595 -1528
rect 629 -1562 663 -1528
rect 697 -1562 731 -1528
rect 765 -1562 799 -1528
rect 833 -1562 867 -1528
rect 901 -1562 935 -1528
rect 969 -1562 1003 -1528
rect 1037 -1562 1071 -1528
rect 1105 -1562 1139 -1528
rect 1173 -1562 1207 -1528
rect 1241 -1562 1275 -1528
rect 1309 -1562 1343 -1528
rect 1377 -1562 1411 -1528
rect 1445 -1562 1479 -1528
<< xpolycontact >>
rect -1466 1000 -1396 1432
rect -1466 -1432 -1396 -1000
rect -1148 1000 -1078 1432
rect -1148 -1432 -1078 -1000
rect -830 1000 -760 1432
rect -830 -1432 -760 -1000
rect -512 1000 -442 1432
rect -512 -1432 -442 -1000
rect -194 1000 -124 1432
rect -194 -1432 -124 -1000
rect 124 1000 194 1432
rect 124 -1432 194 -1000
rect 442 1000 512 1432
rect 442 -1432 512 -1000
rect 760 1000 830 1432
rect 760 -1432 830 -1000
rect 1078 1000 1148 1432
rect 1078 -1432 1148 -1000
rect 1396 1000 1466 1432
rect 1396 -1432 1466 -1000
<< ppolyres >>
rect -1466 -1000 -1396 1000
rect -1148 -1000 -1078 1000
rect -830 -1000 -760 1000
rect -512 -1000 -442 1000
rect -194 -1000 -124 1000
rect 124 -1000 194 1000
rect 442 -1000 512 1000
rect 760 -1000 830 1000
rect 1078 -1000 1148 1000
rect 1396 -1000 1466 1000
<< locali >>
rect -1596 1528 -1479 1562
rect -1445 1528 -1411 1562
rect -1377 1528 -1343 1562
rect -1309 1528 -1275 1562
rect -1241 1528 -1207 1562
rect -1173 1528 -1139 1562
rect -1105 1528 -1071 1562
rect -1037 1528 -1003 1562
rect -969 1528 -935 1562
rect -901 1528 -867 1562
rect -833 1528 -799 1562
rect -765 1528 -731 1562
rect -697 1528 -663 1562
rect -629 1528 -595 1562
rect -561 1528 -527 1562
rect -493 1528 -459 1562
rect -425 1528 -391 1562
rect -357 1528 -323 1562
rect -289 1528 -255 1562
rect -221 1528 -187 1562
rect -153 1528 -119 1562
rect -85 1528 -51 1562
rect -17 1528 17 1562
rect 51 1528 85 1562
rect 119 1528 153 1562
rect 187 1528 221 1562
rect 255 1528 289 1562
rect 323 1528 357 1562
rect 391 1528 425 1562
rect 459 1528 493 1562
rect 527 1528 561 1562
rect 595 1528 629 1562
rect 663 1528 697 1562
rect 731 1528 765 1562
rect 799 1528 833 1562
rect 867 1528 901 1562
rect 935 1528 969 1562
rect 1003 1528 1037 1562
rect 1071 1528 1105 1562
rect 1139 1528 1173 1562
rect 1207 1528 1241 1562
rect 1275 1528 1309 1562
rect 1343 1528 1377 1562
rect 1411 1528 1445 1562
rect 1479 1528 1596 1562
rect -1596 1445 -1562 1528
rect 1562 1445 1596 1528
rect -1596 1377 -1562 1411
rect -1596 1309 -1562 1343
rect -1596 1241 -1562 1275
rect -1596 1173 -1562 1207
rect -1596 1105 -1562 1139
rect -1596 1037 -1562 1071
rect -1596 969 -1562 1003
rect 1562 1377 1596 1411
rect 1562 1309 1596 1343
rect 1562 1241 1596 1275
rect 1562 1173 1596 1207
rect 1562 1105 1596 1139
rect 1562 1037 1596 1071
rect -1596 901 -1562 935
rect -1596 833 -1562 867
rect -1596 765 -1562 799
rect -1596 697 -1562 731
rect -1596 629 -1562 663
rect -1596 561 -1562 595
rect -1596 493 -1562 527
rect -1596 425 -1562 459
rect -1596 357 -1562 391
rect -1596 289 -1562 323
rect -1596 221 -1562 255
rect -1596 153 -1562 187
rect -1596 85 -1562 119
rect -1596 17 -1562 51
rect -1596 -51 -1562 -17
rect -1596 -119 -1562 -85
rect -1596 -187 -1562 -153
rect -1596 -255 -1562 -221
rect -1596 -323 -1562 -289
rect -1596 -391 -1562 -357
rect -1596 -459 -1562 -425
rect -1596 -527 -1562 -493
rect -1596 -595 -1562 -561
rect -1596 -663 -1562 -629
rect -1596 -731 -1562 -697
rect -1596 -799 -1562 -765
rect -1596 -867 -1562 -833
rect -1596 -935 -1562 -901
rect -1596 -1003 -1562 -969
rect 1562 969 1596 1003
rect 1562 901 1596 935
rect 1562 833 1596 867
rect 1562 765 1596 799
rect 1562 697 1596 731
rect 1562 629 1596 663
rect 1562 561 1596 595
rect 1562 493 1596 527
rect 1562 425 1596 459
rect 1562 357 1596 391
rect 1562 289 1596 323
rect 1562 221 1596 255
rect 1562 153 1596 187
rect 1562 85 1596 119
rect 1562 17 1596 51
rect 1562 -51 1596 -17
rect 1562 -119 1596 -85
rect 1562 -187 1596 -153
rect 1562 -255 1596 -221
rect 1562 -323 1596 -289
rect 1562 -391 1596 -357
rect 1562 -459 1596 -425
rect 1562 -527 1596 -493
rect 1562 -595 1596 -561
rect 1562 -663 1596 -629
rect 1562 -731 1596 -697
rect 1562 -799 1596 -765
rect 1562 -867 1596 -833
rect 1562 -935 1596 -901
rect -1596 -1071 -1562 -1037
rect -1596 -1139 -1562 -1105
rect -1596 -1207 -1562 -1173
rect -1596 -1275 -1562 -1241
rect -1596 -1343 -1562 -1309
rect -1596 -1411 -1562 -1377
rect 1562 -1003 1596 -969
rect 1562 -1071 1596 -1037
rect 1562 -1139 1596 -1105
rect 1562 -1207 1596 -1173
rect 1562 -1275 1596 -1241
rect 1562 -1343 1596 -1309
rect 1562 -1411 1596 -1377
rect -1596 -1528 -1562 -1445
rect 1562 -1528 1596 -1445
rect -1596 -1562 -1479 -1528
rect -1445 -1562 -1411 -1528
rect -1377 -1562 -1343 -1528
rect -1309 -1562 -1275 -1528
rect -1241 -1562 -1207 -1528
rect -1173 -1562 -1139 -1528
rect -1105 -1562 -1071 -1528
rect -1037 -1562 -1003 -1528
rect -969 -1562 -935 -1528
rect -901 -1562 -867 -1528
rect -833 -1562 -799 -1528
rect -765 -1562 -731 -1528
rect -697 -1562 -663 -1528
rect -629 -1562 -595 -1528
rect -561 -1562 -527 -1528
rect -493 -1562 -459 -1528
rect -425 -1562 -391 -1528
rect -357 -1562 -323 -1528
rect -289 -1562 -255 -1528
rect -221 -1562 -187 -1528
rect -153 -1562 -119 -1528
rect -85 -1562 -51 -1528
rect -17 -1562 17 -1528
rect 51 -1562 85 -1528
rect 119 -1562 153 -1528
rect 187 -1562 221 -1528
rect 255 -1562 289 -1528
rect 323 -1562 357 -1528
rect 391 -1562 425 -1528
rect 459 -1562 493 -1528
rect 527 -1562 561 -1528
rect 595 -1562 629 -1528
rect 663 -1562 697 -1528
rect 731 -1562 765 -1528
rect 799 -1562 833 -1528
rect 867 -1562 901 -1528
rect 935 -1562 969 -1528
rect 1003 -1562 1037 -1528
rect 1071 -1562 1105 -1528
rect 1139 -1562 1173 -1528
rect 1207 -1562 1241 -1528
rect 1275 -1562 1309 -1528
rect 1343 -1562 1377 -1528
rect 1411 -1562 1445 -1528
rect 1479 -1562 1596 -1528
<< properties >>
string FIXED_BBOX -1578 -1544 1578 1544
<< end >>
