magic
tech sky130A
magscale 1 2
timestamp 1608071797
<< nwell >>
rect -1770 -919 1770 919
<< pmos >>
rect -1574 -700 -1174 700
rect -1116 -700 -716 700
rect -658 -700 -258 700
rect -200 -700 200 700
rect 258 -700 658 700
rect 716 -700 1116 700
rect 1174 -700 1574 700
<< pdiff >>
rect -1632 138 -1574 700
rect -1632 -138 -1620 138
rect -1586 -138 -1574 138
rect -1632 -700 -1574 -138
rect -1174 138 -1116 700
rect -1174 -138 -1162 138
rect -1128 -138 -1116 138
rect -1174 -700 -1116 -138
rect -716 138 -658 700
rect -716 -138 -704 138
rect -670 -138 -658 138
rect -716 -700 -658 -138
rect -258 138 -200 700
rect -258 -138 -246 138
rect -212 -138 -200 138
rect -258 -700 -200 -138
rect 200 138 258 700
rect 200 -138 212 138
rect 246 -138 258 138
rect 200 -700 258 -138
rect 658 138 716 700
rect 658 -138 670 138
rect 704 -138 716 138
rect 658 -700 716 -138
rect 1116 138 1174 700
rect 1116 -138 1128 138
rect 1162 -138 1174 138
rect 1116 -700 1174 -138
rect 1574 138 1632 700
rect 1574 -138 1586 138
rect 1620 -138 1632 138
rect 1574 -700 1632 -138
<< pdiffc >>
rect -1620 -138 -1586 138
rect -1162 -138 -1128 138
rect -704 -138 -670 138
rect -246 -138 -212 138
rect 212 -138 246 138
rect 670 -138 704 138
rect 1128 -138 1162 138
rect 1586 -138 1620 138
<< nsubdiff >>
rect -1734 849 -1638 883
rect 1638 849 1734 883
rect -1734 787 -1700 849
rect 1700 787 1734 849
rect -1734 -849 -1700 -787
rect 1700 -849 1734 -787
rect -1734 -883 -1638 -849
rect 1638 -883 1734 -849
<< nsubdiffcont >>
rect -1638 849 1638 883
rect -1734 -787 -1700 787
rect 1700 -787 1734 787
rect -1638 -883 1638 -849
<< poly >>
rect -1427 781 -1321 797
rect -1427 764 -1411 781
rect -1574 747 -1411 764
rect -1337 764 -1321 781
rect -969 781 -863 797
rect -969 764 -953 781
rect -1337 747 -1174 764
rect -1574 700 -1174 747
rect -1116 747 -953 764
rect -879 764 -863 781
rect -511 781 -405 797
rect -511 764 -495 781
rect -879 747 -716 764
rect -1116 700 -716 747
rect -658 747 -495 764
rect -421 764 -405 781
rect -53 781 53 797
rect -53 764 -37 781
rect -421 747 -258 764
rect -658 700 -258 747
rect -200 747 -37 764
rect 37 764 53 781
rect 405 781 511 797
rect 405 764 421 781
rect 37 747 200 764
rect -200 700 200 747
rect 258 747 421 764
rect 495 764 511 781
rect 863 781 969 797
rect 863 764 879 781
rect 495 747 658 764
rect 258 700 658 747
rect 716 747 879 764
rect 953 764 969 781
rect 1321 781 1427 797
rect 1321 764 1337 781
rect 953 747 1116 764
rect 716 700 1116 747
rect 1174 747 1337 764
rect 1411 764 1427 781
rect 1411 747 1574 764
rect 1174 700 1574 747
rect -1574 -747 -1174 -700
rect -1574 -764 -1411 -747
rect -1427 -781 -1411 -764
rect -1337 -764 -1174 -747
rect -1116 -747 -716 -700
rect -1116 -764 -953 -747
rect -1337 -781 -1321 -764
rect -1427 -797 -1321 -781
rect -969 -781 -953 -764
rect -879 -764 -716 -747
rect -658 -747 -258 -700
rect -658 -764 -495 -747
rect -879 -781 -863 -764
rect -969 -797 -863 -781
rect -511 -781 -495 -764
rect -421 -764 -258 -747
rect -200 -747 200 -700
rect -200 -764 -37 -747
rect -421 -781 -405 -764
rect -511 -797 -405 -781
rect -53 -781 -37 -764
rect 37 -764 200 -747
rect 258 -747 658 -700
rect 258 -764 421 -747
rect 37 -781 53 -764
rect -53 -797 53 -781
rect 405 -781 421 -764
rect 495 -764 658 -747
rect 716 -747 1116 -700
rect 716 -764 879 -747
rect 495 -781 511 -764
rect 405 -797 511 -781
rect 863 -781 879 -764
rect 953 -764 1116 -747
rect 1174 -747 1574 -700
rect 1174 -764 1337 -747
rect 953 -781 969 -764
rect 863 -797 969 -781
rect 1321 -781 1337 -764
rect 1411 -764 1574 -747
rect 1411 -781 1427 -764
rect 1321 -797 1427 -781
<< polycont >>
rect -1411 747 -1337 781
rect -953 747 -879 781
rect -495 747 -421 781
rect -37 747 37 781
rect 421 747 495 781
rect 879 747 953 781
rect 1337 747 1411 781
rect -1411 -781 -1337 -747
rect -953 -781 -879 -747
rect -495 -781 -421 -747
rect -37 -781 37 -747
rect 421 -781 495 -747
rect 879 -781 953 -747
rect 1337 -781 1411 -747
<< locali >>
rect -1734 849 -1638 883
rect 1638 849 1734 883
rect -1734 787 -1700 849
rect 1700 787 1734 849
rect -1427 747 -1411 781
rect -1337 747 -1321 781
rect -969 747 -953 781
rect -879 747 -863 781
rect -511 747 -495 781
rect -421 747 -405 781
rect -53 747 -37 781
rect 37 747 53 781
rect 405 747 421 781
rect 495 747 511 781
rect 863 747 879 781
rect 953 747 969 781
rect 1321 747 1337 781
rect 1411 747 1427 781
rect -1620 138 -1586 154
rect -1620 -154 -1586 -138
rect -1162 138 -1128 154
rect -1162 -154 -1128 -138
rect -704 138 -670 154
rect -704 -154 -670 -138
rect -246 138 -212 154
rect -246 -154 -212 -138
rect 212 138 246 154
rect 212 -154 246 -138
rect 670 138 704 154
rect 670 -154 704 -138
rect 1128 138 1162 154
rect 1128 -154 1162 -138
rect 1586 138 1620 154
rect 1586 -154 1620 -138
rect -1427 -781 -1411 -747
rect -1337 -781 -1321 -747
rect -969 -781 -953 -747
rect -879 -781 -863 -747
rect -511 -781 -495 -747
rect -421 -781 -405 -747
rect -53 -781 -37 -747
rect 37 -781 53 -747
rect 405 -781 421 -747
rect 495 -781 511 -747
rect 863 -781 879 -747
rect 953 -781 969 -747
rect 1321 -781 1337 -747
rect 1411 -781 1427 -747
rect -1734 -849 -1700 -787
rect 1700 -849 1734 -787
rect -1734 -883 -1638 -849
rect 1638 -883 1734 -849
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1717 -866 1717 866
string parameters w 7 l 2 m 1 nf 7 diffcov 20 polycov 20 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 0 viadrn 0 viasrc 0
string library sky130
<< end >>
