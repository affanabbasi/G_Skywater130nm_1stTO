magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect -211 -319 211 319
<< pmos >>
rect -15 -100 15 100
<< pdiff >>
rect -73 85 -15 100
rect -73 51 -61 85
rect -27 51 -15 85
rect -73 17 -15 51
rect -73 -17 -61 17
rect -27 -17 -15 17
rect -73 -51 -15 -17
rect -73 -85 -61 -51
rect -27 -85 -15 -51
rect -73 -100 -15 -85
rect 15 85 73 100
rect 15 51 27 85
rect 61 51 73 85
rect 15 17 73 51
rect 15 -17 27 17
rect 61 -17 73 17
rect 15 -51 73 -17
rect 15 -85 27 -51
rect 61 -85 73 -51
rect 15 -100 73 -85
<< pdiffc >>
rect -61 51 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -51
rect 27 51 61 85
rect 27 -17 61 17
rect 27 -85 61 -51
<< nsubdiff >>
rect -175 249 -51 283
rect -17 249 17 283
rect 51 249 175 283
rect -175 187 -141 249
rect -175 119 -141 153
rect 141 187 175 249
rect 141 119 175 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -153 -141 -119
rect -175 -249 -141 -187
rect 141 -153 175 -119
rect 141 -249 175 -187
rect -175 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 175 -249
<< nsubdiffcont >>
rect -51 249 -17 283
rect 17 249 51 283
rect -175 153 -141 187
rect 141 153 175 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect -175 -187 -141 -153
rect 141 -187 175 -153
rect -51 -283 -17 -249
rect 17 -283 51 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -15 100 15 131
rect -15 -131 15 -100
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
<< polycont >>
rect -17 147 17 181
rect -17 -181 17 -147
<< locali >>
rect -175 249 -51 283
rect -17 249 17 283
rect 51 249 175 283
rect -175 187 -141 249
rect 141 187 175 249
rect -175 119 -141 153
rect -33 147 -17 181
rect 17 147 33 181
rect 141 119 175 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -61 85 -27 104
rect -61 17 -27 51
rect -61 -51 -27 -17
rect -61 -104 -27 -85
rect 27 85 61 104
rect 27 17 61 51
rect 27 -51 61 -17
rect 27 -104 61 -85
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -153 -141 -119
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect 141 -153 175 -119
rect -175 -249 -141 -187
rect 141 -249 175 -187
rect -175 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 175 -249
<< properties >>
string FIXED_BBOX -158 -266 158 266
<< end >>
