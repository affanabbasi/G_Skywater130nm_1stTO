magic
tech sky130A
timestamp 1606508276
<< pwell >>
rect -105 -126 105 126
<< nmos >>
rect -7 -21 7 21
<< ndiff >>
rect -36 15 -7 21
rect -36 -15 -30 15
rect -13 -15 -7 15
rect -36 -21 -7 -15
rect 7 15 36 21
rect 7 -15 13 15
rect 30 -15 36 15
rect 7 -21 36 -15
<< ndiffc >>
rect -30 -15 -13 15
rect 13 -15 30 15
<< psubdiff >>
rect -87 91 -39 108
rect 39 91 87 108
rect -87 60 -70 91
rect 70 60 87 91
rect -87 -91 -70 -60
rect 70 -91 87 -60
rect -87 -108 -39 -91
rect 39 -108 87 -91
<< psubdiffcont >>
rect -39 91 39 108
rect -87 -60 -70 60
rect 70 -60 87 60
rect -39 -108 39 -91
<< poly >>
rect -16 57 16 65
rect -16 40 -8 57
rect 8 40 16 57
rect -16 32 16 40
rect -7 21 7 32
rect -7 -32 7 -21
rect -16 -40 16 -32
rect -16 -57 -8 -40
rect 8 -57 16 -40
rect -16 -65 16 -57
<< polycont >>
rect -8 40 8 57
rect -8 -57 8 -40
<< locali >>
rect -87 91 -39 108
rect 39 91 87 108
rect -87 60 -70 91
rect 70 60 87 91
rect -16 40 -8 57
rect 8 40 16 57
rect -30 15 -13 23
rect -30 -23 -13 -15
rect 13 15 30 23
rect 13 -23 30 -15
rect -16 -57 -8 -40
rect 8 -57 16 -40
rect -87 -91 -70 -60
rect 70 -91 87 -60
rect -87 -108 -39 -91
rect 39 -108 87 -91
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -79 -99 79 99
string parameters w 0.420 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1
string library sky130
<< end >>
