magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect -696 -969 696 969
<< pmoslvt >>
rect -500 -750 500 750
<< pdiff >>
rect -558 731 -500 750
rect -558 697 -546 731
rect -512 697 -500 731
rect -558 663 -500 697
rect -558 629 -546 663
rect -512 629 -500 663
rect -558 595 -500 629
rect -558 561 -546 595
rect -512 561 -500 595
rect -558 527 -500 561
rect -558 493 -546 527
rect -512 493 -500 527
rect -558 459 -500 493
rect -558 425 -546 459
rect -512 425 -500 459
rect -558 391 -500 425
rect -558 357 -546 391
rect -512 357 -500 391
rect -558 323 -500 357
rect -558 289 -546 323
rect -512 289 -500 323
rect -558 255 -500 289
rect -558 221 -546 255
rect -512 221 -500 255
rect -558 187 -500 221
rect -558 153 -546 187
rect -512 153 -500 187
rect -558 119 -500 153
rect -558 85 -546 119
rect -512 85 -500 119
rect -558 51 -500 85
rect -558 17 -546 51
rect -512 17 -500 51
rect -558 -17 -500 17
rect -558 -51 -546 -17
rect -512 -51 -500 -17
rect -558 -85 -500 -51
rect -558 -119 -546 -85
rect -512 -119 -500 -85
rect -558 -153 -500 -119
rect -558 -187 -546 -153
rect -512 -187 -500 -153
rect -558 -221 -500 -187
rect -558 -255 -546 -221
rect -512 -255 -500 -221
rect -558 -289 -500 -255
rect -558 -323 -546 -289
rect -512 -323 -500 -289
rect -558 -357 -500 -323
rect -558 -391 -546 -357
rect -512 -391 -500 -357
rect -558 -425 -500 -391
rect -558 -459 -546 -425
rect -512 -459 -500 -425
rect -558 -493 -500 -459
rect -558 -527 -546 -493
rect -512 -527 -500 -493
rect -558 -561 -500 -527
rect -558 -595 -546 -561
rect -512 -595 -500 -561
rect -558 -629 -500 -595
rect -558 -663 -546 -629
rect -512 -663 -500 -629
rect -558 -697 -500 -663
rect -558 -731 -546 -697
rect -512 -731 -500 -697
rect -558 -750 -500 -731
rect 500 731 558 750
rect 500 697 512 731
rect 546 697 558 731
rect 500 663 558 697
rect 500 629 512 663
rect 546 629 558 663
rect 500 595 558 629
rect 500 561 512 595
rect 546 561 558 595
rect 500 527 558 561
rect 500 493 512 527
rect 546 493 558 527
rect 500 459 558 493
rect 500 425 512 459
rect 546 425 558 459
rect 500 391 558 425
rect 500 357 512 391
rect 546 357 558 391
rect 500 323 558 357
rect 500 289 512 323
rect 546 289 558 323
rect 500 255 558 289
rect 500 221 512 255
rect 546 221 558 255
rect 500 187 558 221
rect 500 153 512 187
rect 546 153 558 187
rect 500 119 558 153
rect 500 85 512 119
rect 546 85 558 119
rect 500 51 558 85
rect 500 17 512 51
rect 546 17 558 51
rect 500 -17 558 17
rect 500 -51 512 -17
rect 546 -51 558 -17
rect 500 -85 558 -51
rect 500 -119 512 -85
rect 546 -119 558 -85
rect 500 -153 558 -119
rect 500 -187 512 -153
rect 546 -187 558 -153
rect 500 -221 558 -187
rect 500 -255 512 -221
rect 546 -255 558 -221
rect 500 -289 558 -255
rect 500 -323 512 -289
rect 546 -323 558 -289
rect 500 -357 558 -323
rect 500 -391 512 -357
rect 546 -391 558 -357
rect 500 -425 558 -391
rect 500 -459 512 -425
rect 546 -459 558 -425
rect 500 -493 558 -459
rect 500 -527 512 -493
rect 546 -527 558 -493
rect 500 -561 558 -527
rect 500 -595 512 -561
rect 546 -595 558 -561
rect 500 -629 558 -595
rect 500 -663 512 -629
rect 546 -663 558 -629
rect 500 -697 558 -663
rect 500 -731 512 -697
rect 546 -731 558 -697
rect 500 -750 558 -731
<< pdiffc >>
rect -546 697 -512 731
rect -546 629 -512 663
rect -546 561 -512 595
rect -546 493 -512 527
rect -546 425 -512 459
rect -546 357 -512 391
rect -546 289 -512 323
rect -546 221 -512 255
rect -546 153 -512 187
rect -546 85 -512 119
rect -546 17 -512 51
rect -546 -51 -512 -17
rect -546 -119 -512 -85
rect -546 -187 -512 -153
rect -546 -255 -512 -221
rect -546 -323 -512 -289
rect -546 -391 -512 -357
rect -546 -459 -512 -425
rect -546 -527 -512 -493
rect -546 -595 -512 -561
rect -546 -663 -512 -629
rect -546 -731 -512 -697
rect 512 697 546 731
rect 512 629 546 663
rect 512 561 546 595
rect 512 493 546 527
rect 512 425 546 459
rect 512 357 546 391
rect 512 289 546 323
rect 512 221 546 255
rect 512 153 546 187
rect 512 85 546 119
rect 512 17 546 51
rect 512 -51 546 -17
rect 512 -119 546 -85
rect 512 -187 546 -153
rect 512 -255 546 -221
rect 512 -323 546 -289
rect 512 -391 546 -357
rect 512 -459 546 -425
rect 512 -527 546 -493
rect 512 -595 546 -561
rect 512 -663 546 -629
rect 512 -731 546 -697
<< nsubdiff >>
rect -660 899 -561 933
rect -527 899 -493 933
rect -459 899 -425 933
rect -391 899 -357 933
rect -323 899 -289 933
rect -255 899 -221 933
rect -187 899 -153 933
rect -119 899 -85 933
rect -51 899 -17 933
rect 17 899 51 933
rect 85 899 119 933
rect 153 899 187 933
rect 221 899 255 933
rect 289 899 323 933
rect 357 899 391 933
rect 425 899 459 933
rect 493 899 527 933
rect 561 899 660 933
rect -660 833 -626 899
rect -660 765 -626 799
rect 626 833 660 899
rect 626 765 660 799
rect -660 697 -626 731
rect -660 629 -626 663
rect -660 561 -626 595
rect -660 493 -626 527
rect -660 425 -626 459
rect -660 357 -626 391
rect -660 289 -626 323
rect -660 221 -626 255
rect -660 153 -626 187
rect -660 85 -626 119
rect -660 17 -626 51
rect -660 -51 -626 -17
rect -660 -119 -626 -85
rect -660 -187 -626 -153
rect -660 -255 -626 -221
rect -660 -323 -626 -289
rect -660 -391 -626 -357
rect -660 -459 -626 -425
rect -660 -527 -626 -493
rect -660 -595 -626 -561
rect -660 -663 -626 -629
rect -660 -731 -626 -697
rect 626 697 660 731
rect 626 629 660 663
rect 626 561 660 595
rect 626 493 660 527
rect 626 425 660 459
rect 626 357 660 391
rect 626 289 660 323
rect 626 221 660 255
rect 626 153 660 187
rect 626 85 660 119
rect 626 17 660 51
rect 626 -51 660 -17
rect 626 -119 660 -85
rect 626 -187 660 -153
rect 626 -255 660 -221
rect 626 -323 660 -289
rect 626 -391 660 -357
rect 626 -459 660 -425
rect 626 -527 660 -493
rect 626 -595 660 -561
rect 626 -663 660 -629
rect 626 -731 660 -697
rect -660 -799 -626 -765
rect -660 -899 -626 -833
rect 626 -799 660 -765
rect 626 -899 660 -833
rect -660 -933 -561 -899
rect -527 -933 -493 -899
rect -459 -933 -425 -899
rect -391 -933 -357 -899
rect -323 -933 -289 -899
rect -255 -933 -221 -899
rect -187 -933 -153 -899
rect -119 -933 -85 -899
rect -51 -933 -17 -899
rect 17 -933 51 -899
rect 85 -933 119 -899
rect 153 -933 187 -899
rect 221 -933 255 -899
rect 289 -933 323 -899
rect 357 -933 391 -899
rect 425 -933 459 -899
rect 493 -933 527 -899
rect 561 -933 660 -899
<< nsubdiffcont >>
rect -561 899 -527 933
rect -493 899 -459 933
rect -425 899 -391 933
rect -357 899 -323 933
rect -289 899 -255 933
rect -221 899 -187 933
rect -153 899 -119 933
rect -85 899 -51 933
rect -17 899 17 933
rect 51 899 85 933
rect 119 899 153 933
rect 187 899 221 933
rect 255 899 289 933
rect 323 899 357 933
rect 391 899 425 933
rect 459 899 493 933
rect 527 899 561 933
rect -660 799 -626 833
rect -660 731 -626 765
rect 626 799 660 833
rect -660 663 -626 697
rect -660 595 -626 629
rect -660 527 -626 561
rect -660 459 -626 493
rect -660 391 -626 425
rect -660 323 -626 357
rect -660 255 -626 289
rect -660 187 -626 221
rect -660 119 -626 153
rect -660 51 -626 85
rect -660 -17 -626 17
rect -660 -85 -626 -51
rect -660 -153 -626 -119
rect -660 -221 -626 -187
rect -660 -289 -626 -255
rect -660 -357 -626 -323
rect -660 -425 -626 -391
rect -660 -493 -626 -459
rect -660 -561 -626 -527
rect -660 -629 -626 -595
rect -660 -697 -626 -663
rect -660 -765 -626 -731
rect 626 731 660 765
rect 626 663 660 697
rect 626 595 660 629
rect 626 527 660 561
rect 626 459 660 493
rect 626 391 660 425
rect 626 323 660 357
rect 626 255 660 289
rect 626 187 660 221
rect 626 119 660 153
rect 626 51 660 85
rect 626 -17 660 17
rect 626 -85 660 -51
rect 626 -153 660 -119
rect 626 -221 660 -187
rect 626 -289 660 -255
rect 626 -357 660 -323
rect 626 -425 660 -391
rect 626 -493 660 -459
rect 626 -561 660 -527
rect 626 -629 660 -595
rect 626 -697 660 -663
rect -660 -833 -626 -799
rect 626 -765 660 -731
rect 626 -833 660 -799
rect -561 -933 -527 -899
rect -493 -933 -459 -899
rect -425 -933 -391 -899
rect -357 -933 -323 -899
rect -289 -933 -255 -899
rect -221 -933 -187 -899
rect -153 -933 -119 -899
rect -85 -933 -51 -899
rect -17 -933 17 -899
rect 51 -933 85 -899
rect 119 -933 153 -899
rect 187 -933 221 -899
rect 255 -933 289 -899
rect 323 -933 357 -899
rect 391 -933 425 -899
rect 459 -933 493 -899
rect 527 -933 561 -899
<< poly >>
rect -500 831 500 847
rect -500 797 -459 831
rect -425 797 -391 831
rect -357 797 -323 831
rect -289 797 -255 831
rect -221 797 -187 831
rect -153 797 -119 831
rect -85 797 -51 831
rect -17 797 17 831
rect 51 797 85 831
rect 119 797 153 831
rect 187 797 221 831
rect 255 797 289 831
rect 323 797 357 831
rect 391 797 425 831
rect 459 797 500 831
rect -500 750 500 797
rect -500 -797 500 -750
rect -500 -831 -459 -797
rect -425 -831 -391 -797
rect -357 -831 -323 -797
rect -289 -831 -255 -797
rect -221 -831 -187 -797
rect -153 -831 -119 -797
rect -85 -831 -51 -797
rect -17 -831 17 -797
rect 51 -831 85 -797
rect 119 -831 153 -797
rect 187 -831 221 -797
rect 255 -831 289 -797
rect 323 -831 357 -797
rect 391 -831 425 -797
rect 459 -831 500 -797
rect -500 -847 500 -831
<< polycont >>
rect -459 797 -425 831
rect -391 797 -357 831
rect -323 797 -289 831
rect -255 797 -221 831
rect -187 797 -153 831
rect -119 797 -85 831
rect -51 797 -17 831
rect 17 797 51 831
rect 85 797 119 831
rect 153 797 187 831
rect 221 797 255 831
rect 289 797 323 831
rect 357 797 391 831
rect 425 797 459 831
rect -459 -831 -425 -797
rect -391 -831 -357 -797
rect -323 -831 -289 -797
rect -255 -831 -221 -797
rect -187 -831 -153 -797
rect -119 -831 -85 -797
rect -51 -831 -17 -797
rect 17 -831 51 -797
rect 85 -831 119 -797
rect 153 -831 187 -797
rect 221 -831 255 -797
rect 289 -831 323 -797
rect 357 -831 391 -797
rect 425 -831 459 -797
<< locali >>
rect -660 899 -561 933
rect -527 899 -493 933
rect -459 899 -425 933
rect -391 899 -357 933
rect -323 899 -289 933
rect -255 899 -221 933
rect -187 899 -153 933
rect -119 899 -85 933
rect -51 899 -17 933
rect 17 899 51 933
rect 85 899 119 933
rect 153 899 187 933
rect 221 899 255 933
rect 289 899 323 933
rect 357 899 391 933
rect 425 899 459 933
rect 493 899 527 933
rect 561 899 660 933
rect -660 833 -626 899
rect 626 833 660 899
rect -660 765 -626 799
rect -500 797 -459 831
rect -415 797 -391 831
rect -343 797 -323 831
rect -271 797 -255 831
rect -199 797 -187 831
rect -127 797 -119 831
rect -55 797 -51 831
rect 51 797 55 831
rect 119 797 127 831
rect 187 797 199 831
rect 255 797 271 831
rect 323 797 343 831
rect 391 797 415 831
rect 459 797 500 831
rect 626 765 660 799
rect -660 697 -626 731
rect -660 629 -626 663
rect -660 561 -626 595
rect -660 493 -626 527
rect -660 425 -626 459
rect -660 357 -626 391
rect -660 289 -626 323
rect -660 221 -626 255
rect -660 153 -626 187
rect -660 85 -626 119
rect -660 17 -626 51
rect -660 -51 -626 -17
rect -660 -119 -626 -85
rect -660 -187 -626 -153
rect -660 -255 -626 -221
rect -660 -323 -626 -289
rect -660 -391 -626 -357
rect -660 -459 -626 -425
rect -660 -527 -626 -493
rect -660 -595 -626 -561
rect -660 -663 -626 -629
rect -660 -731 -626 -697
rect -546 737 -512 754
rect -546 665 -512 697
rect -546 595 -512 629
rect -546 527 -512 559
rect -546 459 -512 487
rect -546 391 -512 415
rect -546 323 -512 343
rect -546 255 -512 271
rect -546 187 -512 199
rect -546 119 -512 127
rect -546 51 -512 55
rect -546 -55 -512 -51
rect -546 -127 -512 -119
rect -546 -199 -512 -187
rect -546 -271 -512 -255
rect -546 -343 -512 -323
rect -546 -415 -512 -391
rect -546 -487 -512 -459
rect -546 -559 -512 -527
rect -546 -629 -512 -595
rect -546 -697 -512 -665
rect -546 -754 -512 -737
rect 512 737 546 754
rect 512 665 546 697
rect 512 595 546 629
rect 512 527 546 559
rect 512 459 546 487
rect 512 391 546 415
rect 512 323 546 343
rect 512 255 546 271
rect 512 187 546 199
rect 512 119 546 127
rect 512 51 546 55
rect 512 -55 546 -51
rect 512 -127 546 -119
rect 512 -199 546 -187
rect 512 -271 546 -255
rect 512 -343 546 -323
rect 512 -415 546 -391
rect 512 -487 546 -459
rect 512 -559 546 -527
rect 512 -629 546 -595
rect 512 -697 546 -665
rect 512 -754 546 -737
rect 626 697 660 731
rect 626 629 660 663
rect 626 561 660 595
rect 626 493 660 527
rect 626 425 660 459
rect 626 357 660 391
rect 626 289 660 323
rect 626 221 660 255
rect 626 153 660 187
rect 626 85 660 119
rect 626 17 660 51
rect 626 -51 660 -17
rect 626 -119 660 -85
rect 626 -187 660 -153
rect 626 -255 660 -221
rect 626 -323 660 -289
rect 626 -391 660 -357
rect 626 -459 660 -425
rect 626 -527 660 -493
rect 626 -595 660 -561
rect 626 -663 660 -629
rect 626 -731 660 -697
rect -660 -799 -626 -765
rect -500 -831 -459 -797
rect -415 -831 -391 -797
rect -343 -831 -323 -797
rect -271 -831 -255 -797
rect -199 -831 -187 -797
rect -127 -831 -119 -797
rect -55 -831 -51 -797
rect 51 -831 55 -797
rect 119 -831 127 -797
rect 187 -831 199 -797
rect 255 -831 271 -797
rect 323 -831 343 -797
rect 391 -831 415 -797
rect 459 -831 500 -797
rect 626 -799 660 -765
rect -660 -899 -626 -833
rect 626 -899 660 -833
rect -660 -933 -561 -899
rect -527 -933 -493 -899
rect -459 -933 -425 -899
rect -391 -933 -357 -899
rect -323 -933 -289 -899
rect -255 -933 -221 -899
rect -187 -933 -153 -899
rect -119 -933 -85 -899
rect -51 -933 -17 -899
rect 17 -933 51 -899
rect 85 -933 119 -899
rect 153 -933 187 -899
rect 221 -933 255 -899
rect 289 -933 323 -899
rect 357 -933 391 -899
rect 425 -933 459 -899
rect 493 -933 527 -899
rect 561 -933 660 -899
<< viali >>
rect -449 797 -425 831
rect -425 797 -415 831
rect -377 797 -357 831
rect -357 797 -343 831
rect -305 797 -289 831
rect -289 797 -271 831
rect -233 797 -221 831
rect -221 797 -199 831
rect -161 797 -153 831
rect -153 797 -127 831
rect -89 797 -85 831
rect -85 797 -55 831
rect -17 797 17 831
rect 55 797 85 831
rect 85 797 89 831
rect 127 797 153 831
rect 153 797 161 831
rect 199 797 221 831
rect 221 797 233 831
rect 271 797 289 831
rect 289 797 305 831
rect 343 797 357 831
rect 357 797 377 831
rect 415 797 425 831
rect 425 797 449 831
rect -546 731 -512 737
rect -546 703 -512 731
rect -546 663 -512 665
rect -546 631 -512 663
rect -546 561 -512 593
rect -546 559 -512 561
rect -546 493 -512 521
rect -546 487 -512 493
rect -546 425 -512 449
rect -546 415 -512 425
rect -546 357 -512 377
rect -546 343 -512 357
rect -546 289 -512 305
rect -546 271 -512 289
rect -546 221 -512 233
rect -546 199 -512 221
rect -546 153 -512 161
rect -546 127 -512 153
rect -546 85 -512 89
rect -546 55 -512 85
rect -546 -17 -512 17
rect -546 -85 -512 -55
rect -546 -89 -512 -85
rect -546 -153 -512 -127
rect -546 -161 -512 -153
rect -546 -221 -512 -199
rect -546 -233 -512 -221
rect -546 -289 -512 -271
rect -546 -305 -512 -289
rect -546 -357 -512 -343
rect -546 -377 -512 -357
rect -546 -425 -512 -415
rect -546 -449 -512 -425
rect -546 -493 -512 -487
rect -546 -521 -512 -493
rect -546 -561 -512 -559
rect -546 -593 -512 -561
rect -546 -663 -512 -631
rect -546 -665 -512 -663
rect -546 -731 -512 -703
rect -546 -737 -512 -731
rect 512 731 546 737
rect 512 703 546 731
rect 512 663 546 665
rect 512 631 546 663
rect 512 561 546 593
rect 512 559 546 561
rect 512 493 546 521
rect 512 487 546 493
rect 512 425 546 449
rect 512 415 546 425
rect 512 357 546 377
rect 512 343 546 357
rect 512 289 546 305
rect 512 271 546 289
rect 512 221 546 233
rect 512 199 546 221
rect 512 153 546 161
rect 512 127 546 153
rect 512 85 546 89
rect 512 55 546 85
rect 512 -17 546 17
rect 512 -85 546 -55
rect 512 -89 546 -85
rect 512 -153 546 -127
rect 512 -161 546 -153
rect 512 -221 546 -199
rect 512 -233 546 -221
rect 512 -289 546 -271
rect 512 -305 546 -289
rect 512 -357 546 -343
rect 512 -377 546 -357
rect 512 -425 546 -415
rect 512 -449 546 -425
rect 512 -493 546 -487
rect 512 -521 546 -493
rect 512 -561 546 -559
rect 512 -593 546 -561
rect 512 -663 546 -631
rect 512 -665 546 -663
rect 512 -731 546 -703
rect 512 -737 546 -731
rect -449 -831 -425 -797
rect -425 -831 -415 -797
rect -377 -831 -357 -797
rect -357 -831 -343 -797
rect -305 -831 -289 -797
rect -289 -831 -271 -797
rect -233 -831 -221 -797
rect -221 -831 -199 -797
rect -161 -831 -153 -797
rect -153 -831 -127 -797
rect -89 -831 -85 -797
rect -85 -831 -55 -797
rect -17 -831 17 -797
rect 55 -831 85 -797
rect 85 -831 89 -797
rect 127 -831 153 -797
rect 153 -831 161 -797
rect 199 -831 221 -797
rect 221 -831 233 -797
rect 271 -831 289 -797
rect 289 -831 305 -797
rect 343 -831 357 -797
rect 357 -831 377 -797
rect 415 -831 425 -797
rect 425 -831 449 -797
<< metal1 >>
rect -496 831 496 837
rect -496 797 -449 831
rect -415 797 -377 831
rect -343 797 -305 831
rect -271 797 -233 831
rect -199 797 -161 831
rect -127 797 -89 831
rect -55 797 -17 831
rect 17 797 55 831
rect 89 797 127 831
rect 161 797 199 831
rect 233 797 271 831
rect 305 797 343 831
rect 377 797 415 831
rect 449 797 496 831
rect -496 791 496 797
rect -552 737 -506 750
rect -552 703 -546 737
rect -512 703 -506 737
rect -552 665 -506 703
rect -552 631 -546 665
rect -512 631 -506 665
rect -552 593 -506 631
rect -552 559 -546 593
rect -512 559 -506 593
rect -552 521 -506 559
rect -552 487 -546 521
rect -512 487 -506 521
rect -552 449 -506 487
rect -552 415 -546 449
rect -512 415 -506 449
rect -552 377 -506 415
rect -552 343 -546 377
rect -512 343 -506 377
rect -552 305 -506 343
rect -552 271 -546 305
rect -512 271 -506 305
rect -552 233 -506 271
rect -552 199 -546 233
rect -512 199 -506 233
rect -552 161 -506 199
rect -552 127 -546 161
rect -512 127 -506 161
rect -552 89 -506 127
rect -552 55 -546 89
rect -512 55 -506 89
rect -552 17 -506 55
rect -552 -17 -546 17
rect -512 -17 -506 17
rect -552 -55 -506 -17
rect -552 -89 -546 -55
rect -512 -89 -506 -55
rect -552 -127 -506 -89
rect -552 -161 -546 -127
rect -512 -161 -506 -127
rect -552 -199 -506 -161
rect -552 -233 -546 -199
rect -512 -233 -506 -199
rect -552 -271 -506 -233
rect -552 -305 -546 -271
rect -512 -305 -506 -271
rect -552 -343 -506 -305
rect -552 -377 -546 -343
rect -512 -377 -506 -343
rect -552 -415 -506 -377
rect -552 -449 -546 -415
rect -512 -449 -506 -415
rect -552 -487 -506 -449
rect -552 -521 -546 -487
rect -512 -521 -506 -487
rect -552 -559 -506 -521
rect -552 -593 -546 -559
rect -512 -593 -506 -559
rect -552 -631 -506 -593
rect -552 -665 -546 -631
rect -512 -665 -506 -631
rect -552 -703 -506 -665
rect -552 -737 -546 -703
rect -512 -737 -506 -703
rect -552 -750 -506 -737
rect 506 737 552 750
rect 506 703 512 737
rect 546 703 552 737
rect 506 665 552 703
rect 506 631 512 665
rect 546 631 552 665
rect 506 593 552 631
rect 506 559 512 593
rect 546 559 552 593
rect 506 521 552 559
rect 506 487 512 521
rect 546 487 552 521
rect 506 449 552 487
rect 506 415 512 449
rect 546 415 552 449
rect 506 377 552 415
rect 506 343 512 377
rect 546 343 552 377
rect 506 305 552 343
rect 506 271 512 305
rect 546 271 552 305
rect 506 233 552 271
rect 506 199 512 233
rect 546 199 552 233
rect 506 161 552 199
rect 506 127 512 161
rect 546 127 552 161
rect 506 89 552 127
rect 506 55 512 89
rect 546 55 552 89
rect 506 17 552 55
rect 506 -17 512 17
rect 546 -17 552 17
rect 506 -55 552 -17
rect 506 -89 512 -55
rect 546 -89 552 -55
rect 506 -127 552 -89
rect 506 -161 512 -127
rect 546 -161 552 -127
rect 506 -199 552 -161
rect 506 -233 512 -199
rect 546 -233 552 -199
rect 506 -271 552 -233
rect 506 -305 512 -271
rect 546 -305 552 -271
rect 506 -343 552 -305
rect 506 -377 512 -343
rect 546 -377 552 -343
rect 506 -415 552 -377
rect 506 -449 512 -415
rect 546 -449 552 -415
rect 506 -487 552 -449
rect 506 -521 512 -487
rect 546 -521 552 -487
rect 506 -559 552 -521
rect 506 -593 512 -559
rect 546 -593 552 -559
rect 506 -631 552 -593
rect 506 -665 512 -631
rect 546 -665 552 -631
rect 506 -703 552 -665
rect 506 -737 512 -703
rect 546 -737 552 -703
rect 506 -750 552 -737
rect -496 -797 496 -791
rect -496 -831 -449 -797
rect -415 -831 -377 -797
rect -343 -831 -305 -797
rect -271 -831 -233 -797
rect -199 -831 -161 -797
rect -127 -831 -89 -797
rect -55 -831 -17 -797
rect 17 -831 55 -797
rect 89 -831 127 -797
rect 161 -831 199 -797
rect 233 -831 271 -797
rect 305 -831 343 -797
rect 377 -831 415 -797
rect 449 -831 496 -797
rect -496 -837 496 -831
<< properties >>
string FIXED_BBOX -643 -916 643 916
<< end >>
