magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -210 1249 210 1283
rect -210 -1249 -176 1249
rect 176 -1249 210 1249
rect -210 -1283 210 -1249
<< nmos >>
rect -50 109 50 1109
rect -50 -1109 50 -109
<< ndiff >>
rect -108 1068 -50 1109
rect -108 1034 -96 1068
rect -62 1034 -50 1068
rect -108 1000 -50 1034
rect -108 966 -96 1000
rect -62 966 -50 1000
rect -108 932 -50 966
rect -108 898 -96 932
rect -62 898 -50 932
rect -108 864 -50 898
rect -108 830 -96 864
rect -62 830 -50 864
rect -108 796 -50 830
rect -108 762 -96 796
rect -62 762 -50 796
rect -108 728 -50 762
rect -108 694 -96 728
rect -62 694 -50 728
rect -108 660 -50 694
rect -108 626 -96 660
rect -62 626 -50 660
rect -108 592 -50 626
rect -108 558 -96 592
rect -62 558 -50 592
rect -108 524 -50 558
rect -108 490 -96 524
rect -62 490 -50 524
rect -108 456 -50 490
rect -108 422 -96 456
rect -62 422 -50 456
rect -108 388 -50 422
rect -108 354 -96 388
rect -62 354 -50 388
rect -108 320 -50 354
rect -108 286 -96 320
rect -62 286 -50 320
rect -108 252 -50 286
rect -108 218 -96 252
rect -62 218 -50 252
rect -108 184 -50 218
rect -108 150 -96 184
rect -62 150 -50 184
rect -108 109 -50 150
rect 50 1068 108 1109
rect 50 1034 62 1068
rect 96 1034 108 1068
rect 50 1000 108 1034
rect 50 966 62 1000
rect 96 966 108 1000
rect 50 932 108 966
rect 50 898 62 932
rect 96 898 108 932
rect 50 864 108 898
rect 50 830 62 864
rect 96 830 108 864
rect 50 796 108 830
rect 50 762 62 796
rect 96 762 108 796
rect 50 728 108 762
rect 50 694 62 728
rect 96 694 108 728
rect 50 660 108 694
rect 50 626 62 660
rect 96 626 108 660
rect 50 592 108 626
rect 50 558 62 592
rect 96 558 108 592
rect 50 524 108 558
rect 50 490 62 524
rect 96 490 108 524
rect 50 456 108 490
rect 50 422 62 456
rect 96 422 108 456
rect 50 388 108 422
rect 50 354 62 388
rect 96 354 108 388
rect 50 320 108 354
rect 50 286 62 320
rect 96 286 108 320
rect 50 252 108 286
rect 50 218 62 252
rect 96 218 108 252
rect 50 184 108 218
rect 50 150 62 184
rect 96 150 108 184
rect 50 109 108 150
rect -108 -150 -50 -109
rect -108 -184 -96 -150
rect -62 -184 -50 -150
rect -108 -218 -50 -184
rect -108 -252 -96 -218
rect -62 -252 -50 -218
rect -108 -286 -50 -252
rect -108 -320 -96 -286
rect -62 -320 -50 -286
rect -108 -354 -50 -320
rect -108 -388 -96 -354
rect -62 -388 -50 -354
rect -108 -422 -50 -388
rect -108 -456 -96 -422
rect -62 -456 -50 -422
rect -108 -490 -50 -456
rect -108 -524 -96 -490
rect -62 -524 -50 -490
rect -108 -558 -50 -524
rect -108 -592 -96 -558
rect -62 -592 -50 -558
rect -108 -626 -50 -592
rect -108 -660 -96 -626
rect -62 -660 -50 -626
rect -108 -694 -50 -660
rect -108 -728 -96 -694
rect -62 -728 -50 -694
rect -108 -762 -50 -728
rect -108 -796 -96 -762
rect -62 -796 -50 -762
rect -108 -830 -50 -796
rect -108 -864 -96 -830
rect -62 -864 -50 -830
rect -108 -898 -50 -864
rect -108 -932 -96 -898
rect -62 -932 -50 -898
rect -108 -966 -50 -932
rect -108 -1000 -96 -966
rect -62 -1000 -50 -966
rect -108 -1034 -50 -1000
rect -108 -1068 -96 -1034
rect -62 -1068 -50 -1034
rect -108 -1109 -50 -1068
rect 50 -150 108 -109
rect 50 -184 62 -150
rect 96 -184 108 -150
rect 50 -218 108 -184
rect 50 -252 62 -218
rect 96 -252 108 -218
rect 50 -286 108 -252
rect 50 -320 62 -286
rect 96 -320 108 -286
rect 50 -354 108 -320
rect 50 -388 62 -354
rect 96 -388 108 -354
rect 50 -422 108 -388
rect 50 -456 62 -422
rect 96 -456 108 -422
rect 50 -490 108 -456
rect 50 -524 62 -490
rect 96 -524 108 -490
rect 50 -558 108 -524
rect 50 -592 62 -558
rect 96 -592 108 -558
rect 50 -626 108 -592
rect 50 -660 62 -626
rect 96 -660 108 -626
rect 50 -694 108 -660
rect 50 -728 62 -694
rect 96 -728 108 -694
rect 50 -762 108 -728
rect 50 -796 62 -762
rect 96 -796 108 -762
rect 50 -830 108 -796
rect 50 -864 62 -830
rect 96 -864 108 -830
rect 50 -898 108 -864
rect 50 -932 62 -898
rect 96 -932 108 -898
rect 50 -966 108 -932
rect 50 -1000 62 -966
rect 96 -1000 108 -966
rect 50 -1034 108 -1000
rect 50 -1068 62 -1034
rect 96 -1068 108 -1034
rect 50 -1109 108 -1068
<< ndiffc >>
rect -96 1034 -62 1068
rect -96 966 -62 1000
rect -96 898 -62 932
rect -96 830 -62 864
rect -96 762 -62 796
rect -96 694 -62 728
rect -96 626 -62 660
rect -96 558 -62 592
rect -96 490 -62 524
rect -96 422 -62 456
rect -96 354 -62 388
rect -96 286 -62 320
rect -96 218 -62 252
rect -96 150 -62 184
rect 62 1034 96 1068
rect 62 966 96 1000
rect 62 898 96 932
rect 62 830 96 864
rect 62 762 96 796
rect 62 694 96 728
rect 62 626 96 660
rect 62 558 96 592
rect 62 490 96 524
rect 62 422 96 456
rect 62 354 96 388
rect 62 286 96 320
rect 62 218 96 252
rect 62 150 96 184
rect -96 -184 -62 -150
rect -96 -252 -62 -218
rect -96 -320 -62 -286
rect -96 -388 -62 -354
rect -96 -456 -62 -422
rect -96 -524 -62 -490
rect -96 -592 -62 -558
rect -96 -660 -62 -626
rect -96 -728 -62 -694
rect -96 -796 -62 -762
rect -96 -864 -62 -830
rect -96 -932 -62 -898
rect -96 -1000 -62 -966
rect -96 -1068 -62 -1034
rect 62 -184 96 -150
rect 62 -252 96 -218
rect 62 -320 96 -286
rect 62 -388 96 -354
rect 62 -456 96 -422
rect 62 -524 96 -490
rect 62 -592 96 -558
rect 62 -660 96 -626
rect 62 -728 96 -694
rect 62 -796 96 -762
rect 62 -864 96 -830
rect 62 -932 96 -898
rect 62 -1000 96 -966
rect 62 -1068 96 -1034
<< psubdiff >>
rect -210 1249 -85 1283
rect -51 1249 -17 1283
rect 17 1249 51 1283
rect 85 1249 210 1283
rect -210 1173 -176 1249
rect -210 1105 -176 1139
rect 176 1173 210 1249
rect -210 1037 -176 1071
rect -210 969 -176 1003
rect -210 901 -176 935
rect -210 833 -176 867
rect -210 765 -176 799
rect -210 697 -176 731
rect -210 629 -176 663
rect -210 561 -176 595
rect -210 493 -176 527
rect -210 425 -176 459
rect -210 357 -176 391
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect 176 1105 210 1139
rect 176 1037 210 1071
rect 176 969 210 1003
rect 176 901 210 935
rect 176 833 210 867
rect 176 765 210 799
rect 176 697 210 731
rect 176 629 210 663
rect 176 561 210 595
rect 176 493 210 527
rect 176 425 210 459
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect -210 17 -176 51
rect 176 85 210 119
rect -210 -51 -176 -17
rect 176 17 210 51
rect -210 -119 -176 -85
rect 176 -51 210 -17
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect -210 -459 -176 -425
rect -210 -527 -176 -493
rect -210 -595 -176 -561
rect -210 -663 -176 -629
rect -210 -731 -176 -697
rect -210 -799 -176 -765
rect -210 -867 -176 -833
rect -210 -935 -176 -901
rect -210 -1003 -176 -969
rect -210 -1071 -176 -1037
rect -210 -1139 -176 -1105
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect 176 -391 210 -357
rect 176 -459 210 -425
rect 176 -527 210 -493
rect 176 -595 210 -561
rect 176 -663 210 -629
rect 176 -731 210 -697
rect 176 -799 210 -765
rect 176 -867 210 -833
rect 176 -935 210 -901
rect 176 -1003 210 -969
rect 176 -1071 210 -1037
rect -210 -1249 -176 -1173
rect 176 -1139 210 -1105
rect 176 -1249 210 -1173
rect -210 -1283 -85 -1249
rect -51 -1283 -17 -1249
rect 17 -1283 51 -1249
rect 85 -1283 210 -1249
<< psubdiffcont >>
rect -85 1249 -51 1283
rect -17 1249 17 1283
rect 51 1249 85 1283
rect -210 1139 -176 1173
rect 176 1139 210 1173
rect -210 1071 -176 1105
rect -210 1003 -176 1037
rect -210 935 -176 969
rect -210 867 -176 901
rect -210 799 -176 833
rect -210 731 -176 765
rect -210 663 -176 697
rect -210 595 -176 629
rect -210 527 -176 561
rect -210 459 -176 493
rect -210 391 -176 425
rect -210 323 -176 357
rect -210 255 -176 289
rect -210 187 -176 221
rect -210 119 -176 153
rect 176 1071 210 1105
rect 176 1003 210 1037
rect 176 935 210 969
rect 176 867 210 901
rect 176 799 210 833
rect 176 731 210 765
rect 176 663 210 697
rect 176 595 210 629
rect 176 527 210 561
rect 176 459 210 493
rect 176 391 210 425
rect 176 323 210 357
rect 176 255 210 289
rect 176 187 210 221
rect 176 119 210 153
rect -210 51 -176 85
rect 176 51 210 85
rect -210 -17 -176 17
rect 176 -17 210 17
rect -210 -85 -176 -51
rect 176 -85 210 -51
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect -210 -289 -176 -255
rect -210 -357 -176 -323
rect -210 -425 -176 -391
rect -210 -493 -176 -459
rect -210 -561 -176 -527
rect -210 -629 -176 -595
rect -210 -697 -176 -663
rect -210 -765 -176 -731
rect -210 -833 -176 -799
rect -210 -901 -176 -867
rect -210 -969 -176 -935
rect -210 -1037 -176 -1003
rect -210 -1105 -176 -1071
rect 176 -153 210 -119
rect 176 -221 210 -187
rect 176 -289 210 -255
rect 176 -357 210 -323
rect 176 -425 210 -391
rect 176 -493 210 -459
rect 176 -561 210 -527
rect 176 -629 210 -595
rect 176 -697 210 -663
rect 176 -765 210 -731
rect 176 -833 210 -799
rect 176 -901 210 -867
rect 176 -969 210 -935
rect 176 -1037 210 -1003
rect 176 -1105 210 -1071
rect -210 -1173 -176 -1139
rect 176 -1173 210 -1139
rect -85 -1283 -51 -1249
rect -17 -1283 17 -1249
rect 51 -1283 85 -1249
<< poly >>
rect -50 1181 50 1197
rect -50 1147 -17 1181
rect 17 1147 50 1181
rect -50 1109 50 1147
rect -50 71 50 109
rect -50 37 -17 71
rect 17 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -17 -37
rect 17 -71 50 -37
rect -50 -109 50 -71
rect -50 -1147 50 -1109
rect -50 -1181 -17 -1147
rect 17 -1181 50 -1147
rect -50 -1197 50 -1181
<< polycont >>
rect -17 1147 17 1181
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -1181 17 -1147
<< locali >>
rect -210 1249 -85 1283
rect -51 1249 -17 1283
rect 17 1249 51 1283
rect 85 1249 210 1283
rect -210 1173 -176 1249
rect -50 1147 -17 1181
rect 17 1147 50 1181
rect 176 1173 210 1249
rect -210 1105 -176 1139
rect -210 1037 -176 1071
rect -210 969 -176 1003
rect -210 901 -176 935
rect -210 833 -176 867
rect -210 765 -176 799
rect -210 697 -176 731
rect -210 629 -176 663
rect -210 561 -176 595
rect -210 493 -176 527
rect -210 425 -176 459
rect -210 357 -176 391
rect -210 289 -176 323
rect -210 221 -176 255
rect -210 153 -176 187
rect -210 85 -176 119
rect -96 1068 -62 1113
rect -96 1000 -62 1034
rect -96 932 -62 966
rect -96 864 -62 898
rect -96 796 -62 830
rect -96 728 -62 762
rect -96 660 -62 694
rect -96 592 -62 626
rect -96 524 -62 558
rect -96 456 -62 490
rect -96 388 -62 422
rect -96 320 -62 354
rect -96 252 -62 286
rect -96 184 -62 218
rect -96 105 -62 150
rect 62 1068 96 1113
rect 62 1000 96 1034
rect 62 932 96 966
rect 62 864 96 898
rect 62 796 96 830
rect 62 728 96 762
rect 62 660 96 694
rect 62 592 96 626
rect 62 524 96 558
rect 62 456 96 490
rect 62 388 96 422
rect 62 320 96 354
rect 62 252 96 286
rect 62 184 96 218
rect 62 105 96 150
rect 176 1105 210 1139
rect 176 1037 210 1071
rect 176 969 210 1003
rect 176 901 210 935
rect 176 833 210 867
rect 176 765 210 799
rect 176 697 210 731
rect 176 629 210 663
rect 176 561 210 595
rect 176 493 210 527
rect 176 425 210 459
rect 176 357 210 391
rect 176 289 210 323
rect 176 221 210 255
rect 176 153 210 187
rect 176 85 210 119
rect -210 17 -176 51
rect -50 37 -17 71
rect 17 37 50 71
rect -210 -51 -176 -17
rect 176 17 210 51
rect -50 -71 -17 -37
rect 17 -71 50 -37
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -255 -176 -221
rect -210 -323 -176 -289
rect -210 -391 -176 -357
rect -210 -459 -176 -425
rect -210 -527 -176 -493
rect -210 -595 -176 -561
rect -210 -663 -176 -629
rect -210 -731 -176 -697
rect -210 -799 -176 -765
rect -210 -867 -176 -833
rect -210 -935 -176 -901
rect -210 -1003 -176 -969
rect -210 -1071 -176 -1037
rect -210 -1139 -176 -1105
rect -96 -150 -62 -105
rect -96 -218 -62 -184
rect -96 -286 -62 -252
rect -96 -354 -62 -320
rect -96 -422 -62 -388
rect -96 -490 -62 -456
rect -96 -558 -62 -524
rect -96 -626 -62 -592
rect -96 -694 -62 -660
rect -96 -762 -62 -728
rect -96 -830 -62 -796
rect -96 -898 -62 -864
rect -96 -966 -62 -932
rect -96 -1034 -62 -1000
rect -96 -1113 -62 -1068
rect 62 -150 96 -105
rect 62 -218 96 -184
rect 62 -286 96 -252
rect 62 -354 96 -320
rect 62 -422 96 -388
rect 62 -490 96 -456
rect 62 -558 96 -524
rect 62 -626 96 -592
rect 62 -694 96 -660
rect 62 -762 96 -728
rect 62 -830 96 -796
rect 62 -898 96 -864
rect 62 -966 96 -932
rect 62 -1034 96 -1000
rect 62 -1113 96 -1068
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -255 210 -221
rect 176 -323 210 -289
rect 176 -391 210 -357
rect 176 -459 210 -425
rect 176 -527 210 -493
rect 176 -595 210 -561
rect 176 -663 210 -629
rect 176 -731 210 -697
rect 176 -799 210 -765
rect 176 -867 210 -833
rect 176 -935 210 -901
rect 176 -1003 210 -969
rect 176 -1071 210 -1037
rect 176 -1139 210 -1105
rect -210 -1249 -176 -1173
rect -50 -1181 -17 -1147
rect 17 -1181 50 -1147
rect 176 -1249 210 -1173
rect -210 -1283 -85 -1249
rect -51 -1283 -17 -1249
rect 17 -1283 51 -1249
rect 85 -1283 210 -1249
<< properties >>
string FIXED_BBOX -193 -1266 193 1266
<< end >>
