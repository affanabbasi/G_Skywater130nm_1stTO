magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< pwell >>
rect -360 1340 360 1374
rect -360 -1340 -326 1340
rect 326 -1340 360 1340
rect -360 -1374 360 -1340
<< nmoslvt >>
rect -200 -1200 200 1200
<< ndiff >>
rect -258 1173 -200 1200
rect -258 1139 -246 1173
rect -212 1139 -200 1173
rect -258 1105 -200 1139
rect -258 1071 -246 1105
rect -212 1071 -200 1105
rect -258 1037 -200 1071
rect -258 1003 -246 1037
rect -212 1003 -200 1037
rect -258 969 -200 1003
rect -258 935 -246 969
rect -212 935 -200 969
rect -258 901 -200 935
rect -258 867 -246 901
rect -212 867 -200 901
rect -258 833 -200 867
rect -258 799 -246 833
rect -212 799 -200 833
rect -258 765 -200 799
rect -258 731 -246 765
rect -212 731 -200 765
rect -258 697 -200 731
rect -258 663 -246 697
rect -212 663 -200 697
rect -258 629 -200 663
rect -258 595 -246 629
rect -212 595 -200 629
rect -258 561 -200 595
rect -258 527 -246 561
rect -212 527 -200 561
rect -258 493 -200 527
rect -258 459 -246 493
rect -212 459 -200 493
rect -258 425 -200 459
rect -258 391 -246 425
rect -212 391 -200 425
rect -258 357 -200 391
rect -258 323 -246 357
rect -212 323 -200 357
rect -258 289 -200 323
rect -258 255 -246 289
rect -212 255 -200 289
rect -258 221 -200 255
rect -258 187 -246 221
rect -212 187 -200 221
rect -258 153 -200 187
rect -258 119 -246 153
rect -212 119 -200 153
rect -258 85 -200 119
rect -258 51 -246 85
rect -212 51 -200 85
rect -258 17 -200 51
rect -258 -17 -246 17
rect -212 -17 -200 17
rect -258 -51 -200 -17
rect -258 -85 -246 -51
rect -212 -85 -200 -51
rect -258 -119 -200 -85
rect -258 -153 -246 -119
rect -212 -153 -200 -119
rect -258 -187 -200 -153
rect -258 -221 -246 -187
rect -212 -221 -200 -187
rect -258 -255 -200 -221
rect -258 -289 -246 -255
rect -212 -289 -200 -255
rect -258 -323 -200 -289
rect -258 -357 -246 -323
rect -212 -357 -200 -323
rect -258 -391 -200 -357
rect -258 -425 -246 -391
rect -212 -425 -200 -391
rect -258 -459 -200 -425
rect -258 -493 -246 -459
rect -212 -493 -200 -459
rect -258 -527 -200 -493
rect -258 -561 -246 -527
rect -212 -561 -200 -527
rect -258 -595 -200 -561
rect -258 -629 -246 -595
rect -212 -629 -200 -595
rect -258 -663 -200 -629
rect -258 -697 -246 -663
rect -212 -697 -200 -663
rect -258 -731 -200 -697
rect -258 -765 -246 -731
rect -212 -765 -200 -731
rect -258 -799 -200 -765
rect -258 -833 -246 -799
rect -212 -833 -200 -799
rect -258 -867 -200 -833
rect -258 -901 -246 -867
rect -212 -901 -200 -867
rect -258 -935 -200 -901
rect -258 -969 -246 -935
rect -212 -969 -200 -935
rect -258 -1003 -200 -969
rect -258 -1037 -246 -1003
rect -212 -1037 -200 -1003
rect -258 -1071 -200 -1037
rect -258 -1105 -246 -1071
rect -212 -1105 -200 -1071
rect -258 -1139 -200 -1105
rect -258 -1173 -246 -1139
rect -212 -1173 -200 -1139
rect -258 -1200 -200 -1173
rect 200 1173 258 1200
rect 200 1139 212 1173
rect 246 1139 258 1173
rect 200 1105 258 1139
rect 200 1071 212 1105
rect 246 1071 258 1105
rect 200 1037 258 1071
rect 200 1003 212 1037
rect 246 1003 258 1037
rect 200 969 258 1003
rect 200 935 212 969
rect 246 935 258 969
rect 200 901 258 935
rect 200 867 212 901
rect 246 867 258 901
rect 200 833 258 867
rect 200 799 212 833
rect 246 799 258 833
rect 200 765 258 799
rect 200 731 212 765
rect 246 731 258 765
rect 200 697 258 731
rect 200 663 212 697
rect 246 663 258 697
rect 200 629 258 663
rect 200 595 212 629
rect 246 595 258 629
rect 200 561 258 595
rect 200 527 212 561
rect 246 527 258 561
rect 200 493 258 527
rect 200 459 212 493
rect 246 459 258 493
rect 200 425 258 459
rect 200 391 212 425
rect 246 391 258 425
rect 200 357 258 391
rect 200 323 212 357
rect 246 323 258 357
rect 200 289 258 323
rect 200 255 212 289
rect 246 255 258 289
rect 200 221 258 255
rect 200 187 212 221
rect 246 187 258 221
rect 200 153 258 187
rect 200 119 212 153
rect 246 119 258 153
rect 200 85 258 119
rect 200 51 212 85
rect 246 51 258 85
rect 200 17 258 51
rect 200 -17 212 17
rect 246 -17 258 17
rect 200 -51 258 -17
rect 200 -85 212 -51
rect 246 -85 258 -51
rect 200 -119 258 -85
rect 200 -153 212 -119
rect 246 -153 258 -119
rect 200 -187 258 -153
rect 200 -221 212 -187
rect 246 -221 258 -187
rect 200 -255 258 -221
rect 200 -289 212 -255
rect 246 -289 258 -255
rect 200 -323 258 -289
rect 200 -357 212 -323
rect 246 -357 258 -323
rect 200 -391 258 -357
rect 200 -425 212 -391
rect 246 -425 258 -391
rect 200 -459 258 -425
rect 200 -493 212 -459
rect 246 -493 258 -459
rect 200 -527 258 -493
rect 200 -561 212 -527
rect 246 -561 258 -527
rect 200 -595 258 -561
rect 200 -629 212 -595
rect 246 -629 258 -595
rect 200 -663 258 -629
rect 200 -697 212 -663
rect 246 -697 258 -663
rect 200 -731 258 -697
rect 200 -765 212 -731
rect 246 -765 258 -731
rect 200 -799 258 -765
rect 200 -833 212 -799
rect 246 -833 258 -799
rect 200 -867 258 -833
rect 200 -901 212 -867
rect 246 -901 258 -867
rect 200 -935 258 -901
rect 200 -969 212 -935
rect 246 -969 258 -935
rect 200 -1003 258 -969
rect 200 -1037 212 -1003
rect 246 -1037 258 -1003
rect 200 -1071 258 -1037
rect 200 -1105 212 -1071
rect 246 -1105 258 -1071
rect 200 -1139 258 -1105
rect 200 -1173 212 -1139
rect 246 -1173 258 -1139
rect 200 -1200 258 -1173
<< ndiffc >>
rect -246 1139 -212 1173
rect -246 1071 -212 1105
rect -246 1003 -212 1037
rect -246 935 -212 969
rect -246 867 -212 901
rect -246 799 -212 833
rect -246 731 -212 765
rect -246 663 -212 697
rect -246 595 -212 629
rect -246 527 -212 561
rect -246 459 -212 493
rect -246 391 -212 425
rect -246 323 -212 357
rect -246 255 -212 289
rect -246 187 -212 221
rect -246 119 -212 153
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect -246 -153 -212 -119
rect -246 -221 -212 -187
rect -246 -289 -212 -255
rect -246 -357 -212 -323
rect -246 -425 -212 -391
rect -246 -493 -212 -459
rect -246 -561 -212 -527
rect -246 -629 -212 -595
rect -246 -697 -212 -663
rect -246 -765 -212 -731
rect -246 -833 -212 -799
rect -246 -901 -212 -867
rect -246 -969 -212 -935
rect -246 -1037 -212 -1003
rect -246 -1105 -212 -1071
rect -246 -1173 -212 -1139
rect 212 1139 246 1173
rect 212 1071 246 1105
rect 212 1003 246 1037
rect 212 935 246 969
rect 212 867 246 901
rect 212 799 246 833
rect 212 731 246 765
rect 212 663 246 697
rect 212 595 246 629
rect 212 527 246 561
rect 212 459 246 493
rect 212 391 246 425
rect 212 323 246 357
rect 212 255 246 289
rect 212 187 246 221
rect 212 119 246 153
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
rect 212 -153 246 -119
rect 212 -221 246 -187
rect 212 -289 246 -255
rect 212 -357 246 -323
rect 212 -425 246 -391
rect 212 -493 246 -459
rect 212 -561 246 -527
rect 212 -629 246 -595
rect 212 -697 246 -663
rect 212 -765 246 -731
rect 212 -833 246 -799
rect 212 -901 246 -867
rect 212 -969 246 -935
rect 212 -1037 246 -1003
rect 212 -1105 246 -1071
rect 212 -1173 246 -1139
<< psubdiff >>
rect -360 1340 -255 1374
rect -221 1340 -187 1374
rect -153 1340 -119 1374
rect -85 1340 -51 1374
rect -17 1340 17 1374
rect 51 1340 85 1374
rect 119 1340 153 1374
rect 187 1340 221 1374
rect 255 1340 360 1374
rect -360 1275 -326 1340
rect -360 1207 -326 1241
rect 326 1275 360 1340
rect 326 1207 360 1241
rect -360 1139 -326 1173
rect -360 1071 -326 1105
rect -360 1003 -326 1037
rect -360 935 -326 969
rect -360 867 -326 901
rect -360 799 -326 833
rect -360 731 -326 765
rect -360 663 -326 697
rect -360 595 -326 629
rect -360 527 -326 561
rect -360 459 -326 493
rect -360 391 -326 425
rect -360 323 -326 357
rect -360 255 -326 289
rect -360 187 -326 221
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
rect -360 -289 -326 -255
rect -360 -357 -326 -323
rect -360 -425 -326 -391
rect -360 -493 -326 -459
rect -360 -561 -326 -527
rect -360 -629 -326 -595
rect -360 -697 -326 -663
rect -360 -765 -326 -731
rect -360 -833 -326 -799
rect -360 -901 -326 -867
rect -360 -969 -326 -935
rect -360 -1037 -326 -1003
rect -360 -1105 -326 -1071
rect -360 -1173 -326 -1139
rect 326 1139 360 1173
rect 326 1071 360 1105
rect 326 1003 360 1037
rect 326 935 360 969
rect 326 867 360 901
rect 326 799 360 833
rect 326 731 360 765
rect 326 663 360 697
rect 326 595 360 629
rect 326 527 360 561
rect 326 459 360 493
rect 326 391 360 425
rect 326 323 360 357
rect 326 255 360 289
rect 326 187 360 221
rect 326 119 360 153
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect 326 -153 360 -119
rect 326 -221 360 -187
rect 326 -289 360 -255
rect 326 -357 360 -323
rect 326 -425 360 -391
rect 326 -493 360 -459
rect 326 -561 360 -527
rect 326 -629 360 -595
rect 326 -697 360 -663
rect 326 -765 360 -731
rect 326 -833 360 -799
rect 326 -901 360 -867
rect 326 -969 360 -935
rect 326 -1037 360 -1003
rect 326 -1105 360 -1071
rect 326 -1173 360 -1139
rect -360 -1241 -326 -1207
rect -360 -1340 -326 -1275
rect 326 -1241 360 -1207
rect 326 -1340 360 -1275
rect -360 -1374 -255 -1340
rect -221 -1374 -187 -1340
rect -153 -1374 -119 -1340
rect -85 -1374 -51 -1340
rect -17 -1374 17 -1340
rect 51 -1374 85 -1340
rect 119 -1374 153 -1340
rect 187 -1374 221 -1340
rect 255 -1374 360 -1340
<< psubdiffcont >>
rect -255 1340 -221 1374
rect -187 1340 -153 1374
rect -119 1340 -85 1374
rect -51 1340 -17 1374
rect 17 1340 51 1374
rect 85 1340 119 1374
rect 153 1340 187 1374
rect 221 1340 255 1374
rect -360 1241 -326 1275
rect -360 1173 -326 1207
rect 326 1241 360 1275
rect -360 1105 -326 1139
rect -360 1037 -326 1071
rect -360 969 -326 1003
rect -360 901 -326 935
rect -360 833 -326 867
rect -360 765 -326 799
rect -360 697 -326 731
rect -360 629 -326 663
rect -360 561 -326 595
rect -360 493 -326 527
rect -360 425 -326 459
rect -360 357 -326 391
rect -360 289 -326 323
rect -360 221 -326 255
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect -360 -255 -326 -221
rect -360 -323 -326 -289
rect -360 -391 -326 -357
rect -360 -459 -326 -425
rect -360 -527 -326 -493
rect -360 -595 -326 -561
rect -360 -663 -326 -629
rect -360 -731 -326 -697
rect -360 -799 -326 -765
rect -360 -867 -326 -833
rect -360 -935 -326 -901
rect -360 -1003 -326 -969
rect -360 -1071 -326 -1037
rect -360 -1139 -326 -1105
rect -360 -1207 -326 -1173
rect 326 1173 360 1207
rect 326 1105 360 1139
rect 326 1037 360 1071
rect 326 969 360 1003
rect 326 901 360 935
rect 326 833 360 867
rect 326 765 360 799
rect 326 697 360 731
rect 326 629 360 663
rect 326 561 360 595
rect 326 493 360 527
rect 326 425 360 459
rect 326 357 360 391
rect 326 289 360 323
rect 326 221 360 255
rect 326 153 360 187
rect 326 85 360 119
rect 326 17 360 51
rect 326 -51 360 -17
rect 326 -119 360 -85
rect 326 -187 360 -153
rect 326 -255 360 -221
rect 326 -323 360 -289
rect 326 -391 360 -357
rect 326 -459 360 -425
rect 326 -527 360 -493
rect 326 -595 360 -561
rect 326 -663 360 -629
rect 326 -731 360 -697
rect 326 -799 360 -765
rect 326 -867 360 -833
rect 326 -935 360 -901
rect 326 -1003 360 -969
rect 326 -1071 360 -1037
rect 326 -1139 360 -1105
rect -360 -1275 -326 -1241
rect 326 -1207 360 -1173
rect 326 -1275 360 -1241
rect -255 -1374 -221 -1340
rect -187 -1374 -153 -1340
rect -119 -1374 -85 -1340
rect -51 -1374 -17 -1340
rect 17 -1374 51 -1340
rect 85 -1374 119 -1340
rect 153 -1374 187 -1340
rect 221 -1374 255 -1340
<< poly >>
rect -200 1272 200 1288
rect -200 1238 -153 1272
rect -119 1238 -85 1272
rect -51 1238 -17 1272
rect 17 1238 51 1272
rect 85 1238 119 1272
rect 153 1238 200 1272
rect -200 1200 200 1238
rect -200 -1238 200 -1200
rect -200 -1272 -153 -1238
rect -119 -1272 -85 -1238
rect -51 -1272 -17 -1238
rect 17 -1272 51 -1238
rect 85 -1272 119 -1238
rect 153 -1272 200 -1238
rect -200 -1288 200 -1272
<< polycont >>
rect -153 1238 -119 1272
rect -85 1238 -51 1272
rect -17 1238 17 1272
rect 51 1238 85 1272
rect 119 1238 153 1272
rect -153 -1272 -119 -1238
rect -85 -1272 -51 -1238
rect -17 -1272 17 -1238
rect 51 -1272 85 -1238
rect 119 -1272 153 -1238
<< locali >>
rect -360 1340 -255 1374
rect -221 1340 -187 1374
rect -153 1340 -119 1374
rect -85 1340 -51 1374
rect -17 1340 17 1374
rect 51 1340 85 1374
rect 119 1340 153 1374
rect 187 1340 221 1374
rect 255 1340 360 1374
rect -360 1275 -326 1340
rect 326 1275 360 1340
rect -360 1207 -326 1241
rect -200 1238 -153 1272
rect -119 1238 -85 1272
rect -51 1238 -17 1272
rect 17 1238 51 1272
rect 85 1238 119 1272
rect 153 1238 200 1272
rect 326 1207 360 1241
rect -360 1139 -326 1173
rect -360 1071 -326 1105
rect -360 1003 -326 1037
rect -360 935 -326 969
rect -360 867 -326 901
rect -360 799 -326 833
rect -360 731 -326 765
rect -360 663 -326 697
rect -360 595 -326 629
rect -360 527 -326 561
rect -360 459 -326 493
rect -360 391 -326 425
rect -360 323 -326 357
rect -360 255 -326 289
rect -360 187 -326 221
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
rect -360 -289 -326 -255
rect -360 -357 -326 -323
rect -360 -425 -326 -391
rect -360 -493 -326 -459
rect -360 -561 -326 -527
rect -360 -629 -326 -595
rect -360 -697 -326 -663
rect -360 -765 -326 -731
rect -360 -833 -326 -799
rect -360 -901 -326 -867
rect -360 -969 -326 -935
rect -360 -1037 -326 -1003
rect -360 -1105 -326 -1071
rect -360 -1173 -326 -1139
rect -246 1173 -212 1204
rect -246 1105 -212 1139
rect -246 1037 -212 1071
rect -246 969 -212 1003
rect -246 901 -212 935
rect -246 833 -212 867
rect -246 765 -212 799
rect -246 697 -212 731
rect -246 629 -212 663
rect -246 561 -212 595
rect -246 493 -212 527
rect -246 425 -212 459
rect -246 357 -212 391
rect -246 289 -212 323
rect -246 221 -212 255
rect -246 153 -212 187
rect -246 85 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -85
rect -246 -187 -212 -153
rect -246 -255 -212 -221
rect -246 -323 -212 -289
rect -246 -391 -212 -357
rect -246 -459 -212 -425
rect -246 -527 -212 -493
rect -246 -595 -212 -561
rect -246 -663 -212 -629
rect -246 -731 -212 -697
rect -246 -799 -212 -765
rect -246 -867 -212 -833
rect -246 -935 -212 -901
rect -246 -1003 -212 -969
rect -246 -1071 -212 -1037
rect -246 -1139 -212 -1105
rect -246 -1204 -212 -1173
rect 212 1173 246 1204
rect 212 1105 246 1139
rect 212 1037 246 1071
rect 212 969 246 1003
rect 212 901 246 935
rect 212 833 246 867
rect 212 765 246 799
rect 212 697 246 731
rect 212 629 246 663
rect 212 561 246 595
rect 212 493 246 527
rect 212 425 246 459
rect 212 357 246 391
rect 212 289 246 323
rect 212 221 246 255
rect 212 153 246 187
rect 212 85 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -85
rect 212 -187 246 -153
rect 212 -255 246 -221
rect 212 -323 246 -289
rect 212 -391 246 -357
rect 212 -459 246 -425
rect 212 -527 246 -493
rect 212 -595 246 -561
rect 212 -663 246 -629
rect 212 -731 246 -697
rect 212 -799 246 -765
rect 212 -867 246 -833
rect 212 -935 246 -901
rect 212 -1003 246 -969
rect 212 -1071 246 -1037
rect 212 -1139 246 -1105
rect 212 -1204 246 -1173
rect 326 1139 360 1173
rect 326 1071 360 1105
rect 326 1003 360 1037
rect 326 935 360 969
rect 326 867 360 901
rect 326 799 360 833
rect 326 731 360 765
rect 326 663 360 697
rect 326 595 360 629
rect 326 527 360 561
rect 326 459 360 493
rect 326 391 360 425
rect 326 323 360 357
rect 326 255 360 289
rect 326 187 360 221
rect 326 119 360 153
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect 326 -153 360 -119
rect 326 -221 360 -187
rect 326 -289 360 -255
rect 326 -357 360 -323
rect 326 -425 360 -391
rect 326 -493 360 -459
rect 326 -561 360 -527
rect 326 -629 360 -595
rect 326 -697 360 -663
rect 326 -765 360 -731
rect 326 -833 360 -799
rect 326 -901 360 -867
rect 326 -969 360 -935
rect 326 -1037 360 -1003
rect 326 -1105 360 -1071
rect 326 -1173 360 -1139
rect -360 -1241 -326 -1207
rect -200 -1272 -153 -1238
rect -119 -1272 -85 -1238
rect -51 -1272 -17 -1238
rect 17 -1272 51 -1238
rect 85 -1272 119 -1238
rect 153 -1272 200 -1238
rect 326 -1241 360 -1207
rect -360 -1340 -326 -1275
rect 326 -1340 360 -1275
rect -360 -1374 -255 -1340
rect -221 -1374 -187 -1340
rect -153 -1374 -119 -1340
rect -85 -1374 -51 -1340
rect -17 -1374 17 -1340
rect 51 -1374 85 -1340
rect 119 -1374 153 -1340
rect 187 -1374 221 -1340
rect 255 -1374 360 -1340
<< properties >>
string FIXED_BBOX -342 -1356 342 1356
<< end >>
