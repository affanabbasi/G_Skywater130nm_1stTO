magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< error_p >>
rect -31 181 31 187
rect -31 147 -17 181
rect -31 141 31 147
rect -31 -147 31 -141
rect -31 -181 -17 -147
rect -31 -187 31 -181
<< nwell >>
rect -231 -319 231 319
<< pmoslvt >>
rect -35 -100 35 100
<< pdiff >>
rect -93 85 -35 100
rect -93 51 -81 85
rect -47 51 -35 85
rect -93 17 -35 51
rect -93 -17 -81 17
rect -47 -17 -35 17
rect -93 -51 -35 -17
rect -93 -85 -81 -51
rect -47 -85 -35 -51
rect -93 -100 -35 -85
rect 35 85 93 100
rect 35 51 47 85
rect 81 51 93 85
rect 35 17 93 51
rect 35 -17 47 17
rect 81 -17 93 17
rect 35 -51 93 -17
rect 35 -85 47 -51
rect 81 -85 93 -51
rect 35 -100 93 -85
<< pdiffc >>
rect -81 51 -47 85
rect -81 -17 -47 17
rect -81 -85 -47 -51
rect 47 51 81 85
rect 47 -17 81 17
rect 47 -85 81 -51
<< nsubdiff >>
rect -195 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 195 283
rect -195 187 -161 249
rect -195 119 -161 153
rect 161 187 195 249
rect 161 119 195 153
rect -195 51 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -51
rect 161 51 195 85
rect 161 -17 195 17
rect 161 -85 195 -51
rect -195 -153 -161 -119
rect -195 -249 -161 -187
rect 161 -153 195 -119
rect 161 -249 195 -187
rect -195 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 195 -249
<< nsubdiffcont >>
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect -195 153 -161 187
rect -195 85 -161 119
rect 161 153 195 187
rect -195 17 -161 51
rect -195 -51 -161 -17
rect -195 -119 -161 -85
rect 161 85 195 119
rect 161 17 195 51
rect 161 -51 195 -17
rect -195 -187 -161 -153
rect 161 -119 195 -85
rect 161 -187 195 -153
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
<< poly >>
rect -35 181 35 197
rect -35 147 -17 181
rect 17 147 35 181
rect -35 100 35 147
rect -35 -147 35 -100
rect -35 -181 -17 -147
rect 17 -181 35 -147
rect -35 -197 35 -181
<< polycont >>
rect -17 147 17 181
rect -17 -181 17 -147
<< locali >>
rect -195 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 195 283
rect -195 187 -161 249
rect 161 187 195 249
rect -195 119 -161 153
rect -35 147 -17 181
rect 17 147 35 181
rect 161 119 195 153
rect -195 51 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -51
rect -81 85 -47 104
rect -81 17 -47 19
rect -81 -19 -47 -17
rect -81 -104 -47 -85
rect 47 85 81 104
rect 47 17 81 19
rect 47 -19 81 -17
rect 47 -104 81 -85
rect 161 51 195 85
rect 161 -17 195 17
rect 161 -85 195 -51
rect -195 -153 -161 -119
rect -35 -181 -17 -147
rect 17 -181 35 -147
rect 161 -153 195 -119
rect -195 -249 -161 -187
rect 161 -249 195 -187
rect -195 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 195 -249
<< viali >>
rect -17 147 17 181
rect -81 51 -47 53
rect -81 19 -47 51
rect -81 -51 -47 -19
rect -81 -53 -47 -51
rect 47 51 81 53
rect 47 19 81 51
rect 47 -51 81 -19
rect 47 -53 81 -51
rect -17 -181 17 -147
<< metal1 >>
rect -31 181 31 187
rect -31 147 -17 181
rect 17 147 31 181
rect -31 141 31 147
rect -87 53 -41 100
rect -87 19 -81 53
rect -47 19 -41 53
rect -87 -19 -41 19
rect -87 -53 -81 -19
rect -47 -53 -41 -19
rect -87 -100 -41 -53
rect 41 53 87 100
rect 41 19 47 53
rect 81 19 87 53
rect 41 -19 87 19
rect 41 -53 47 -19
rect 81 -53 87 -19
rect 41 -100 87 -53
rect -31 -147 31 -141
rect -31 -181 -17 -147
rect 17 -181 31 -147
rect -31 -187 31 -181
<< properties >>
string FIXED_BBOX -178 -266 178 266
<< end >>
