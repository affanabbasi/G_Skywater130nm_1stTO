magic
tech sky130A
magscale 1 2
timestamp 1611881054
<< nwell >>
rect -1312 -1019 1312 1019
<< pmoslvt >>
rect -1116 -800 -716 800
rect -658 -800 -258 800
rect -200 -800 200 800
rect 258 -800 658 800
rect 716 -800 1116 800
<< pdiff >>
rect -1174 765 -1116 800
rect -1174 731 -1162 765
rect -1128 731 -1116 765
rect -1174 697 -1116 731
rect -1174 663 -1162 697
rect -1128 663 -1116 697
rect -1174 629 -1116 663
rect -1174 595 -1162 629
rect -1128 595 -1116 629
rect -1174 561 -1116 595
rect -1174 527 -1162 561
rect -1128 527 -1116 561
rect -1174 493 -1116 527
rect -1174 459 -1162 493
rect -1128 459 -1116 493
rect -1174 425 -1116 459
rect -1174 391 -1162 425
rect -1128 391 -1116 425
rect -1174 357 -1116 391
rect -1174 323 -1162 357
rect -1128 323 -1116 357
rect -1174 289 -1116 323
rect -1174 255 -1162 289
rect -1128 255 -1116 289
rect -1174 221 -1116 255
rect -1174 187 -1162 221
rect -1128 187 -1116 221
rect -1174 153 -1116 187
rect -1174 119 -1162 153
rect -1128 119 -1116 153
rect -1174 85 -1116 119
rect -1174 51 -1162 85
rect -1128 51 -1116 85
rect -1174 17 -1116 51
rect -1174 -17 -1162 17
rect -1128 -17 -1116 17
rect -1174 -51 -1116 -17
rect -1174 -85 -1162 -51
rect -1128 -85 -1116 -51
rect -1174 -119 -1116 -85
rect -1174 -153 -1162 -119
rect -1128 -153 -1116 -119
rect -1174 -187 -1116 -153
rect -1174 -221 -1162 -187
rect -1128 -221 -1116 -187
rect -1174 -255 -1116 -221
rect -1174 -289 -1162 -255
rect -1128 -289 -1116 -255
rect -1174 -323 -1116 -289
rect -1174 -357 -1162 -323
rect -1128 -357 -1116 -323
rect -1174 -391 -1116 -357
rect -1174 -425 -1162 -391
rect -1128 -425 -1116 -391
rect -1174 -459 -1116 -425
rect -1174 -493 -1162 -459
rect -1128 -493 -1116 -459
rect -1174 -527 -1116 -493
rect -1174 -561 -1162 -527
rect -1128 -561 -1116 -527
rect -1174 -595 -1116 -561
rect -1174 -629 -1162 -595
rect -1128 -629 -1116 -595
rect -1174 -663 -1116 -629
rect -1174 -697 -1162 -663
rect -1128 -697 -1116 -663
rect -1174 -731 -1116 -697
rect -1174 -765 -1162 -731
rect -1128 -765 -1116 -731
rect -1174 -800 -1116 -765
rect -716 765 -658 800
rect -716 731 -704 765
rect -670 731 -658 765
rect -716 697 -658 731
rect -716 663 -704 697
rect -670 663 -658 697
rect -716 629 -658 663
rect -716 595 -704 629
rect -670 595 -658 629
rect -716 561 -658 595
rect -716 527 -704 561
rect -670 527 -658 561
rect -716 493 -658 527
rect -716 459 -704 493
rect -670 459 -658 493
rect -716 425 -658 459
rect -716 391 -704 425
rect -670 391 -658 425
rect -716 357 -658 391
rect -716 323 -704 357
rect -670 323 -658 357
rect -716 289 -658 323
rect -716 255 -704 289
rect -670 255 -658 289
rect -716 221 -658 255
rect -716 187 -704 221
rect -670 187 -658 221
rect -716 153 -658 187
rect -716 119 -704 153
rect -670 119 -658 153
rect -716 85 -658 119
rect -716 51 -704 85
rect -670 51 -658 85
rect -716 17 -658 51
rect -716 -17 -704 17
rect -670 -17 -658 17
rect -716 -51 -658 -17
rect -716 -85 -704 -51
rect -670 -85 -658 -51
rect -716 -119 -658 -85
rect -716 -153 -704 -119
rect -670 -153 -658 -119
rect -716 -187 -658 -153
rect -716 -221 -704 -187
rect -670 -221 -658 -187
rect -716 -255 -658 -221
rect -716 -289 -704 -255
rect -670 -289 -658 -255
rect -716 -323 -658 -289
rect -716 -357 -704 -323
rect -670 -357 -658 -323
rect -716 -391 -658 -357
rect -716 -425 -704 -391
rect -670 -425 -658 -391
rect -716 -459 -658 -425
rect -716 -493 -704 -459
rect -670 -493 -658 -459
rect -716 -527 -658 -493
rect -716 -561 -704 -527
rect -670 -561 -658 -527
rect -716 -595 -658 -561
rect -716 -629 -704 -595
rect -670 -629 -658 -595
rect -716 -663 -658 -629
rect -716 -697 -704 -663
rect -670 -697 -658 -663
rect -716 -731 -658 -697
rect -716 -765 -704 -731
rect -670 -765 -658 -731
rect -716 -800 -658 -765
rect -258 765 -200 800
rect -258 731 -246 765
rect -212 731 -200 765
rect -258 697 -200 731
rect -258 663 -246 697
rect -212 663 -200 697
rect -258 629 -200 663
rect -258 595 -246 629
rect -212 595 -200 629
rect -258 561 -200 595
rect -258 527 -246 561
rect -212 527 -200 561
rect -258 493 -200 527
rect -258 459 -246 493
rect -212 459 -200 493
rect -258 425 -200 459
rect -258 391 -246 425
rect -212 391 -200 425
rect -258 357 -200 391
rect -258 323 -246 357
rect -212 323 -200 357
rect -258 289 -200 323
rect -258 255 -246 289
rect -212 255 -200 289
rect -258 221 -200 255
rect -258 187 -246 221
rect -212 187 -200 221
rect -258 153 -200 187
rect -258 119 -246 153
rect -212 119 -200 153
rect -258 85 -200 119
rect -258 51 -246 85
rect -212 51 -200 85
rect -258 17 -200 51
rect -258 -17 -246 17
rect -212 -17 -200 17
rect -258 -51 -200 -17
rect -258 -85 -246 -51
rect -212 -85 -200 -51
rect -258 -119 -200 -85
rect -258 -153 -246 -119
rect -212 -153 -200 -119
rect -258 -187 -200 -153
rect -258 -221 -246 -187
rect -212 -221 -200 -187
rect -258 -255 -200 -221
rect -258 -289 -246 -255
rect -212 -289 -200 -255
rect -258 -323 -200 -289
rect -258 -357 -246 -323
rect -212 -357 -200 -323
rect -258 -391 -200 -357
rect -258 -425 -246 -391
rect -212 -425 -200 -391
rect -258 -459 -200 -425
rect -258 -493 -246 -459
rect -212 -493 -200 -459
rect -258 -527 -200 -493
rect -258 -561 -246 -527
rect -212 -561 -200 -527
rect -258 -595 -200 -561
rect -258 -629 -246 -595
rect -212 -629 -200 -595
rect -258 -663 -200 -629
rect -258 -697 -246 -663
rect -212 -697 -200 -663
rect -258 -731 -200 -697
rect -258 -765 -246 -731
rect -212 -765 -200 -731
rect -258 -800 -200 -765
rect 200 765 258 800
rect 200 731 212 765
rect 246 731 258 765
rect 200 697 258 731
rect 200 663 212 697
rect 246 663 258 697
rect 200 629 258 663
rect 200 595 212 629
rect 246 595 258 629
rect 200 561 258 595
rect 200 527 212 561
rect 246 527 258 561
rect 200 493 258 527
rect 200 459 212 493
rect 246 459 258 493
rect 200 425 258 459
rect 200 391 212 425
rect 246 391 258 425
rect 200 357 258 391
rect 200 323 212 357
rect 246 323 258 357
rect 200 289 258 323
rect 200 255 212 289
rect 246 255 258 289
rect 200 221 258 255
rect 200 187 212 221
rect 246 187 258 221
rect 200 153 258 187
rect 200 119 212 153
rect 246 119 258 153
rect 200 85 258 119
rect 200 51 212 85
rect 246 51 258 85
rect 200 17 258 51
rect 200 -17 212 17
rect 246 -17 258 17
rect 200 -51 258 -17
rect 200 -85 212 -51
rect 246 -85 258 -51
rect 200 -119 258 -85
rect 200 -153 212 -119
rect 246 -153 258 -119
rect 200 -187 258 -153
rect 200 -221 212 -187
rect 246 -221 258 -187
rect 200 -255 258 -221
rect 200 -289 212 -255
rect 246 -289 258 -255
rect 200 -323 258 -289
rect 200 -357 212 -323
rect 246 -357 258 -323
rect 200 -391 258 -357
rect 200 -425 212 -391
rect 246 -425 258 -391
rect 200 -459 258 -425
rect 200 -493 212 -459
rect 246 -493 258 -459
rect 200 -527 258 -493
rect 200 -561 212 -527
rect 246 -561 258 -527
rect 200 -595 258 -561
rect 200 -629 212 -595
rect 246 -629 258 -595
rect 200 -663 258 -629
rect 200 -697 212 -663
rect 246 -697 258 -663
rect 200 -731 258 -697
rect 200 -765 212 -731
rect 246 -765 258 -731
rect 200 -800 258 -765
rect 658 765 716 800
rect 658 731 670 765
rect 704 731 716 765
rect 658 697 716 731
rect 658 663 670 697
rect 704 663 716 697
rect 658 629 716 663
rect 658 595 670 629
rect 704 595 716 629
rect 658 561 716 595
rect 658 527 670 561
rect 704 527 716 561
rect 658 493 716 527
rect 658 459 670 493
rect 704 459 716 493
rect 658 425 716 459
rect 658 391 670 425
rect 704 391 716 425
rect 658 357 716 391
rect 658 323 670 357
rect 704 323 716 357
rect 658 289 716 323
rect 658 255 670 289
rect 704 255 716 289
rect 658 221 716 255
rect 658 187 670 221
rect 704 187 716 221
rect 658 153 716 187
rect 658 119 670 153
rect 704 119 716 153
rect 658 85 716 119
rect 658 51 670 85
rect 704 51 716 85
rect 658 17 716 51
rect 658 -17 670 17
rect 704 -17 716 17
rect 658 -51 716 -17
rect 658 -85 670 -51
rect 704 -85 716 -51
rect 658 -119 716 -85
rect 658 -153 670 -119
rect 704 -153 716 -119
rect 658 -187 716 -153
rect 658 -221 670 -187
rect 704 -221 716 -187
rect 658 -255 716 -221
rect 658 -289 670 -255
rect 704 -289 716 -255
rect 658 -323 716 -289
rect 658 -357 670 -323
rect 704 -357 716 -323
rect 658 -391 716 -357
rect 658 -425 670 -391
rect 704 -425 716 -391
rect 658 -459 716 -425
rect 658 -493 670 -459
rect 704 -493 716 -459
rect 658 -527 716 -493
rect 658 -561 670 -527
rect 704 -561 716 -527
rect 658 -595 716 -561
rect 658 -629 670 -595
rect 704 -629 716 -595
rect 658 -663 716 -629
rect 658 -697 670 -663
rect 704 -697 716 -663
rect 658 -731 716 -697
rect 658 -765 670 -731
rect 704 -765 716 -731
rect 658 -800 716 -765
rect 1116 765 1174 800
rect 1116 731 1128 765
rect 1162 731 1174 765
rect 1116 697 1174 731
rect 1116 663 1128 697
rect 1162 663 1174 697
rect 1116 629 1174 663
rect 1116 595 1128 629
rect 1162 595 1174 629
rect 1116 561 1174 595
rect 1116 527 1128 561
rect 1162 527 1174 561
rect 1116 493 1174 527
rect 1116 459 1128 493
rect 1162 459 1174 493
rect 1116 425 1174 459
rect 1116 391 1128 425
rect 1162 391 1174 425
rect 1116 357 1174 391
rect 1116 323 1128 357
rect 1162 323 1174 357
rect 1116 289 1174 323
rect 1116 255 1128 289
rect 1162 255 1174 289
rect 1116 221 1174 255
rect 1116 187 1128 221
rect 1162 187 1174 221
rect 1116 153 1174 187
rect 1116 119 1128 153
rect 1162 119 1174 153
rect 1116 85 1174 119
rect 1116 51 1128 85
rect 1162 51 1174 85
rect 1116 17 1174 51
rect 1116 -17 1128 17
rect 1162 -17 1174 17
rect 1116 -51 1174 -17
rect 1116 -85 1128 -51
rect 1162 -85 1174 -51
rect 1116 -119 1174 -85
rect 1116 -153 1128 -119
rect 1162 -153 1174 -119
rect 1116 -187 1174 -153
rect 1116 -221 1128 -187
rect 1162 -221 1174 -187
rect 1116 -255 1174 -221
rect 1116 -289 1128 -255
rect 1162 -289 1174 -255
rect 1116 -323 1174 -289
rect 1116 -357 1128 -323
rect 1162 -357 1174 -323
rect 1116 -391 1174 -357
rect 1116 -425 1128 -391
rect 1162 -425 1174 -391
rect 1116 -459 1174 -425
rect 1116 -493 1128 -459
rect 1162 -493 1174 -459
rect 1116 -527 1174 -493
rect 1116 -561 1128 -527
rect 1162 -561 1174 -527
rect 1116 -595 1174 -561
rect 1116 -629 1128 -595
rect 1162 -629 1174 -595
rect 1116 -663 1174 -629
rect 1116 -697 1128 -663
rect 1162 -697 1174 -663
rect 1116 -731 1174 -697
rect 1116 -765 1128 -731
rect 1162 -765 1174 -731
rect 1116 -800 1174 -765
<< pdiffc >>
rect -1162 731 -1128 765
rect -1162 663 -1128 697
rect -1162 595 -1128 629
rect -1162 527 -1128 561
rect -1162 459 -1128 493
rect -1162 391 -1128 425
rect -1162 323 -1128 357
rect -1162 255 -1128 289
rect -1162 187 -1128 221
rect -1162 119 -1128 153
rect -1162 51 -1128 85
rect -1162 -17 -1128 17
rect -1162 -85 -1128 -51
rect -1162 -153 -1128 -119
rect -1162 -221 -1128 -187
rect -1162 -289 -1128 -255
rect -1162 -357 -1128 -323
rect -1162 -425 -1128 -391
rect -1162 -493 -1128 -459
rect -1162 -561 -1128 -527
rect -1162 -629 -1128 -595
rect -1162 -697 -1128 -663
rect -1162 -765 -1128 -731
rect -704 731 -670 765
rect -704 663 -670 697
rect -704 595 -670 629
rect -704 527 -670 561
rect -704 459 -670 493
rect -704 391 -670 425
rect -704 323 -670 357
rect -704 255 -670 289
rect -704 187 -670 221
rect -704 119 -670 153
rect -704 51 -670 85
rect -704 -17 -670 17
rect -704 -85 -670 -51
rect -704 -153 -670 -119
rect -704 -221 -670 -187
rect -704 -289 -670 -255
rect -704 -357 -670 -323
rect -704 -425 -670 -391
rect -704 -493 -670 -459
rect -704 -561 -670 -527
rect -704 -629 -670 -595
rect -704 -697 -670 -663
rect -704 -765 -670 -731
rect -246 731 -212 765
rect -246 663 -212 697
rect -246 595 -212 629
rect -246 527 -212 561
rect -246 459 -212 493
rect -246 391 -212 425
rect -246 323 -212 357
rect -246 255 -212 289
rect -246 187 -212 221
rect -246 119 -212 153
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect -246 -153 -212 -119
rect -246 -221 -212 -187
rect -246 -289 -212 -255
rect -246 -357 -212 -323
rect -246 -425 -212 -391
rect -246 -493 -212 -459
rect -246 -561 -212 -527
rect -246 -629 -212 -595
rect -246 -697 -212 -663
rect -246 -765 -212 -731
rect 212 731 246 765
rect 212 663 246 697
rect 212 595 246 629
rect 212 527 246 561
rect 212 459 246 493
rect 212 391 246 425
rect 212 323 246 357
rect 212 255 246 289
rect 212 187 246 221
rect 212 119 246 153
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
rect 212 -153 246 -119
rect 212 -221 246 -187
rect 212 -289 246 -255
rect 212 -357 246 -323
rect 212 -425 246 -391
rect 212 -493 246 -459
rect 212 -561 246 -527
rect 212 -629 246 -595
rect 212 -697 246 -663
rect 212 -765 246 -731
rect 670 731 704 765
rect 670 663 704 697
rect 670 595 704 629
rect 670 527 704 561
rect 670 459 704 493
rect 670 391 704 425
rect 670 323 704 357
rect 670 255 704 289
rect 670 187 704 221
rect 670 119 704 153
rect 670 51 704 85
rect 670 -17 704 17
rect 670 -85 704 -51
rect 670 -153 704 -119
rect 670 -221 704 -187
rect 670 -289 704 -255
rect 670 -357 704 -323
rect 670 -425 704 -391
rect 670 -493 704 -459
rect 670 -561 704 -527
rect 670 -629 704 -595
rect 670 -697 704 -663
rect 670 -765 704 -731
rect 1128 731 1162 765
rect 1128 663 1162 697
rect 1128 595 1162 629
rect 1128 527 1162 561
rect 1128 459 1162 493
rect 1128 391 1162 425
rect 1128 323 1162 357
rect 1128 255 1162 289
rect 1128 187 1162 221
rect 1128 119 1162 153
rect 1128 51 1162 85
rect 1128 -17 1162 17
rect 1128 -85 1162 -51
rect 1128 -153 1162 -119
rect 1128 -221 1162 -187
rect 1128 -289 1162 -255
rect 1128 -357 1162 -323
rect 1128 -425 1162 -391
rect 1128 -493 1162 -459
rect 1128 -561 1162 -527
rect 1128 -629 1162 -595
rect 1128 -697 1162 -663
rect 1128 -765 1162 -731
<< nsubdiff >>
rect -1276 949 -1173 983
rect -1139 949 -1105 983
rect -1071 949 -1037 983
rect -1003 949 -969 983
rect -935 949 -901 983
rect -867 949 -833 983
rect -799 949 -765 983
rect -731 949 -697 983
rect -663 949 -629 983
rect -595 949 -561 983
rect -527 949 -493 983
rect -459 949 -425 983
rect -391 949 -357 983
rect -323 949 -289 983
rect -255 949 -221 983
rect -187 949 -153 983
rect -119 949 -85 983
rect -51 949 -17 983
rect 17 949 51 983
rect 85 949 119 983
rect 153 949 187 983
rect 221 949 255 983
rect 289 949 323 983
rect 357 949 391 983
rect 425 949 459 983
rect 493 949 527 983
rect 561 949 595 983
rect 629 949 663 983
rect 697 949 731 983
rect 765 949 799 983
rect 833 949 867 983
rect 901 949 935 983
rect 969 949 1003 983
rect 1037 949 1071 983
rect 1105 949 1139 983
rect 1173 949 1276 983
rect -1276 867 -1242 949
rect -1276 799 -1242 833
rect 1242 867 1276 949
rect -1276 731 -1242 765
rect -1276 663 -1242 697
rect -1276 595 -1242 629
rect -1276 527 -1242 561
rect -1276 459 -1242 493
rect -1276 391 -1242 425
rect -1276 323 -1242 357
rect -1276 255 -1242 289
rect -1276 187 -1242 221
rect -1276 119 -1242 153
rect -1276 51 -1242 85
rect -1276 -17 -1242 17
rect -1276 -85 -1242 -51
rect -1276 -153 -1242 -119
rect -1276 -221 -1242 -187
rect -1276 -289 -1242 -255
rect -1276 -357 -1242 -323
rect -1276 -425 -1242 -391
rect -1276 -493 -1242 -459
rect -1276 -561 -1242 -527
rect -1276 -629 -1242 -595
rect -1276 -697 -1242 -663
rect -1276 -765 -1242 -731
rect -1276 -833 -1242 -799
rect 1242 799 1276 833
rect 1242 731 1276 765
rect 1242 663 1276 697
rect 1242 595 1276 629
rect 1242 527 1276 561
rect 1242 459 1276 493
rect 1242 391 1276 425
rect 1242 323 1276 357
rect 1242 255 1276 289
rect 1242 187 1276 221
rect 1242 119 1276 153
rect 1242 51 1276 85
rect 1242 -17 1276 17
rect 1242 -85 1276 -51
rect 1242 -153 1276 -119
rect 1242 -221 1276 -187
rect 1242 -289 1276 -255
rect 1242 -357 1276 -323
rect 1242 -425 1276 -391
rect 1242 -493 1276 -459
rect 1242 -561 1276 -527
rect 1242 -629 1276 -595
rect 1242 -697 1276 -663
rect 1242 -765 1276 -731
rect -1276 -949 -1242 -867
rect 1242 -833 1276 -799
rect 1242 -949 1276 -867
rect -1276 -983 -1173 -949
rect -1139 -983 -1105 -949
rect -1071 -983 -1037 -949
rect -1003 -983 -969 -949
rect -935 -983 -901 -949
rect -867 -983 -833 -949
rect -799 -983 -765 -949
rect -731 -983 -697 -949
rect -663 -983 -629 -949
rect -595 -983 -561 -949
rect -527 -983 -493 -949
rect -459 -983 -425 -949
rect -391 -983 -357 -949
rect -323 -983 -289 -949
rect -255 -983 -221 -949
rect -187 -983 -153 -949
rect -119 -983 -85 -949
rect -51 -983 -17 -949
rect 17 -983 51 -949
rect 85 -983 119 -949
rect 153 -983 187 -949
rect 221 -983 255 -949
rect 289 -983 323 -949
rect 357 -983 391 -949
rect 425 -983 459 -949
rect 493 -983 527 -949
rect 561 -983 595 -949
rect 629 -983 663 -949
rect 697 -983 731 -949
rect 765 -983 799 -949
rect 833 -983 867 -949
rect 901 -983 935 -949
rect 969 -983 1003 -949
rect 1037 -983 1071 -949
rect 1105 -983 1139 -949
rect 1173 -983 1276 -949
<< nsubdiffcont >>
rect -1173 949 -1139 983
rect -1105 949 -1071 983
rect -1037 949 -1003 983
rect -969 949 -935 983
rect -901 949 -867 983
rect -833 949 -799 983
rect -765 949 -731 983
rect -697 949 -663 983
rect -629 949 -595 983
rect -561 949 -527 983
rect -493 949 -459 983
rect -425 949 -391 983
rect -357 949 -323 983
rect -289 949 -255 983
rect -221 949 -187 983
rect -153 949 -119 983
rect -85 949 -51 983
rect -17 949 17 983
rect 51 949 85 983
rect 119 949 153 983
rect 187 949 221 983
rect 255 949 289 983
rect 323 949 357 983
rect 391 949 425 983
rect 459 949 493 983
rect 527 949 561 983
rect 595 949 629 983
rect 663 949 697 983
rect 731 949 765 983
rect 799 949 833 983
rect 867 949 901 983
rect 935 949 969 983
rect 1003 949 1037 983
rect 1071 949 1105 983
rect 1139 949 1173 983
rect -1276 833 -1242 867
rect 1242 833 1276 867
rect -1276 765 -1242 799
rect -1276 697 -1242 731
rect -1276 629 -1242 663
rect -1276 561 -1242 595
rect -1276 493 -1242 527
rect -1276 425 -1242 459
rect -1276 357 -1242 391
rect -1276 289 -1242 323
rect -1276 221 -1242 255
rect -1276 153 -1242 187
rect -1276 85 -1242 119
rect -1276 17 -1242 51
rect -1276 -51 -1242 -17
rect -1276 -119 -1242 -85
rect -1276 -187 -1242 -153
rect -1276 -255 -1242 -221
rect -1276 -323 -1242 -289
rect -1276 -391 -1242 -357
rect -1276 -459 -1242 -425
rect -1276 -527 -1242 -493
rect -1276 -595 -1242 -561
rect -1276 -663 -1242 -629
rect -1276 -731 -1242 -697
rect -1276 -799 -1242 -765
rect 1242 765 1276 799
rect 1242 697 1276 731
rect 1242 629 1276 663
rect 1242 561 1276 595
rect 1242 493 1276 527
rect 1242 425 1276 459
rect 1242 357 1276 391
rect 1242 289 1276 323
rect 1242 221 1276 255
rect 1242 153 1276 187
rect 1242 85 1276 119
rect 1242 17 1276 51
rect 1242 -51 1276 -17
rect 1242 -119 1276 -85
rect 1242 -187 1276 -153
rect 1242 -255 1276 -221
rect 1242 -323 1276 -289
rect 1242 -391 1276 -357
rect 1242 -459 1276 -425
rect 1242 -527 1276 -493
rect 1242 -595 1276 -561
rect 1242 -663 1276 -629
rect 1242 -731 1276 -697
rect 1242 -799 1276 -765
rect -1276 -867 -1242 -833
rect 1242 -867 1276 -833
rect -1173 -983 -1139 -949
rect -1105 -983 -1071 -949
rect -1037 -983 -1003 -949
rect -969 -983 -935 -949
rect -901 -983 -867 -949
rect -833 -983 -799 -949
rect -765 -983 -731 -949
rect -697 -983 -663 -949
rect -629 -983 -595 -949
rect -561 -983 -527 -949
rect -493 -983 -459 -949
rect -425 -983 -391 -949
rect -357 -983 -323 -949
rect -289 -983 -255 -949
rect -221 -983 -187 -949
rect -153 -983 -119 -949
rect -85 -983 -51 -949
rect -17 -983 17 -949
rect 51 -983 85 -949
rect 119 -983 153 -949
rect 187 -983 221 -949
rect 255 -983 289 -949
rect 323 -983 357 -949
rect 391 -983 425 -949
rect 459 -983 493 -949
rect 527 -983 561 -949
rect 595 -983 629 -949
rect 663 -983 697 -949
rect 731 -983 765 -949
rect 799 -983 833 -949
rect 867 -983 901 -949
rect 935 -983 969 -949
rect 1003 -983 1037 -949
rect 1071 -983 1105 -949
rect 1139 -983 1173 -949
<< poly >>
rect -969 881 -863 897
rect -969 864 -933 881
rect -1116 847 -933 864
rect -899 864 -863 881
rect -511 881 -405 897
rect -511 864 -475 881
rect -899 847 -716 864
rect -1116 800 -716 847
rect -658 847 -475 864
rect -441 864 -405 881
rect -53 881 53 897
rect -53 864 -17 881
rect -441 847 -258 864
rect -658 800 -258 847
rect -200 847 -17 864
rect 17 864 53 881
rect 405 881 511 897
rect 405 864 441 881
rect 17 847 200 864
rect -200 800 200 847
rect 258 847 441 864
rect 475 864 511 881
rect 863 881 969 897
rect 863 864 899 881
rect 475 847 658 864
rect 258 800 658 847
rect 716 847 899 864
rect 933 864 969 881
rect 933 847 1116 864
rect 716 800 1116 847
rect -1116 -847 -716 -800
rect -1116 -864 -933 -847
rect -969 -881 -933 -864
rect -899 -864 -716 -847
rect -658 -847 -258 -800
rect -658 -864 -475 -847
rect -899 -881 -863 -864
rect -969 -897 -863 -881
rect -511 -881 -475 -864
rect -441 -864 -258 -847
rect -200 -847 200 -800
rect -200 -864 -17 -847
rect -441 -881 -405 -864
rect -511 -897 -405 -881
rect -53 -881 -17 -864
rect 17 -864 200 -847
rect 258 -847 658 -800
rect 258 -864 441 -847
rect 17 -881 53 -864
rect -53 -897 53 -881
rect 405 -881 441 -864
rect 475 -864 658 -847
rect 716 -847 1116 -800
rect 716 -864 899 -847
rect 475 -881 511 -864
rect 405 -897 511 -881
rect 863 -881 899 -864
rect 933 -864 1116 -847
rect 933 -881 969 -864
rect 863 -897 969 -881
<< polycont >>
rect -933 847 -899 881
rect -475 847 -441 881
rect -17 847 17 881
rect 441 847 475 881
rect 899 847 933 881
rect -933 -881 -899 -847
rect -475 -881 -441 -847
rect -17 -881 17 -847
rect 441 -881 475 -847
rect 899 -881 933 -847
<< locali >>
rect -1276 949 -1241 983
rect -1207 949 -1173 983
rect -1135 949 -1105 983
rect -1063 949 -1037 983
rect -991 949 -969 983
rect -919 949 -901 983
rect -847 949 -833 983
rect -775 949 -765 983
rect -703 949 -697 983
rect -631 949 -629 983
rect -595 949 -593 983
rect -527 949 -521 983
rect -459 949 -449 983
rect -391 949 -377 983
rect -323 949 -305 983
rect -255 949 -233 983
rect -187 949 -161 983
rect -119 949 -89 983
rect -51 949 -17 983
rect 17 949 51 983
rect 89 949 119 983
rect 161 949 187 983
rect 233 949 255 983
rect 305 949 323 983
rect 377 949 391 983
rect 449 949 459 983
rect 521 949 527 983
rect 593 949 595 983
rect 629 949 631 983
rect 697 949 703 983
rect 765 949 775 983
rect 833 949 847 983
rect 901 949 919 983
rect 969 949 991 983
rect 1037 949 1063 983
rect 1105 949 1135 983
rect 1173 949 1207 983
rect 1241 949 1276 983
rect -1276 867 -1242 949
rect -969 847 -933 881
rect -899 847 -863 881
rect -511 847 -475 881
rect -441 847 -405 881
rect -53 847 -17 881
rect 17 847 53 881
rect 405 847 441 881
rect 475 847 511 881
rect 863 847 899 881
rect 933 847 969 881
rect 1242 867 1276 949
rect -1276 799 -1242 833
rect -1276 731 -1242 765
rect -1276 663 -1242 697
rect -1276 595 -1242 629
rect -1276 527 -1242 561
rect -1276 459 -1242 493
rect -1276 391 -1242 425
rect -1276 323 -1242 357
rect -1276 255 -1242 289
rect -1276 187 -1242 221
rect -1276 119 -1242 153
rect -1276 51 -1242 85
rect -1276 -17 -1242 17
rect -1276 -85 -1242 -51
rect -1276 -153 -1242 -119
rect -1276 -221 -1242 -187
rect -1276 -289 -1242 -255
rect -1276 -357 -1242 -323
rect -1276 -425 -1242 -391
rect -1276 -493 -1242 -459
rect -1276 -561 -1242 -527
rect -1276 -629 -1242 -595
rect -1276 -697 -1242 -663
rect -1276 -765 -1242 -731
rect -1276 -833 -1242 -799
rect -1162 773 -1128 804
rect -1162 701 -1128 731
rect -1162 629 -1128 663
rect -1162 561 -1128 595
rect -1162 493 -1128 523
rect -1162 425 -1128 451
rect -1162 357 -1128 379
rect -1162 289 -1128 307
rect -1162 221 -1128 235
rect -1162 153 -1128 163
rect -1162 85 -1128 91
rect -1162 17 -1128 19
rect -1162 -19 -1128 -17
rect -1162 -91 -1128 -85
rect -1162 -163 -1128 -153
rect -1162 -235 -1128 -221
rect -1162 -307 -1128 -289
rect -1162 -379 -1128 -357
rect -1162 -451 -1128 -425
rect -1162 -523 -1128 -493
rect -1162 -595 -1128 -561
rect -1162 -663 -1128 -629
rect -1162 -731 -1128 -701
rect -1162 -804 -1128 -773
rect -704 773 -670 804
rect -704 701 -670 731
rect -704 629 -670 663
rect -704 561 -670 595
rect -704 493 -670 523
rect -704 425 -670 451
rect -704 357 -670 379
rect -704 289 -670 307
rect -704 221 -670 235
rect -704 153 -670 163
rect -704 85 -670 91
rect -704 17 -670 19
rect -704 -19 -670 -17
rect -704 -91 -670 -85
rect -704 -163 -670 -153
rect -704 -235 -670 -221
rect -704 -307 -670 -289
rect -704 -379 -670 -357
rect -704 -451 -670 -425
rect -704 -523 -670 -493
rect -704 -595 -670 -561
rect -704 -663 -670 -629
rect -704 -731 -670 -701
rect -704 -804 -670 -773
rect -246 773 -212 804
rect -246 701 -212 731
rect -246 629 -212 663
rect -246 561 -212 595
rect -246 493 -212 523
rect -246 425 -212 451
rect -246 357 -212 379
rect -246 289 -212 307
rect -246 221 -212 235
rect -246 153 -212 163
rect -246 85 -212 91
rect -246 17 -212 19
rect -246 -19 -212 -17
rect -246 -91 -212 -85
rect -246 -163 -212 -153
rect -246 -235 -212 -221
rect -246 -307 -212 -289
rect -246 -379 -212 -357
rect -246 -451 -212 -425
rect -246 -523 -212 -493
rect -246 -595 -212 -561
rect -246 -663 -212 -629
rect -246 -731 -212 -701
rect -246 -804 -212 -773
rect 212 773 246 804
rect 212 701 246 731
rect 212 629 246 663
rect 212 561 246 595
rect 212 493 246 523
rect 212 425 246 451
rect 212 357 246 379
rect 212 289 246 307
rect 212 221 246 235
rect 212 153 246 163
rect 212 85 246 91
rect 212 17 246 19
rect 212 -19 246 -17
rect 212 -91 246 -85
rect 212 -163 246 -153
rect 212 -235 246 -221
rect 212 -307 246 -289
rect 212 -379 246 -357
rect 212 -451 246 -425
rect 212 -523 246 -493
rect 212 -595 246 -561
rect 212 -663 246 -629
rect 212 -731 246 -701
rect 212 -804 246 -773
rect 670 773 704 804
rect 670 701 704 731
rect 670 629 704 663
rect 670 561 704 595
rect 670 493 704 523
rect 670 425 704 451
rect 670 357 704 379
rect 670 289 704 307
rect 670 221 704 235
rect 670 153 704 163
rect 670 85 704 91
rect 670 17 704 19
rect 670 -19 704 -17
rect 670 -91 704 -85
rect 670 -163 704 -153
rect 670 -235 704 -221
rect 670 -307 704 -289
rect 670 -379 704 -357
rect 670 -451 704 -425
rect 670 -523 704 -493
rect 670 -595 704 -561
rect 670 -663 704 -629
rect 670 -731 704 -701
rect 670 -804 704 -773
rect 1128 773 1162 804
rect 1128 701 1162 731
rect 1128 629 1162 663
rect 1128 561 1162 595
rect 1128 493 1162 523
rect 1128 425 1162 451
rect 1128 357 1162 379
rect 1128 289 1162 307
rect 1128 221 1162 235
rect 1128 153 1162 163
rect 1128 85 1162 91
rect 1128 17 1162 19
rect 1128 -19 1162 -17
rect 1128 -91 1162 -85
rect 1128 -163 1162 -153
rect 1128 -235 1162 -221
rect 1128 -307 1162 -289
rect 1128 -379 1162 -357
rect 1128 -451 1162 -425
rect 1128 -523 1162 -493
rect 1128 -595 1162 -561
rect 1128 -663 1162 -629
rect 1128 -731 1162 -701
rect 1128 -804 1162 -773
rect 1242 799 1276 833
rect 1242 731 1276 765
rect 1242 663 1276 697
rect 1242 595 1276 629
rect 1242 527 1276 561
rect 1242 459 1276 493
rect 1242 391 1276 425
rect 1242 323 1276 357
rect 1242 255 1276 289
rect 1242 187 1276 221
rect 1242 119 1276 153
rect 1242 51 1276 85
rect 1242 -17 1276 17
rect 1242 -85 1276 -51
rect 1242 -153 1276 -119
rect 1242 -221 1276 -187
rect 1242 -289 1276 -255
rect 1242 -357 1276 -323
rect 1242 -425 1276 -391
rect 1242 -493 1276 -459
rect 1242 -561 1276 -527
rect 1242 -629 1276 -595
rect 1242 -697 1276 -663
rect 1242 -765 1276 -731
rect 1242 -833 1276 -799
rect -1276 -949 -1242 -867
rect -969 -881 -933 -847
rect -899 -881 -863 -847
rect -511 -881 -475 -847
rect -441 -881 -405 -847
rect -53 -881 -17 -847
rect 17 -881 53 -847
rect 405 -881 441 -847
rect 475 -881 511 -847
rect 863 -881 899 -847
rect 933 -881 969 -847
rect 1242 -949 1276 -867
rect -1276 -983 -1173 -949
rect -1139 -983 -1105 -949
rect -1071 -983 -1037 -949
rect -1003 -983 -969 -949
rect -935 -983 -901 -949
rect -867 -983 -833 -949
rect -799 -983 -765 -949
rect -731 -983 -697 -949
rect -663 -983 -629 -949
rect -595 -983 -561 -949
rect -527 -983 -493 -949
rect -459 -983 -425 -949
rect -391 -983 -357 -949
rect -323 -983 -289 -949
rect -255 -983 -221 -949
rect -187 -983 -153 -949
rect -119 -983 -85 -949
rect -51 -983 -17 -949
rect 17 -983 51 -949
rect 85 -983 119 -949
rect 153 -983 187 -949
rect 221 -983 255 -949
rect 289 -983 323 -949
rect 357 -983 391 -949
rect 425 -983 459 -949
rect 493 -983 527 -949
rect 561 -983 595 -949
rect 629 -983 663 -949
rect 697 -983 731 -949
rect 765 -983 799 -949
rect 833 -983 867 -949
rect 901 -983 935 -949
rect 969 -983 1003 -949
rect 1037 -983 1071 -949
rect 1105 -983 1139 -949
rect 1173 -983 1276 -949
<< viali >>
rect -1241 949 -1207 983
rect -1169 949 -1139 983
rect -1139 949 -1135 983
rect -1097 949 -1071 983
rect -1071 949 -1063 983
rect -1025 949 -1003 983
rect -1003 949 -991 983
rect -953 949 -935 983
rect -935 949 -919 983
rect -881 949 -867 983
rect -867 949 -847 983
rect -809 949 -799 983
rect -799 949 -775 983
rect -737 949 -731 983
rect -731 949 -703 983
rect -665 949 -663 983
rect -663 949 -631 983
rect -593 949 -561 983
rect -561 949 -559 983
rect -521 949 -493 983
rect -493 949 -487 983
rect -449 949 -425 983
rect -425 949 -415 983
rect -377 949 -357 983
rect -357 949 -343 983
rect -305 949 -289 983
rect -289 949 -271 983
rect -233 949 -221 983
rect -221 949 -199 983
rect -161 949 -153 983
rect -153 949 -127 983
rect -89 949 -85 983
rect -85 949 -55 983
rect -17 949 17 983
rect 55 949 85 983
rect 85 949 89 983
rect 127 949 153 983
rect 153 949 161 983
rect 199 949 221 983
rect 221 949 233 983
rect 271 949 289 983
rect 289 949 305 983
rect 343 949 357 983
rect 357 949 377 983
rect 415 949 425 983
rect 425 949 449 983
rect 487 949 493 983
rect 493 949 521 983
rect 559 949 561 983
rect 561 949 593 983
rect 631 949 663 983
rect 663 949 665 983
rect 703 949 731 983
rect 731 949 737 983
rect 775 949 799 983
rect 799 949 809 983
rect 847 949 867 983
rect 867 949 881 983
rect 919 949 935 983
rect 935 949 953 983
rect 991 949 1003 983
rect 1003 949 1025 983
rect 1063 949 1071 983
rect 1071 949 1097 983
rect 1135 949 1139 983
rect 1139 949 1169 983
rect 1207 949 1241 983
rect -1162 765 -1128 773
rect -1162 739 -1128 765
rect -1162 697 -1128 701
rect -1162 667 -1128 697
rect -1162 595 -1128 629
rect -1162 527 -1128 557
rect -1162 523 -1128 527
rect -1162 459 -1128 485
rect -1162 451 -1128 459
rect -1162 391 -1128 413
rect -1162 379 -1128 391
rect -1162 323 -1128 341
rect -1162 307 -1128 323
rect -1162 255 -1128 269
rect -1162 235 -1128 255
rect -1162 187 -1128 197
rect -1162 163 -1128 187
rect -1162 119 -1128 125
rect -1162 91 -1128 119
rect -1162 51 -1128 53
rect -1162 19 -1128 51
rect -1162 -51 -1128 -19
rect -1162 -53 -1128 -51
rect -1162 -119 -1128 -91
rect -1162 -125 -1128 -119
rect -1162 -187 -1128 -163
rect -1162 -197 -1128 -187
rect -1162 -255 -1128 -235
rect -1162 -269 -1128 -255
rect -1162 -323 -1128 -307
rect -1162 -341 -1128 -323
rect -1162 -391 -1128 -379
rect -1162 -413 -1128 -391
rect -1162 -459 -1128 -451
rect -1162 -485 -1128 -459
rect -1162 -527 -1128 -523
rect -1162 -557 -1128 -527
rect -1162 -629 -1128 -595
rect -1162 -697 -1128 -667
rect -1162 -701 -1128 -697
rect -1162 -765 -1128 -739
rect -1162 -773 -1128 -765
rect -704 765 -670 773
rect -704 739 -670 765
rect -704 697 -670 701
rect -704 667 -670 697
rect -704 595 -670 629
rect -704 527 -670 557
rect -704 523 -670 527
rect -704 459 -670 485
rect -704 451 -670 459
rect -704 391 -670 413
rect -704 379 -670 391
rect -704 323 -670 341
rect -704 307 -670 323
rect -704 255 -670 269
rect -704 235 -670 255
rect -704 187 -670 197
rect -704 163 -670 187
rect -704 119 -670 125
rect -704 91 -670 119
rect -704 51 -670 53
rect -704 19 -670 51
rect -704 -51 -670 -19
rect -704 -53 -670 -51
rect -704 -119 -670 -91
rect -704 -125 -670 -119
rect -704 -187 -670 -163
rect -704 -197 -670 -187
rect -704 -255 -670 -235
rect -704 -269 -670 -255
rect -704 -323 -670 -307
rect -704 -341 -670 -323
rect -704 -391 -670 -379
rect -704 -413 -670 -391
rect -704 -459 -670 -451
rect -704 -485 -670 -459
rect -704 -527 -670 -523
rect -704 -557 -670 -527
rect -704 -629 -670 -595
rect -704 -697 -670 -667
rect -704 -701 -670 -697
rect -704 -765 -670 -739
rect -704 -773 -670 -765
rect -246 765 -212 773
rect -246 739 -212 765
rect -246 697 -212 701
rect -246 667 -212 697
rect -246 595 -212 629
rect -246 527 -212 557
rect -246 523 -212 527
rect -246 459 -212 485
rect -246 451 -212 459
rect -246 391 -212 413
rect -246 379 -212 391
rect -246 323 -212 341
rect -246 307 -212 323
rect -246 255 -212 269
rect -246 235 -212 255
rect -246 187 -212 197
rect -246 163 -212 187
rect -246 119 -212 125
rect -246 91 -212 119
rect -246 51 -212 53
rect -246 19 -212 51
rect -246 -51 -212 -19
rect -246 -53 -212 -51
rect -246 -119 -212 -91
rect -246 -125 -212 -119
rect -246 -187 -212 -163
rect -246 -197 -212 -187
rect -246 -255 -212 -235
rect -246 -269 -212 -255
rect -246 -323 -212 -307
rect -246 -341 -212 -323
rect -246 -391 -212 -379
rect -246 -413 -212 -391
rect -246 -459 -212 -451
rect -246 -485 -212 -459
rect -246 -527 -212 -523
rect -246 -557 -212 -527
rect -246 -629 -212 -595
rect -246 -697 -212 -667
rect -246 -701 -212 -697
rect -246 -765 -212 -739
rect -246 -773 -212 -765
rect 212 765 246 773
rect 212 739 246 765
rect 212 697 246 701
rect 212 667 246 697
rect 212 595 246 629
rect 212 527 246 557
rect 212 523 246 527
rect 212 459 246 485
rect 212 451 246 459
rect 212 391 246 413
rect 212 379 246 391
rect 212 323 246 341
rect 212 307 246 323
rect 212 255 246 269
rect 212 235 246 255
rect 212 187 246 197
rect 212 163 246 187
rect 212 119 246 125
rect 212 91 246 119
rect 212 51 246 53
rect 212 19 246 51
rect 212 -51 246 -19
rect 212 -53 246 -51
rect 212 -119 246 -91
rect 212 -125 246 -119
rect 212 -187 246 -163
rect 212 -197 246 -187
rect 212 -255 246 -235
rect 212 -269 246 -255
rect 212 -323 246 -307
rect 212 -341 246 -323
rect 212 -391 246 -379
rect 212 -413 246 -391
rect 212 -459 246 -451
rect 212 -485 246 -459
rect 212 -527 246 -523
rect 212 -557 246 -527
rect 212 -629 246 -595
rect 212 -697 246 -667
rect 212 -701 246 -697
rect 212 -765 246 -739
rect 212 -773 246 -765
rect 670 765 704 773
rect 670 739 704 765
rect 670 697 704 701
rect 670 667 704 697
rect 670 595 704 629
rect 670 527 704 557
rect 670 523 704 527
rect 670 459 704 485
rect 670 451 704 459
rect 670 391 704 413
rect 670 379 704 391
rect 670 323 704 341
rect 670 307 704 323
rect 670 255 704 269
rect 670 235 704 255
rect 670 187 704 197
rect 670 163 704 187
rect 670 119 704 125
rect 670 91 704 119
rect 670 51 704 53
rect 670 19 704 51
rect 670 -51 704 -19
rect 670 -53 704 -51
rect 670 -119 704 -91
rect 670 -125 704 -119
rect 670 -187 704 -163
rect 670 -197 704 -187
rect 670 -255 704 -235
rect 670 -269 704 -255
rect 670 -323 704 -307
rect 670 -341 704 -323
rect 670 -391 704 -379
rect 670 -413 704 -391
rect 670 -459 704 -451
rect 670 -485 704 -459
rect 670 -527 704 -523
rect 670 -557 704 -527
rect 670 -629 704 -595
rect 670 -697 704 -667
rect 670 -701 704 -697
rect 670 -765 704 -739
rect 670 -773 704 -765
rect 1128 765 1162 773
rect 1128 739 1162 765
rect 1128 697 1162 701
rect 1128 667 1162 697
rect 1128 595 1162 629
rect 1128 527 1162 557
rect 1128 523 1162 527
rect 1128 459 1162 485
rect 1128 451 1162 459
rect 1128 391 1162 413
rect 1128 379 1162 391
rect 1128 323 1162 341
rect 1128 307 1162 323
rect 1128 255 1162 269
rect 1128 235 1162 255
rect 1128 187 1162 197
rect 1128 163 1162 187
rect 1128 119 1162 125
rect 1128 91 1162 119
rect 1128 51 1162 53
rect 1128 19 1162 51
rect 1128 -51 1162 -19
rect 1128 -53 1162 -51
rect 1128 -119 1162 -91
rect 1128 -125 1162 -119
rect 1128 -187 1162 -163
rect 1128 -197 1162 -187
rect 1128 -255 1162 -235
rect 1128 -269 1162 -255
rect 1128 -323 1162 -307
rect 1128 -341 1162 -323
rect 1128 -391 1162 -379
rect 1128 -413 1162 -391
rect 1128 -459 1162 -451
rect 1128 -485 1162 -459
rect 1128 -527 1162 -523
rect 1128 -557 1162 -527
rect 1128 -629 1162 -595
rect 1128 -697 1162 -667
rect 1128 -701 1162 -697
rect 1128 -765 1162 -739
rect 1128 -773 1162 -765
<< metal1 >>
rect -1254 983 1254 989
rect -1254 949 -1241 983
rect -1207 949 -1169 983
rect -1135 949 -1097 983
rect -1063 949 -1025 983
rect -991 949 -953 983
rect -919 949 -881 983
rect -847 949 -809 983
rect -775 949 -737 983
rect -703 949 -665 983
rect -631 949 -593 983
rect -559 949 -521 983
rect -487 949 -449 983
rect -415 949 -377 983
rect -343 949 -305 983
rect -271 949 -233 983
rect -199 949 -161 983
rect -127 949 -89 983
rect -55 949 -17 983
rect 17 949 55 983
rect 89 949 127 983
rect 161 949 199 983
rect 233 949 271 983
rect 305 949 343 983
rect 377 949 415 983
rect 449 949 487 983
rect 521 949 559 983
rect 593 949 631 983
rect 665 949 703 983
rect 737 949 775 983
rect 809 949 847 983
rect 881 949 919 983
rect 953 949 991 983
rect 1025 949 1063 983
rect 1097 949 1135 983
rect 1169 949 1207 983
rect 1241 949 1254 983
rect -1254 943 1254 949
rect -1168 773 -1122 800
rect -1168 739 -1162 773
rect -1128 739 -1122 773
rect -1168 701 -1122 739
rect -1168 667 -1162 701
rect -1128 667 -1122 701
rect -1168 629 -1122 667
rect -1168 595 -1162 629
rect -1128 595 -1122 629
rect -1168 557 -1122 595
rect -1168 523 -1162 557
rect -1128 523 -1122 557
rect -1168 485 -1122 523
rect -1168 451 -1162 485
rect -1128 451 -1122 485
rect -1168 413 -1122 451
rect -1168 379 -1162 413
rect -1128 379 -1122 413
rect -1168 341 -1122 379
rect -1168 307 -1162 341
rect -1128 307 -1122 341
rect -1168 269 -1122 307
rect -1168 235 -1162 269
rect -1128 235 -1122 269
rect -1168 197 -1122 235
rect -1168 163 -1162 197
rect -1128 163 -1122 197
rect -1168 125 -1122 163
rect -1168 91 -1162 125
rect -1128 91 -1122 125
rect -1168 53 -1122 91
rect -1168 19 -1162 53
rect -1128 19 -1122 53
rect -1168 -19 -1122 19
rect -1168 -53 -1162 -19
rect -1128 -53 -1122 -19
rect -1168 -91 -1122 -53
rect -1168 -125 -1162 -91
rect -1128 -125 -1122 -91
rect -1168 -163 -1122 -125
rect -1168 -197 -1162 -163
rect -1128 -197 -1122 -163
rect -1168 -235 -1122 -197
rect -1168 -269 -1162 -235
rect -1128 -269 -1122 -235
rect -1168 -307 -1122 -269
rect -1168 -341 -1162 -307
rect -1128 -341 -1122 -307
rect -1168 -379 -1122 -341
rect -1168 -413 -1162 -379
rect -1128 -413 -1122 -379
rect -1168 -451 -1122 -413
rect -1168 -485 -1162 -451
rect -1128 -485 -1122 -451
rect -1168 -523 -1122 -485
rect -1168 -557 -1162 -523
rect -1128 -557 -1122 -523
rect -1168 -595 -1122 -557
rect -1168 -629 -1162 -595
rect -1128 -629 -1122 -595
rect -1168 -667 -1122 -629
rect -1168 -701 -1162 -667
rect -1128 -701 -1122 -667
rect -1168 -739 -1122 -701
rect -1168 -773 -1162 -739
rect -1128 -773 -1122 -739
rect -1168 -800 -1122 -773
rect -710 773 -664 800
rect -710 739 -704 773
rect -670 739 -664 773
rect -710 701 -664 739
rect -710 667 -704 701
rect -670 667 -664 701
rect -710 629 -664 667
rect -710 595 -704 629
rect -670 595 -664 629
rect -710 557 -664 595
rect -710 523 -704 557
rect -670 523 -664 557
rect -710 485 -664 523
rect -710 451 -704 485
rect -670 451 -664 485
rect -710 413 -664 451
rect -710 379 -704 413
rect -670 379 -664 413
rect -710 341 -664 379
rect -710 307 -704 341
rect -670 307 -664 341
rect -710 269 -664 307
rect -710 235 -704 269
rect -670 235 -664 269
rect -710 197 -664 235
rect -710 163 -704 197
rect -670 163 -664 197
rect -710 125 -664 163
rect -710 91 -704 125
rect -670 91 -664 125
rect -710 53 -664 91
rect -710 19 -704 53
rect -670 19 -664 53
rect -710 -19 -664 19
rect -710 -53 -704 -19
rect -670 -53 -664 -19
rect -710 -91 -664 -53
rect -710 -125 -704 -91
rect -670 -125 -664 -91
rect -710 -163 -664 -125
rect -710 -197 -704 -163
rect -670 -197 -664 -163
rect -710 -235 -664 -197
rect -710 -269 -704 -235
rect -670 -269 -664 -235
rect -710 -307 -664 -269
rect -710 -341 -704 -307
rect -670 -341 -664 -307
rect -710 -379 -664 -341
rect -710 -413 -704 -379
rect -670 -413 -664 -379
rect -710 -451 -664 -413
rect -710 -485 -704 -451
rect -670 -485 -664 -451
rect -710 -523 -664 -485
rect -710 -557 -704 -523
rect -670 -557 -664 -523
rect -710 -595 -664 -557
rect -710 -629 -704 -595
rect -670 -629 -664 -595
rect -710 -667 -664 -629
rect -710 -701 -704 -667
rect -670 -701 -664 -667
rect -710 -739 -664 -701
rect -710 -773 -704 -739
rect -670 -773 -664 -739
rect -710 -800 -664 -773
rect -252 773 -206 800
rect -252 739 -246 773
rect -212 739 -206 773
rect -252 701 -206 739
rect -252 667 -246 701
rect -212 667 -206 701
rect -252 629 -206 667
rect -252 595 -246 629
rect -212 595 -206 629
rect -252 557 -206 595
rect -252 523 -246 557
rect -212 523 -206 557
rect -252 485 -206 523
rect -252 451 -246 485
rect -212 451 -206 485
rect -252 413 -206 451
rect -252 379 -246 413
rect -212 379 -206 413
rect -252 341 -206 379
rect -252 307 -246 341
rect -212 307 -206 341
rect -252 269 -206 307
rect -252 235 -246 269
rect -212 235 -206 269
rect -252 197 -206 235
rect -252 163 -246 197
rect -212 163 -206 197
rect -252 125 -206 163
rect -252 91 -246 125
rect -212 91 -206 125
rect -252 53 -206 91
rect -252 19 -246 53
rect -212 19 -206 53
rect -252 -19 -206 19
rect -252 -53 -246 -19
rect -212 -53 -206 -19
rect -252 -91 -206 -53
rect -252 -125 -246 -91
rect -212 -125 -206 -91
rect -252 -163 -206 -125
rect -252 -197 -246 -163
rect -212 -197 -206 -163
rect -252 -235 -206 -197
rect -252 -269 -246 -235
rect -212 -269 -206 -235
rect -252 -307 -206 -269
rect -252 -341 -246 -307
rect -212 -341 -206 -307
rect -252 -379 -206 -341
rect -252 -413 -246 -379
rect -212 -413 -206 -379
rect -252 -451 -206 -413
rect -252 -485 -246 -451
rect -212 -485 -206 -451
rect -252 -523 -206 -485
rect -252 -557 -246 -523
rect -212 -557 -206 -523
rect -252 -595 -206 -557
rect -252 -629 -246 -595
rect -212 -629 -206 -595
rect -252 -667 -206 -629
rect -252 -701 -246 -667
rect -212 -701 -206 -667
rect -252 -739 -206 -701
rect -252 -773 -246 -739
rect -212 -773 -206 -739
rect -252 -800 -206 -773
rect 206 773 252 800
rect 206 739 212 773
rect 246 739 252 773
rect 206 701 252 739
rect 206 667 212 701
rect 246 667 252 701
rect 206 629 252 667
rect 206 595 212 629
rect 246 595 252 629
rect 206 557 252 595
rect 206 523 212 557
rect 246 523 252 557
rect 206 485 252 523
rect 206 451 212 485
rect 246 451 252 485
rect 206 413 252 451
rect 206 379 212 413
rect 246 379 252 413
rect 206 341 252 379
rect 206 307 212 341
rect 246 307 252 341
rect 206 269 252 307
rect 206 235 212 269
rect 246 235 252 269
rect 206 197 252 235
rect 206 163 212 197
rect 246 163 252 197
rect 206 125 252 163
rect 206 91 212 125
rect 246 91 252 125
rect 206 53 252 91
rect 206 19 212 53
rect 246 19 252 53
rect 206 -19 252 19
rect 206 -53 212 -19
rect 246 -53 252 -19
rect 206 -91 252 -53
rect 206 -125 212 -91
rect 246 -125 252 -91
rect 206 -163 252 -125
rect 206 -197 212 -163
rect 246 -197 252 -163
rect 206 -235 252 -197
rect 206 -269 212 -235
rect 246 -269 252 -235
rect 206 -307 252 -269
rect 206 -341 212 -307
rect 246 -341 252 -307
rect 206 -379 252 -341
rect 206 -413 212 -379
rect 246 -413 252 -379
rect 206 -451 252 -413
rect 206 -485 212 -451
rect 246 -485 252 -451
rect 206 -523 252 -485
rect 206 -557 212 -523
rect 246 -557 252 -523
rect 206 -595 252 -557
rect 206 -629 212 -595
rect 246 -629 252 -595
rect 206 -667 252 -629
rect 206 -701 212 -667
rect 246 -701 252 -667
rect 206 -739 252 -701
rect 206 -773 212 -739
rect 246 -773 252 -739
rect 206 -800 252 -773
rect 664 773 710 800
rect 664 739 670 773
rect 704 739 710 773
rect 664 701 710 739
rect 664 667 670 701
rect 704 667 710 701
rect 664 629 710 667
rect 664 595 670 629
rect 704 595 710 629
rect 664 557 710 595
rect 664 523 670 557
rect 704 523 710 557
rect 664 485 710 523
rect 664 451 670 485
rect 704 451 710 485
rect 664 413 710 451
rect 664 379 670 413
rect 704 379 710 413
rect 664 341 710 379
rect 664 307 670 341
rect 704 307 710 341
rect 664 269 710 307
rect 664 235 670 269
rect 704 235 710 269
rect 664 197 710 235
rect 664 163 670 197
rect 704 163 710 197
rect 664 125 710 163
rect 664 91 670 125
rect 704 91 710 125
rect 664 53 710 91
rect 664 19 670 53
rect 704 19 710 53
rect 664 -19 710 19
rect 664 -53 670 -19
rect 704 -53 710 -19
rect 664 -91 710 -53
rect 664 -125 670 -91
rect 704 -125 710 -91
rect 664 -163 710 -125
rect 664 -197 670 -163
rect 704 -197 710 -163
rect 664 -235 710 -197
rect 664 -269 670 -235
rect 704 -269 710 -235
rect 664 -307 710 -269
rect 664 -341 670 -307
rect 704 -341 710 -307
rect 664 -379 710 -341
rect 664 -413 670 -379
rect 704 -413 710 -379
rect 664 -451 710 -413
rect 664 -485 670 -451
rect 704 -485 710 -451
rect 664 -523 710 -485
rect 664 -557 670 -523
rect 704 -557 710 -523
rect 664 -595 710 -557
rect 664 -629 670 -595
rect 704 -629 710 -595
rect 664 -667 710 -629
rect 664 -701 670 -667
rect 704 -701 710 -667
rect 664 -739 710 -701
rect 664 -773 670 -739
rect 704 -773 710 -739
rect 664 -800 710 -773
rect 1122 773 1168 800
rect 1122 739 1128 773
rect 1162 739 1168 773
rect 1122 701 1168 739
rect 1122 667 1128 701
rect 1162 667 1168 701
rect 1122 629 1168 667
rect 1122 595 1128 629
rect 1162 595 1168 629
rect 1122 557 1168 595
rect 1122 523 1128 557
rect 1162 523 1168 557
rect 1122 485 1168 523
rect 1122 451 1128 485
rect 1162 451 1168 485
rect 1122 413 1168 451
rect 1122 379 1128 413
rect 1162 379 1168 413
rect 1122 341 1168 379
rect 1122 307 1128 341
rect 1162 307 1168 341
rect 1122 269 1168 307
rect 1122 235 1128 269
rect 1162 235 1168 269
rect 1122 197 1168 235
rect 1122 163 1128 197
rect 1162 163 1168 197
rect 1122 125 1168 163
rect 1122 91 1128 125
rect 1162 91 1168 125
rect 1122 53 1168 91
rect 1122 19 1128 53
rect 1162 19 1168 53
rect 1122 -19 1168 19
rect 1122 -53 1128 -19
rect 1162 -53 1168 -19
rect 1122 -91 1168 -53
rect 1122 -125 1128 -91
rect 1162 -125 1168 -91
rect 1122 -163 1168 -125
rect 1122 -197 1128 -163
rect 1162 -197 1168 -163
rect 1122 -235 1168 -197
rect 1122 -269 1128 -235
rect 1162 -269 1168 -235
rect 1122 -307 1168 -269
rect 1122 -341 1128 -307
rect 1162 -341 1168 -307
rect 1122 -379 1168 -341
rect 1122 -413 1128 -379
rect 1162 -413 1168 -379
rect 1122 -451 1168 -413
rect 1122 -485 1128 -451
rect 1162 -485 1168 -451
rect 1122 -523 1168 -485
rect 1122 -557 1128 -523
rect 1162 -557 1168 -523
rect 1122 -595 1168 -557
rect 1122 -629 1128 -595
rect 1162 -629 1168 -595
rect 1122 -667 1168 -629
rect 1122 -701 1128 -667
rect 1162 -701 1168 -667
rect 1122 -739 1168 -701
rect 1122 -773 1128 -739
rect 1162 -773 1168 -739
rect 1122 -800 1168 -773
<< properties >>
string FIXED_BBOX -1259 -966 1259 966
<< end >>
