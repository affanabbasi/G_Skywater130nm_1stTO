magic
tech sky130A
timestamp 1608072493
<< error_p >>
rect 8 -352 9 352
<< pwell >>
rect -1228 -455 1228 455
<< nmoslvt >>
rect -1130 -350 -930 350
rect -901 -350 -701 350
rect -672 -350 -472 350
rect -443 -350 -243 350
rect -214 -350 -14 350
rect 14 -350 214 350
rect 243 -350 443 350
rect 472 -350 672 350
rect 701 -350 901 350
rect 930 -350 1130 350
<< ndiff >>
rect -1159 344 -1130 350
rect -1159 -344 -1153 344
rect -1136 -344 -1130 344
rect -1159 -350 -1130 -344
rect -930 344 -901 350
rect -930 -344 -924 344
rect -907 -344 -901 344
rect -930 -350 -901 -344
rect -701 344 -672 350
rect -701 -344 -695 344
rect -678 -344 -672 344
rect -701 -350 -672 -344
rect -472 344 -443 350
rect -472 -344 -466 344
rect -449 -344 -443 344
rect -472 -350 -443 -344
rect -243 344 -214 350
rect -243 -344 -237 344
rect -220 -344 -214 344
rect -243 -350 -214 -344
rect -14 344 14 350
rect -14 -344 -8 344
rect 8 -344 14 344
rect -14 -350 14 -344
rect 214 344 243 350
rect 214 -344 220 344
rect 237 -344 243 344
rect 214 -350 243 -344
rect 443 344 472 350
rect 443 -344 449 344
rect 466 -344 472 344
rect 443 -350 472 -344
rect 672 344 701 350
rect 672 -344 678 344
rect 695 -344 701 344
rect 672 -350 701 -344
rect 901 344 930 350
rect 901 -344 907 344
rect 924 -344 930 344
rect 901 -350 930 -344
rect 1130 344 1159 350
rect 1130 -344 1136 344
rect 1153 -344 1159 344
rect 1130 -350 1159 -344
<< ndiffc >>
rect -1153 -344 -1136 344
rect -924 -344 -907 344
rect -695 -344 -678 344
rect -466 -344 -449 344
rect -237 -344 -220 344
rect -8 -344 8 344
rect 220 -344 237 344
rect 449 -344 466 344
rect 678 -344 695 344
rect 907 -344 924 344
rect 1136 -344 1153 344
<< psubdiff >>
rect -1210 420 -1162 437
rect 1162 420 1210 437
rect -1210 389 -1193 420
rect 1193 389 1210 420
rect -1210 -420 -1193 -389
rect 1193 -420 1210 -389
rect -1210 -437 -1162 -420
rect 1162 -437 1210 -420
<< psubdiffcont >>
rect -1162 420 1162 437
rect -1210 -389 -1193 389
rect 1193 -389 1210 389
rect -1162 -437 1162 -420
<< poly >>
rect -1130 386 -930 394
rect -1130 369 -1122 386
rect -938 369 -930 386
rect -1130 350 -930 369
rect -901 386 -701 394
rect -901 369 -893 386
rect -709 369 -701 386
rect -901 350 -701 369
rect -672 386 -472 394
rect -672 369 -664 386
rect -480 369 -472 386
rect -672 350 -472 369
rect -443 386 -243 394
rect -443 369 -435 386
rect -251 369 -243 386
rect -443 350 -243 369
rect -214 386 -14 394
rect -214 369 -206 386
rect -22 369 -14 386
rect -214 350 -14 369
rect 14 386 214 394
rect 14 369 22 386
rect 206 369 214 386
rect 14 350 214 369
rect 243 386 443 394
rect 243 369 251 386
rect 435 369 443 386
rect 243 350 443 369
rect 472 386 672 394
rect 472 369 480 386
rect 664 369 672 386
rect 472 350 672 369
rect 701 386 901 394
rect 701 369 709 386
rect 893 369 901 386
rect 701 350 901 369
rect 930 386 1130 394
rect 930 369 938 386
rect 1122 369 1130 386
rect 930 350 1130 369
rect -1130 -369 -930 -350
rect -1130 -386 -1122 -369
rect -938 -386 -930 -369
rect -1130 -394 -930 -386
rect -901 -369 -701 -350
rect -901 -386 -893 -369
rect -709 -386 -701 -369
rect -901 -394 -701 -386
rect -672 -369 -472 -350
rect -672 -386 -664 -369
rect -480 -386 -472 -369
rect -672 -394 -472 -386
rect -443 -369 -243 -350
rect -443 -386 -435 -369
rect -251 -386 -243 -369
rect -443 -394 -243 -386
rect -214 -369 -14 -350
rect -214 -386 -206 -369
rect -22 -386 -14 -369
rect -214 -394 -14 -386
rect 14 -369 214 -350
rect 14 -386 22 -369
rect 206 -386 214 -369
rect 14 -394 214 -386
rect 243 -369 443 -350
rect 243 -386 251 -369
rect 435 -386 443 -369
rect 243 -394 443 -386
rect 472 -369 672 -350
rect 472 -386 480 -369
rect 664 -386 672 -369
rect 472 -394 672 -386
rect 701 -369 901 -350
rect 701 -386 709 -369
rect 893 -386 901 -369
rect 701 -394 901 -386
rect 930 -369 1130 -350
rect 930 -386 938 -369
rect 1122 -386 1130 -369
rect 930 -394 1130 -386
<< polycont >>
rect -1122 369 -938 386
rect -893 369 -709 386
rect -664 369 -480 386
rect -435 369 -251 386
rect -206 369 -22 386
rect 22 369 206 386
rect 251 369 435 386
rect 480 369 664 386
rect 709 369 893 386
rect 938 369 1122 386
rect -1122 -386 -938 -369
rect -893 -386 -709 -369
rect -664 -386 -480 -369
rect -435 -386 -251 -369
rect -206 -386 -22 -369
rect 22 -386 206 -369
rect 251 -386 435 -369
rect 480 -386 664 -369
rect 709 -386 893 -369
rect 938 -386 1122 -369
<< locali >>
rect -1210 420 -1162 437
rect 1162 420 1210 437
rect -1210 389 -1193 420
rect 1193 389 1210 420
rect -1130 369 -1122 386
rect -938 369 -930 386
rect -901 369 -893 386
rect -709 369 -701 386
rect -672 369 -664 386
rect -480 369 -472 386
rect -443 369 -435 386
rect -251 369 -243 386
rect -214 369 -206 386
rect -22 369 -14 386
rect 14 369 22 386
rect 206 369 214 386
rect 243 369 251 386
rect 435 369 443 386
rect 472 369 480 386
rect 664 369 672 386
rect 701 369 709 386
rect 893 369 901 386
rect 930 369 938 386
rect 1122 369 1130 386
rect -1153 344 -1136 352
rect -1153 -352 -1136 -344
rect -924 344 -907 352
rect -924 -352 -907 -344
rect -695 344 -678 352
rect -695 -352 -678 -344
rect -466 344 -449 352
rect -466 -352 -449 -344
rect -237 344 -220 352
rect -237 -352 -220 -344
rect -8 344 8 352
rect -8 -352 8 -344
rect 220 344 237 352
rect 220 -352 237 -344
rect 449 344 466 352
rect 449 -352 466 -344
rect 678 344 695 352
rect 678 -352 695 -344
rect 907 344 924 352
rect 907 -352 924 -344
rect 1136 344 1153 352
rect 1136 -352 1153 -344
rect -1130 -386 -1122 -369
rect -938 -386 -930 -369
rect -901 -386 -893 -369
rect -709 -386 -701 -369
rect -672 -386 -664 -369
rect -480 -386 -472 -369
rect -443 -386 -435 -369
rect -251 -386 -243 -369
rect -214 -386 -206 -369
rect -22 -386 -14 -369
rect 14 -386 22 -369
rect 206 -386 214 -369
rect 243 -386 251 -369
rect 435 -386 443 -369
rect 472 -386 480 -369
rect 664 -386 672 -369
rect 701 -386 709 -369
rect 893 -386 901 -369
rect 930 -386 938 -369
rect 1122 -386 1130 -369
rect -1210 -420 -1193 -389
rect 1193 -420 1210 -389
rect -1210 -437 -1162 -420
rect 1162 -437 1210 -420
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -1202 -428 1202 428
string parameters w 7 l 2 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1
string library sky130
<< end >>
