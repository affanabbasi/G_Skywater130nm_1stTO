magic
tech sky130A
magscale 1 2
timestamp 1607661548
<< metal1 >>
rect -32 140 32 192
rect -32 -188 32 -136
use sky130_fd_pr__pfet_01v8_lvt_YTP334  sky130_fd_pr__pfet_01v8_lvt_YTP334_0
timestamp 1607661548
transform 1 0 1 0 1 1
box -231 -319 231 319
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -178 -266 178 266
string parameters w 1 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
